
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_pc, ABINPUT, ABINPUT000, ABINPUT001, ABINPUT002, ABINPUT003, ABINPUT004, ABINPUT005, ABINPUT006, ABINPUT007, ABINPUT008, ABINPUT009);
  wire _00000_;
  wire [7:0] _00001_;
  wire _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire [7:0] _29726_;
  wire [7:0] _29727_;
  wire [7:0] _29728_;
  wire [7:0] _29729_;
  wire [7:0] _29730_;
  input [34:0] ABINPUT;
  input [7:0] ABINPUT000;
  input [7:0] ABINPUT001;
  input [7:0] ABINPUT002;
  input [7:0] ABINPUT003;
  input [7:0] ABINPUT004;
  input [7:0] ABINPUT005;
  input [7:0] ABINPUT006;
  input [7:0] ABINPUT007;
  input [7:0] ABINPUT008;
  input [127:0] ABINPUT009;
  wire [7:0] ACC_gm;
  wire [7:0] B_gm;
  wire [7:0] DPH_gm;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IP_gm;
  wire [127:0] IRAM_gm;
  wire [7:0] P0_gm;
  wire [7:0] P1_gm;
  wire [7:0] P2_gm;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PSW_gm;
  wire [7:0] PSW_gm_next;
  wire [7:0] SBUF_gm;
  wire [7:0] SCON_gm;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TH0_gm;
  wire [7:0] TH1_gm;
  wire [7:0] TL0_gm;
  wire [7:0] TL1_gm;
  wire [7:0] TMOD_gm;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire eq_state;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT000 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT001 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT002 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT003 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT004 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT005 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT006 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT007 ;
  wire [127:0] \oc8051_golden_model_1.ABINPUT008 ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_next ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.B_next ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPH_next ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.DPL_next ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [127:0] \oc8051_golden_model_1.IRAM_full ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P0_next ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P1_next ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P2_next ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [7:0] \oc8051_golden_model_1.P3_next ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_fa ;
  wire [7:0] \oc8051_golden_model_1.PSW_fb ;
  wire [7:0] \oc8051_golden_model_1.PSW_fc ;
  wire [7:0] \oc8051_golden_model_1.PSW_fd ;
  wire [7:0] \oc8051_golden_model_1.PSW_fe ;
  wire [7:0] \oc8051_golden_model_1.PSW_ff ;
  wire [7:0] \oc8051_golden_model_1.PSW_next ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0573 ;
  wire [7:0] \oc8051_golden_model_1.n0606 ;
  wire [15:0] \oc8051_golden_model_1.n0713 ;
  wire [15:0] \oc8051_golden_model_1.n0745 ;
  wire [15:0] \oc8051_golden_model_1.n1004 ;
  wire [6:0] \oc8051_golden_model_1.n1008 ;
  wire \oc8051_golden_model_1.n1009 ;
  wire \oc8051_golden_model_1.n1010 ;
  wire \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1023 ;
  wire [7:0] \oc8051_golden_model_1.n1024 ;
  wire [7:0] \oc8051_golden_model_1.n1031 ;
  wire \oc8051_golden_model_1.n1032 ;
  wire \oc8051_golden_model_1.n1033 ;
  wire \oc8051_golden_model_1.n1034 ;
  wire \oc8051_golden_model_1.n1035 ;
  wire \oc8051_golden_model_1.n1036 ;
  wire \oc8051_golden_model_1.n1037 ;
  wire \oc8051_golden_model_1.n1038 ;
  wire \oc8051_golden_model_1.n1039 ;
  wire [7:0] \oc8051_golden_model_1.n1047 ;
  wire [7:0] \oc8051_golden_model_1.n1064 ;
  wire [3:0] \oc8051_golden_model_1.n1157 ;
  wire [3:0] \oc8051_golden_model_1.n1159 ;
  wire [3:0] \oc8051_golden_model_1.n1161 ;
  wire [3:0] \oc8051_golden_model_1.n1162 ;
  wire [3:0] \oc8051_golden_model_1.n1163 ;
  wire [3:0] \oc8051_golden_model_1.n1164 ;
  wire [3:0] \oc8051_golden_model_1.n1165 ;
  wire [3:0] \oc8051_golden_model_1.n1166 ;
  wire [3:0] \oc8051_golden_model_1.n1167 ;
  wire \oc8051_golden_model_1.n1214 ;
  wire \oc8051_golden_model_1.n1259 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [8:0] \oc8051_golden_model_1.n1261 ;
  wire [7:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [2:0] \oc8051_golden_model_1.n1264 ;
  wire \oc8051_golden_model_1.n1265 ;
  wire [1:0] \oc8051_golden_model_1.n1266 ;
  wire [7:0] \oc8051_golden_model_1.n1267 ;
  wire [6:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1269 ;
  wire \oc8051_golden_model_1.n1270 ;
  wire \oc8051_golden_model_1.n1271 ;
  wire \oc8051_golden_model_1.n1272 ;
  wire \oc8051_golden_model_1.n1273 ;
  wire \oc8051_golden_model_1.n1274 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire \oc8051_golden_model_1.n1276 ;
  wire [7:0] \oc8051_golden_model_1.n1284 ;
  wire [7:0] \oc8051_golden_model_1.n1301 ;
  wire [15:0] \oc8051_golden_model_1.n1343 ;
  wire [7:0] \oc8051_golden_model_1.n1345 ;
  wire \oc8051_golden_model_1.n1346 ;
  wire \oc8051_golden_model_1.n1347 ;
  wire \oc8051_golden_model_1.n1348 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire \oc8051_golden_model_1.n1350 ;
  wire \oc8051_golden_model_1.n1351 ;
  wire \oc8051_golden_model_1.n1352 ;
  wire \oc8051_golden_model_1.n1353 ;
  wire \oc8051_golden_model_1.n1360 ;
  wire [7:0] \oc8051_golden_model_1.n1361 ;
  wire [8:0] \oc8051_golden_model_1.n1363 ;
  wire [8:0] \oc8051_golden_model_1.n1367 ;
  wire \oc8051_golden_model_1.n1368 ;
  wire [3:0] \oc8051_golden_model_1.n1369 ;
  wire [4:0] \oc8051_golden_model_1.n1370 ;
  wire [4:0] \oc8051_golden_model_1.n1374 ;
  wire \oc8051_golden_model_1.n1375 ;
  wire [8:0] \oc8051_golden_model_1.n1376 ;
  wire \oc8051_golden_model_1.n1384 ;
  wire [7:0] \oc8051_golden_model_1.n1385 ;
  wire [6:0] \oc8051_golden_model_1.n1386 ;
  wire \oc8051_golden_model_1.n1401 ;
  wire [7:0] \oc8051_golden_model_1.n1402 ;
  wire [8:0] \oc8051_golden_model_1.n1424 ;
  wire \oc8051_golden_model_1.n1425 ;
  wire [4:0] \oc8051_golden_model_1.n1430 ;
  wire \oc8051_golden_model_1.n1431 ;
  wire \oc8051_golden_model_1.n1439 ;
  wire [7:0] \oc8051_golden_model_1.n1440 ;
  wire [6:0] \oc8051_golden_model_1.n1441 ;
  wire \oc8051_golden_model_1.n1456 ;
  wire [7:0] \oc8051_golden_model_1.n1457 ;
  wire [8:0] \oc8051_golden_model_1.n1459 ;
  wire [3:0] \oc8051_golden_model_1.n1463 ;
  wire [4:0] \oc8051_golden_model_1.n1464 ;
  wire [4:0] \oc8051_golden_model_1.n1466 ;
  wire \oc8051_golden_model_1.n1467 ;
  wire [8:0] \oc8051_golden_model_1.n1468 ;
  wire [7:0] \oc8051_golden_model_1.n1476 ;
  wire [6:0] \oc8051_golden_model_1.n1477 ;
  wire \oc8051_golden_model_1.n1492 ;
  wire [7:0] \oc8051_golden_model_1.n1493 ;
  wire [7:0] \oc8051_golden_model_1.n1505 ;
  wire [6:0] \oc8051_golden_model_1.n1506 ;
  wire [7:0] \oc8051_golden_model_1.n1507 ;
  wire [8:0] \oc8051_golden_model_1.n1509 ;
  wire [8:0] \oc8051_golden_model_1.n1511 ;
  wire \oc8051_golden_model_1.n1512 ;
  wire [4:0] \oc8051_golden_model_1.n1513 ;
  wire [4:0] \oc8051_golden_model_1.n1515 ;
  wire \oc8051_golden_model_1.n1516 ;
  wire [8:0] \oc8051_golden_model_1.n1517 ;
  wire \oc8051_golden_model_1.n1524 ;
  wire [7:0] \oc8051_golden_model_1.n1525 ;
  wire [6:0] \oc8051_golden_model_1.n1526 ;
  wire \oc8051_golden_model_1.n1541 ;
  wire [7:0] \oc8051_golden_model_1.n1542 ;
  wire [4:0] \oc8051_golden_model_1.n1544 ;
  wire \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [6:0] \oc8051_golden_model_1.n1547 ;
  wire [7:0] \oc8051_golden_model_1.n1548 ;
  wire [8:0] \oc8051_golden_model_1.n1550 ;
  wire \oc8051_golden_model_1.n1551 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire [7:0] \oc8051_golden_model_1.n1559 ;
  wire [6:0] \oc8051_golden_model_1.n1560 ;
  wire [7:0] \oc8051_golden_model_1.n1561 ;
  wire [7:0] \oc8051_golden_model_1.n1562 ;
  wire [6:0] \oc8051_golden_model_1.n1563 ;
  wire [7:0] \oc8051_golden_model_1.n1564 ;
  wire [8:0] \oc8051_golden_model_1.n1567 ;
  wire [8:0] \oc8051_golden_model_1.n1568 ;
  wire [7:0] \oc8051_golden_model_1.n1569 ;
  wire [7:0] \oc8051_golden_model_1.n1570 ;
  wire [6:0] \oc8051_golden_model_1.n1571 ;
  wire \oc8051_golden_model_1.n1572 ;
  wire \oc8051_golden_model_1.n1573 ;
  wire \oc8051_golden_model_1.n1574 ;
  wire \oc8051_golden_model_1.n1575 ;
  wire \oc8051_golden_model_1.n1576 ;
  wire \oc8051_golden_model_1.n1577 ;
  wire \oc8051_golden_model_1.n1578 ;
  wire \oc8051_golden_model_1.n1579 ;
  wire [7:0] \oc8051_golden_model_1.n1587 ;
  wire [7:0] \oc8051_golden_model_1.n1588 ;
  wire [8:0] \oc8051_golden_model_1.n1591 ;
  wire [4:0] \oc8051_golden_model_1.n1595 ;
  wire [7:0] \oc8051_golden_model_1.n1606 ;
  wire [6:0] \oc8051_golden_model_1.n1607 ;
  wire [7:0] \oc8051_golden_model_1.n1623 ;
  wire [7:0] \oc8051_golden_model_1.n1639 ;
  wire [6:0] \oc8051_golden_model_1.n1640 ;
  wire [7:0] \oc8051_golden_model_1.n1656 ;
  wire [8:0] \oc8051_golden_model_1.n1660 ;
  wire \oc8051_golden_model_1.n1661 ;
  wire [4:0] \oc8051_golden_model_1.n1663 ;
  wire \oc8051_golden_model_1.n1664 ;
  wire \oc8051_golden_model_1.n1671 ;
  wire [7:0] \oc8051_golden_model_1.n1672 ;
  wire [6:0] \oc8051_golden_model_1.n1673 ;
  wire \oc8051_golden_model_1.n1688 ;
  wire [7:0] \oc8051_golden_model_1.n1689 ;
  wire [8:0] \oc8051_golden_model_1.n1693 ;
  wire \oc8051_golden_model_1.n1694 ;
  wire [4:0] \oc8051_golden_model_1.n1696 ;
  wire \oc8051_golden_model_1.n1697 ;
  wire \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1705 ;
  wire [6:0] \oc8051_golden_model_1.n1706 ;
  wire \oc8051_golden_model_1.n1721 ;
  wire [7:0] \oc8051_golden_model_1.n1722 ;
  wire [7:0] \oc8051_golden_model_1.n1749 ;
  wire [7:0] \oc8051_golden_model_1.n1805 ;
  wire [7:0] \oc8051_golden_model_1.n1822 ;
  wire \oc8051_golden_model_1.n1838 ;
  wire [7:0] \oc8051_golden_model_1.n1839 ;
  wire \oc8051_golden_model_1.n1855 ;
  wire [7:0] \oc8051_golden_model_1.n1856 ;
  wire [7:0] \oc8051_golden_model_1.n1881 ;
  wire [7:0] \oc8051_golden_model_1.n1937 ;
  wire [7:0] \oc8051_golden_model_1.n1954 ;
  wire \oc8051_golden_model_1.n1970 ;
  wire [7:0] \oc8051_golden_model_1.n1971 ;
  wire \oc8051_golden_model_1.n1987 ;
  wire [7:0] \oc8051_golden_model_1.n1988 ;
  wire \oc8051_golden_model_1.n2085 ;
  wire [7:0] \oc8051_golden_model_1.n2086 ;
  wire \oc8051_golden_model_1.n2102 ;
  wire [7:0] \oc8051_golden_model_1.n2103 ;
  wire \oc8051_golden_model_1.n2119 ;
  wire [7:0] \oc8051_golden_model_1.n2120 ;
  wire \oc8051_golden_model_1.n2136 ;
  wire [7:0] \oc8051_golden_model_1.n2137 ;
  wire \oc8051_golden_model_1.n2141 ;
  wire [6:0] \oc8051_golden_model_1.n2142 ;
  wire [7:0] \oc8051_golden_model_1.n2143 ;
  wire [6:0] \oc8051_golden_model_1.n2144 ;
  wire [7:0] \oc8051_golden_model_1.n2145 ;
  wire \oc8051_golden_model_1.n2160 ;
  wire [7:0] \oc8051_golden_model_1.n2161 ;
  wire [7:0] \oc8051_golden_model_1.n2201 ;
  wire [6:0] \oc8051_golden_model_1.n2202 ;
  wire [7:0] \oc8051_golden_model_1.n2203 ;
  wire [3:0] \oc8051_golden_model_1.n2210 ;
  wire \oc8051_golden_model_1.n2211 ;
  wire [7:0] \oc8051_golden_model_1.n2212 ;
  wire [6:0] \oc8051_golden_model_1.n2213 ;
  wire \oc8051_golden_model_1.n2228 ;
  wire [7:0] \oc8051_golden_model_1.n2229 ;
  wire [7:0] \oc8051_golden_model_1.n2441 ;
  wire [7:0] \oc8051_golden_model_1.n2453 ;
  wire [6:0] \oc8051_golden_model_1.n2454 ;
  wire \oc8051_golden_model_1.n2469 ;
  wire [7:0] \oc8051_golden_model_1.n2470 ;
  wire \oc8051_golden_model_1.n2474 ;
  wire \oc8051_golden_model_1.n2476 ;
  wire \oc8051_golden_model_1.n2482 ;
  wire [7:0] \oc8051_golden_model_1.n2483 ;
  wire [6:0] \oc8051_golden_model_1.n2484 ;
  wire \oc8051_golden_model_1.n2499 ;
  wire [7:0] \oc8051_golden_model_1.n2500 ;
  wire \oc8051_golden_model_1.n2504 ;
  wire \oc8051_golden_model_1.n2506 ;
  wire \oc8051_golden_model_1.n2512 ;
  wire [7:0] \oc8051_golden_model_1.n2513 ;
  wire [6:0] \oc8051_golden_model_1.n2514 ;
  wire \oc8051_golden_model_1.n2529 ;
  wire [7:0] \oc8051_golden_model_1.n2530 ;
  wire \oc8051_golden_model_1.n2534 ;
  wire \oc8051_golden_model_1.n2536 ;
  wire \oc8051_golden_model_1.n2542 ;
  wire [7:0] \oc8051_golden_model_1.n2543 ;
  wire [6:0] \oc8051_golden_model_1.n2544 ;
  wire \oc8051_golden_model_1.n2559 ;
  wire [7:0] \oc8051_golden_model_1.n2560 ;
  wire \oc8051_golden_model_1.n2562 ;
  wire [7:0] \oc8051_golden_model_1.n2563 ;
  wire [6:0] \oc8051_golden_model_1.n2564 ;
  wire [7:0] \oc8051_golden_model_1.n2565 ;
  wire [7:0] \oc8051_golden_model_1.n2566 ;
  wire [6:0] \oc8051_golden_model_1.n2567 ;
  wire [7:0] \oc8051_golden_model_1.n2568 ;
  wire [15:0] \oc8051_golden_model_1.n2572 ;
  wire \oc8051_golden_model_1.n2578 ;
  wire [7:0] \oc8051_golden_model_1.n2579 ;
  wire [6:0] \oc8051_golden_model_1.n2580 ;
  wire \oc8051_golden_model_1.n2595 ;
  wire [7:0] \oc8051_golden_model_1.n2596 ;
  wire \oc8051_golden_model_1.n2599 ;
  wire [7:0] \oc8051_golden_model_1.n2600 ;
  wire [6:0] \oc8051_golden_model_1.n2601 ;
  wire [7:0] \oc8051_golden_model_1.n2602 ;
  wire \oc8051_golden_model_1.n2634 ;
  wire [7:0] \oc8051_golden_model_1.n2635 ;
  wire [6:0] \oc8051_golden_model_1.n2636 ;
  wire [7:0] \oc8051_golden_model_1.n2637 ;
  wire [7:0] \oc8051_golden_model_1.n2643 ;
  wire [6:0] \oc8051_golden_model_1.n2644 ;
  wire [7:0] \oc8051_golden_model_1.n2645 ;
  wire [7:0] \oc8051_golden_model_1.n2651 ;
  wire [6:0] \oc8051_golden_model_1.n2652 ;
  wire [7:0] \oc8051_golden_model_1.n2653 ;
  wire \oc8051_golden_model_1.n2658 ;
  wire [7:0] \oc8051_golden_model_1.n2659 ;
  wire [6:0] \oc8051_golden_model_1.n2660 ;
  wire [7:0] \oc8051_golden_model_1.n2661 ;
  wire \oc8051_golden_model_1.n2666 ;
  wire [7:0] \oc8051_golden_model_1.n2667 ;
  wire [6:0] \oc8051_golden_model_1.n2668 ;
  wire [7:0] \oc8051_golden_model_1.n2669 ;
  wire [7:0] \oc8051_golden_model_1.n2694 ;
  wire [6:0] \oc8051_golden_model_1.n2695 ;
  wire [7:0] \oc8051_golden_model_1.n2696 ;
  wire [3:0] \oc8051_golden_model_1.n2697 ;
  wire [7:0] \oc8051_golden_model_1.n2698 ;
  wire \oc8051_golden_model_1.n2699 ;
  wire \oc8051_golden_model_1.n2700 ;
  wire \oc8051_golden_model_1.n2701 ;
  wire \oc8051_golden_model_1.n2702 ;
  wire \oc8051_golden_model_1.n2703 ;
  wire \oc8051_golden_model_1.n2704 ;
  wire \oc8051_golden_model_1.n2705 ;
  wire \oc8051_golden_model_1.n2706 ;
  wire \oc8051_golden_model_1.n2713 ;
  wire [7:0] \oc8051_golden_model_1.n2714 ;
  wire \oc8051_golden_model_1.n2752 ;
  wire \oc8051_golden_model_1.n2753 ;
  wire \oc8051_golden_model_1.n2754 ;
  wire \oc8051_golden_model_1.n2755 ;
  wire \oc8051_golden_model_1.n2756 ;
  wire \oc8051_golden_model_1.n2757 ;
  wire \oc8051_golden_model_1.n2758 ;
  wire \oc8051_golden_model_1.n2759 ;
  wire \oc8051_golden_model_1.n2766 ;
  wire [7:0] \oc8051_golden_model_1.n2767 ;
  wire \oc8051_golden_model_1.n2768 ;
  wire \oc8051_golden_model_1.n2769 ;
  wire \oc8051_golden_model_1.n2770 ;
  wire \oc8051_golden_model_1.n2771 ;
  wire \oc8051_golden_model_1.n2772 ;
  wire \oc8051_golden_model_1.n2773 ;
  wire \oc8051_golden_model_1.n2774 ;
  wire \oc8051_golden_model_1.n2775 ;
  wire \oc8051_golden_model_1.n2782 ;
  wire [7:0] \oc8051_golden_model_1.n2783 ;
  wire [7:0] \oc8051_golden_model_1.n2815 ;
  wire [6:0] \oc8051_golden_model_1.n2816 ;
  wire [7:0] \oc8051_golden_model_1.n2817 ;
  wire \oc8051_golden_model_1.n2836 ;
  wire [7:0] \oc8051_golden_model_1.n2837 ;
  wire [6:0] \oc8051_golden_model_1.n2838 ;
  wire [7:0] \oc8051_golden_model_1.n2854 ;
  wire [7:0] \oc8051_golden_model_1.n2858 ;
  wire [3:0] \oc8051_golden_model_1.n2859 ;
  wire [7:0] \oc8051_golden_model_1.n2860 ;
  wire \oc8051_golden_model_1.n2861 ;
  wire \oc8051_golden_model_1.n2862 ;
  wire \oc8051_golden_model_1.n2863 ;
  wire \oc8051_golden_model_1.n2864 ;
  wire \oc8051_golden_model_1.n2865 ;
  wire \oc8051_golden_model_1.n2866 ;
  wire \oc8051_golden_model_1.n2867 ;
  wire \oc8051_golden_model_1.n2868 ;
  wire [7:0] \oc8051_golden_model_1.n2876 ;
  wire \oc8051_golden_model_1.n2894 ;
  wire [7:0] \oc8051_golden_model_1.n2895 ;
  wire [7:0] \oc8051_golden_model_1.n2896 ;
  wire \oc8051_golden_model_1.n2912 ;
  wire [7:0] \oc8051_golden_model_1.n2913 ;
  wire \oc8051_golden_model_1.rst ;
  wire [34:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.des1 ;
  wire [7:0] \oc8051_top_1.des2 ;
  wire \oc8051_top_1.desAc ;
  wire \oc8051_top_1.desCy ;
  wire \oc8051_top_1.desOv ;
  wire [7:0] \oc8051_top_1.des_acc ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire [7:0] \oc8051_top_1.ie ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.des ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.data_in ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.alu ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des1 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des2 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des_acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.wr_dat ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_data_in ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat2 ;
  wire \oc8051_top_1.oc8051_sfr1.desAc ;
  wire \oc8051_top_1.oc8051_sfr1.desOv ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.des_acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.cy_in ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire [7:0] \oc8051_top_1.sub_result ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire [7:0] \oc8051_top_1.wr_dat ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  wire p12_equal;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire p1_valid_r;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_pc;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  wire regs_always_zero;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_25964_, rst);
  not (_15509_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_15520_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15540_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _15520_);
  and (_15541_, _15540_, _15509_);
  and (_15552_, \oc8051_top_1.oc8051_decoder1.wr , _15520_);
  not (_15563_, _15552_);
  nor (_15574_, _15563_, _15541_);
  and (_15585_, _15574_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_15596_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_15607_, _15596_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_15617_, _15607_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_15628_, _15617_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_15639_, _15628_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_15650_, _15639_);
  and (_15661_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _15520_);
  and (_15672_, _15661_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_15683_, _15672_, _15509_);
  not (_15694_, _15683_);
  nor (_15704_, _15628_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_15715_, _15704_, _15694_);
  and (_15726_, _15715_, _15650_);
  not (_15737_, _15726_);
  and (_15748_, _15672_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_15759_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_15770_, _15661_, _15759_);
  and (_15781_, _15770_, _15509_);
  and (_15791_, _15781_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_15802_, _15791_, _15748_);
  not (_15813_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_15824_, _15541_, _15813_);
  and (_15835_, _15824_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_15846_, _15770_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_15857_, _15846_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_15868_, _15857_, _15835_);
  and (_15878_, _15868_, _15802_);
  and (_15889_, _15878_, _15737_);
  and (_15900_, _15639_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_15911_, _15900_);
  nor (_15922_, _15639_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_15933_, _15922_, _15694_);
  and (_15944_, _15933_, _15911_);
  not (_15955_, _15944_);
  and (_15965_, _15781_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_15976_, _15965_, _15748_);
  and (_15987_, _15824_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_15998_, _15846_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_16009_, _15998_, _15987_);
  and (_16020_, _16009_, _15976_);
  and (_16031_, _16020_, _15955_);
  nor (_16042_, _16031_, _15889_);
  not (_16052_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_16063_, _15900_, _16052_);
  and (_16074_, _15900_, _16052_);
  nor (_16085_, _16074_, _16063_);
  nor (_16096_, _16085_, _15694_);
  not (_16107_, _16096_);
  and (_16118_, _15824_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_16129_, _16118_);
  not (_16139_, _15748_);
  and (_16150_, _15781_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_16171_, _15846_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_16172_, _16171_, _16150_);
  and (_16183_, _16172_, _16139_);
  and (_16194_, _16183_, _16129_);
  and (_16205_, _16194_, _16107_);
  not (_16216_, _16205_);
  and (_16226_, _15846_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_16237_, _15781_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_16248_, _16237_, _16226_);
  not (_16259_, _15617_);
  nor (_16270_, _15607_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_16281_, _16270_, _15694_);
  and (_16292_, _16281_, _16259_);
  or (_16303_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_16313_, _16303_, _15520_);
  nor (_16324_, _16313_, _15661_);
  and (_16335_, _16324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_16346_, _15824_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_16357_, _16346_, _16335_);
  not (_16368_, _16357_);
  nor (_16379_, _16368_, _16292_);
  and (_16390_, _16379_, _16248_);
  not (_16400_, _16390_);
  and (_16411_, _15824_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_16422_, _16411_, _15748_);
  and (_16433_, _15846_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_16444_, _16433_);
  and (_16455_, _16444_, _16422_);
  nor (_16466_, _15617_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_16477_, _16466_);
  nor (_16497_, _15694_, _15628_);
  and (_16498_, _16497_, _16477_);
  and (_16509_, _15781_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and (_16520_, _16324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor (_16531_, _16520_, _16509_);
  not (_16542_, _16531_);
  nor (_16553_, _16542_, _16498_);
  and (_16564_, _16553_, _16455_);
  nor (_16574_, _16564_, _16400_);
  and (_16585_, _16574_, _16216_);
  and (_16596_, _16585_, _16042_);
  nor (_16607_, _15596_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_16618_, _16607_, _15607_);
  and (_16629_, _16618_, _15683_);
  and (_16640_, _15824_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_16651_, _16640_, _16629_);
  and (_16661_, _15846_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_16672_, _15781_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and (_16683_, _16324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_16694_, _16683_, _16672_);
  nor (_16705_, _16694_, _16661_);
  and (_16716_, _16705_, _16651_);
  not (_16727_, _16716_);
  not (_16738_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_16748_, _15683_, _16738_);
  and (_16759_, _15781_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_16770_, _16759_, _16748_);
  and (_16781_, _16324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  not (_16792_, _16781_);
  and (_16803_, _15846_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_16814_, _15824_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_16825_, _16814_, _16803_);
  and (_16835_, _16825_, _16792_);
  and (_16846_, _16835_, _16770_);
  nor (_16867_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_16868_, _16867_, _15596_);
  and (_16879_, _16868_, _15683_);
  and (_16890_, _15824_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_16901_, _16890_, _16879_);
  and (_16912_, _15846_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_16922_, _15781_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_16933_, _16324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_16944_, _16933_, _16922_);
  nor (_16955_, _16944_, _16912_);
  and (_16966_, _16955_, _16901_);
  nor (_16977_, _16966_, _16846_);
  and (_16988_, _16977_, _16727_);
  and (_16999_, _16988_, _16596_);
  or (_17009_, _16999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  not (_17020_, ABINPUT[0]);
  nand (_17031_, _16999_, _17020_);
  and (_17042_, _17031_, _17009_);
  and (_17053_, _17042_, _15585_);
  not (_17064_, _15574_);
  and (_17075_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  not (_17086_, ABINPUT[26]);
  and (_17096_, _16966_, _16846_);
  and (_17107_, _17096_, _16716_);
  and (_17118_, _17107_, _16596_);
  nand (_17129_, _17118_, _17086_);
  not (_17140_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_17151_, _15574_, _17140_);
  or (_17162_, _17118_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_17172_, _17162_, _17151_);
  and (_17183_, _17172_, _17129_);
  or (_17194_, _17183_, _17075_);
  or (_17205_, _17194_, _17053_);
  and (_05323_, _17205_, _25964_);
  not (_17226_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor (_17237_, _17118_, _17226_);
  and (_17248_, _17107_, ABINPUT[0]);
  and (_17258_, _17248_, _16596_);
  or (_17269_, _17258_, _17237_);
  and (_17280_, _17269_, _15585_);
  nor (_17291_, _15574_, _17226_);
  and (_17302_, _17118_, ABINPUT[19]);
  or (_17313_, _17302_, _17237_);
  and (_17324_, _17313_, _17151_);
  or (_17335_, _17324_, _17291_);
  or (_17345_, _17335_, _17280_);
  and (_23586_, _17345_, _25964_);
  not (_17366_, _16846_);
  and (_17377_, _16966_, _17366_);
  and (_17388_, _17377_, _16716_);
  nand (_17399_, _17388_, _16596_);
  and (_17410_, _17399_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_17421_, _17388_, ABINPUT[0]);
  and (_17431_, _17421_, _16596_);
  or (_17442_, _17431_, _17410_);
  and (_17453_, _17442_, _15585_);
  and (_17464_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  not (_17475_, ABINPUT[20]);
  nand (_17486_, _17118_, _17475_);
  or (_17497_, _17118_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_17508_, _17497_, _17151_);
  and (_17518_, _17508_, _17486_);
  or (_17529_, _17518_, _17464_);
  or (_17540_, _17529_, _17453_);
  and (_23596_, _17540_, _25964_);
  not (_17561_, _16966_);
  and (_17572_, _17561_, _16846_);
  and (_17583_, _17572_, _16716_);
  nand (_17594_, _17583_, _16596_);
  and (_17604_, _17594_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_17625_, _17583_, ABINPUT[0]);
  and (_17626_, _17625_, _16596_);
  or (_17637_, _17626_, _17604_);
  and (_17648_, _17637_, _15585_);
  and (_17659_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_17670_, ABINPUT[21]);
  nand (_17681_, _17118_, _17670_);
  or (_17692_, _17118_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_17703_, _17692_, _17151_);
  and (_17714_, _17703_, _17681_);
  or (_17725_, _17714_, _17659_);
  or (_17736_, _17725_, _17648_);
  and (_23606_, _17736_, _25964_);
  and (_17757_, _16977_, _16716_);
  nand (_17768_, _17757_, _16596_);
  and (_17779_, _17768_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_17790_, _17757_, ABINPUT[0]);
  and (_17801_, _17790_, _16596_);
  or (_17812_, _17801_, _17779_);
  and (_17823_, _17812_, _15585_);
  and (_17834_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not (_17845_, ABINPUT[22]);
  nand (_17856_, _17118_, _17845_);
  or (_17867_, _17118_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_17877_, _17867_, _17151_);
  and (_17888_, _17877_, _17856_);
  or (_17899_, _17888_, _17834_);
  or (_17910_, _17899_, _17823_);
  and (_23617_, _17910_, _25964_);
  and (_17931_, _17096_, _16727_);
  nand (_17942_, _17931_, _16596_);
  and (_17953_, _17942_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_17964_, _17931_, ABINPUT[0]);
  and (_17975_, _17964_, _16596_);
  or (_17986_, _17975_, _17953_);
  and (_17997_, _17986_, _15585_);
  and (_18008_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_18019_, ABINPUT[23]);
  nand (_18030_, _17118_, _18019_);
  or (_18051_, _17118_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_18052_, _18051_, _17151_);
  and (_18063_, _18052_, _18030_);
  or (_18074_, _18063_, _18008_);
  or (_18095_, _18074_, _17997_);
  and (_23627_, _18095_, _25964_);
  and (_18106_, _17377_, _16727_);
  nand (_18117_, _18106_, _16596_);
  and (_18128_, _18117_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_18139_, _18106_, ABINPUT[0]);
  and (_18150_, _18139_, _16596_);
  or (_18161_, _18150_, _18128_);
  and (_18172_, _18161_, _15585_);
  and (_18183_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_18194_, ABINPUT[24]);
  nand (_18205_, _17118_, _18194_);
  or (_18216_, _17118_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_18227_, _18216_, _17151_);
  and (_18238_, _18227_, _18205_);
  or (_18249_, _18238_, _18183_);
  or (_18260_, _18249_, _18172_);
  and (_23637_, _18260_, _25964_);
  and (_18281_, _17572_, _16727_);
  nand (_18292_, _18281_, _16596_);
  and (_18302_, _18292_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_18313_, _18281_, ABINPUT[0]);
  and (_18324_, _18313_, _16596_);
  or (_18335_, _18324_, _18302_);
  and (_18346_, _18335_, _15585_);
  and (_18357_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  not (_18368_, ABINPUT[25]);
  nand (_18379_, _17118_, _18368_);
  or (_18390_, _17118_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_18401_, _18390_, _17151_);
  and (_18412_, _18401_, _18379_);
  or (_18423_, _18412_, _18357_);
  or (_18434_, _18423_, _18346_);
  and (_23647_, _18434_, _25964_);
  and (_18455_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_18466_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_18477_, _18466_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_18488_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_18499_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_18510_, _18499_, _18488_);
  and (_18521_, _18466_, _15520_);
  and (_18532_, _18521_, _18510_);
  and (_18543_, _18510_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_18554_, _18543_, _18532_);
  and (_18565_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_18576_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_18587_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_18598_, _18587_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_18609_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  not (_18620_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not (_18631_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_18642_, _18631_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_18653_, _18642_, _18620_);
  and (_18664_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_18675_, _18664_, _18609_);
  and (_18685_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_18696_, _18685_, _18620_);
  and (_18707_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  not (_18718_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_18729_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _18718_);
  and (_18740_, _18729_, _18620_);
  and (_18751_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_18762_, _18751_, _18707_);
  and (_18773_, _18762_, _18675_);
  nor (_18784_, _18587_, _18620_);
  and (_18795_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_18806_, _18587_, _18620_);
  and (_18817_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_18828_, _18817_, _18795_);
  and (_18839_, _18828_, _18773_);
  and (_18850_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_18861_, _18850_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_18872_, _18861_, _18839_);
  nor (_18883_, _18872_, _18576_);
  nor (_18894_, _18883_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_18905_, _18894_, _18565_);
  and (_18916_, _18905_, _18532_);
  nor (_18927_, _18916_, _18554_);
  and (_18938_, _18510_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_18949_, _18938_, _18532_);
  and (_18960_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_18971_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_18992_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_18993_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_19004_, _18993_, _18992_);
  and (_19015_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_19026_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_19037_, _19026_, _19015_);
  and (_19047_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_19058_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_19069_, _19058_, _19047_);
  and (_19080_, _19069_, _19037_);
  and (_19091_, _19080_, _19004_);
  nor (_19102_, _19091_, _18861_);
  nor (_19113_, _19102_, _18971_);
  nor (_19124_, _19113_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_19135_, _19124_, _18960_);
  and (_19146_, _19135_, _18532_);
  nor (_19157_, _19146_, _18949_);
  not (_19168_, _19157_);
  nor (_19179_, _19168_, _18927_);
  and (_19190_, _18510_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_19201_, _19190_, _18532_);
  not (_19212_, _18532_);
  not (_19223_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_19234_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_19245_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_19256_, _19245_, _19234_);
  and (_19267_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_19278_, _18850_, _19267_);
  and (_19289_, _19278_, _19256_);
  and (_19300_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not (_19311_, _19300_);
  and (_19322_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_19333_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_19344_, _19333_, _19322_);
  and (_19355_, _19344_, _19311_);
  and (_19366_, _19355_, _19289_);
  and (_19377_, _19366_, _19223_);
  nor (_19388_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _19223_);
  nor (_19399_, _19388_, _19377_);
  nor (_19409_, _19399_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_19420_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_19431_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _19420_);
  nor (_19442_, _19431_, _19409_);
  nor (_19453_, _19442_, _19212_);
  nor (_19464_, _19453_, _19201_);
  not (_19475_, _19464_);
  and (_19497_, _18510_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_19498_, _19497_, _18532_);
  and (_19520_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_19521_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_19543_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_19544_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_19566_, _19544_, _19543_);
  and (_19567_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_19578_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_19589_, _19578_, _19567_);
  and (_19600_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_19611_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_19622_, _19611_, _19600_);
  and (_19633_, _19622_, _19589_);
  and (_19644_, _19633_, _19566_);
  nor (_19655_, _19644_, _18850_);
  and (_19666_, _19655_, _19223_);
  nor (_19677_, _19666_, _19521_);
  nor (_19688_, _19677_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_19699_, _19688_, _19520_);
  and (_19710_, _19699_, _18532_);
  nor (_19721_, _19710_, _19498_);
  and (_19732_, _19721_, _19475_);
  and (_19743_, _19732_, _19179_);
  and (_19754_, _18510_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_19765_, _19754_, _18532_);
  and (_19775_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_19786_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_19797_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_19808_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_19819_, _19808_, _19797_);
  and (_19830_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_19841_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_19852_, _19841_, _19830_);
  and (_19863_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_19874_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_19885_, _19874_, _19863_);
  and (_19896_, _19885_, _19852_);
  and (_19907_, _19896_, _19819_);
  nor (_19918_, _19907_, _18850_);
  and (_19929_, _19918_, _19223_);
  or (_19940_, _19929_, _19786_);
  and (_19951_, _19940_, _19420_);
  nor (_19962_, _19951_, _19775_);
  and (_19973_, _19962_, _18532_);
  nor (_19984_, _19973_, _19765_);
  and (_19995_, _18510_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_20006_, _19995_, _18532_);
  and (_20017_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  not (_20028_, _20017_);
  and (_20039_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_20050_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_20061_, _20050_, _20039_);
  and (_20072_, _20061_, _20028_);
  and (_20083_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_20094_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_20105_, _20094_, _20083_);
  and (_20116_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_20127_, _20116_, _18850_);
  and (_20137_, _20127_, _20105_);
  and (_20148_, _20137_, _20072_);
  and (_20159_, _20148_, _19223_);
  nor (_20170_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _19223_);
  nor (_20181_, _20170_, _20159_);
  nor (_20192_, _20181_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_20203_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _19420_);
  nor (_20214_, _20203_, _20192_);
  nor (_20225_, _20214_, _19212_);
  nor (_20236_, _20225_, _20006_);
  and (_20247_, _18510_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_20258_, _20247_, _18532_);
  and (_20269_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_20280_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_20291_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_20302_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_20313_, _20302_, _20291_);
  and (_20324_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_20335_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_20346_, _20335_, _20324_);
  and (_20357_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_20368_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_20379_, _20368_, _20357_);
  and (_20390_, _20379_, _20346_);
  and (_20401_, _20390_, _20313_);
  nor (_20412_, _20401_, _18861_);
  nor (_20423_, _20412_, _20280_);
  nor (_20434_, _20423_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_20445_, _20434_, _20269_);
  and (_20456_, _20445_, _18532_);
  nor (_20467_, _20456_, _20258_);
  and (_20478_, _18510_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_20489_, _20478_, _18532_);
  and (_20500_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_20510_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_20521_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_20532_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_20543_, _20532_, _20521_);
  and (_20554_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_20565_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_20576_, _20565_, _20554_);
  and (_20587_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_20598_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_20609_, _20598_, _20587_);
  and (_20620_, _20609_, _20576_);
  and (_20631_, _20620_, _20543_);
  nor (_20642_, _20631_, _18850_);
  and (_20653_, _20642_, _19223_);
  or (_20664_, _20653_, _20510_);
  and (_20675_, _20664_, _19420_);
  nor (_20686_, _20675_, _20500_);
  and (_20697_, _20686_, _18532_);
  nor (_20708_, _20697_, _20489_);
  nor (_20719_, _20708_, _20467_);
  and (_20730_, _20719_, _20236_);
  and (_20741_, _20730_, _19984_);
  and (_20752_, _20741_, _19743_);
  not (_20763_, _20752_);
  not (_20774_, _19721_);
  and (_20785_, _20774_, _19179_);
  and (_20796_, _20785_, _19464_);
  and (_20807_, _20741_, _20796_);
  and (_20818_, _19721_, _18927_);
  and (_20829_, _20818_, _19168_);
  and (_20840_, _20829_, _19464_);
  and (_20850_, _20741_, _20840_);
  nor (_20861_, _20850_, _20807_);
  and (_20872_, _20861_, _20763_);
  nor (_20883_, _20872_, _18477_);
  not (_20894_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_20905_, \oc8051_top_1.oc8051_decoder1.state [1], _15520_);
  and (_20916_, _20905_, _20894_);
  and (_20927_, _19168_, _18927_);
  nor (_20938_, _20236_, _19984_);
  and (_20949_, _20938_, _20719_);
  and (_20960_, _20949_, _20927_);
  and (_20971_, _20960_, _20916_);
  not (_20982_, _20971_);
  and (_20993_, _20785_, _19475_);
  not (_21004_, _20708_);
  and (_21015_, _21004_, _20467_);
  and (_21026_, _20938_, _21015_);
  and (_21037_, _21026_, _20993_);
  and (_21048_, _21026_, _19743_);
  nor (_21059_, _21048_, _21037_);
  and (_21070_, _21059_, _20982_);
  not (_21081_, _21070_);
  nor (_21092_, _21081_, _20883_);
  nor (_21103_, _21092_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_21114_, _21103_, _18455_);
  and (_21125_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_21136_, _19984_);
  and (_21147_, _20730_, _21136_);
  and (_21158_, _21147_, _20993_);
  and (_21169_, _20774_, _18927_);
  and (_21180_, _21169_, _19168_);
  and (_21190_, _21180_, _19464_);
  and (_21201_, _21190_, _20730_);
  nor (_21212_, _21201_, _21158_);
  and (_21223_, _20796_, _21147_);
  not (_21234_, _20236_);
  and (_21245_, _21234_, _19984_);
  and (_21256_, _21245_, _21015_);
  and (_21267_, _21256_, _20993_);
  nor (_21278_, _21267_, _21223_);
  and (_21289_, _21278_, _21212_);
  and (_21300_, _19157_, _18927_);
  and (_21311_, _21300_, _20774_);
  and (_21322_, _21311_, _19464_);
  and (_21333_, _21322_, _21147_);
  and (_21344_, _19743_, _21147_);
  nor (_21355_, _21344_, _21333_);
  nor (_21366_, _19157_, _18927_);
  and (_21377_, _21366_, _19721_);
  and (_21388_, _21377_, _20949_);
  and (_21399_, _21388_, _19475_);
  and (_21410_, _19721_, _19464_);
  and (_21421_, _21410_, _21366_);
  and (_21432_, _21366_, _20774_);
  and (_21443_, _21432_, _19464_);
  or (_21454_, _21443_, _21421_);
  and (_21465_, _21454_, _20949_);
  nor (_21476_, _21465_, _21399_);
  and (_21487_, _21476_, _21355_);
  and (_21498_, _21487_, _21289_);
  and (_21508_, _19721_, _19179_);
  and (_21519_, _20467_, _20236_);
  and (_21530_, _21519_, _21004_);
  and (_21541_, _21530_, _19475_);
  and (_21552_, _21541_, _21508_);
  not (_21563_, _21552_);
  and (_21574_, _21377_, _21147_);
  and (_21585_, _20708_, _19475_);
  and (_21596_, _21585_, _21508_);
  nor (_21607_, _21596_, _21574_);
  and (_21618_, _21607_, _21563_);
  and (_21629_, _21311_, _19475_);
  and (_21640_, _21629_, _21256_);
  and (_21651_, _20829_, _19475_);
  and (_21662_, _21651_, _21256_);
  nor (_21673_, _21662_, _21640_);
  and (_21684_, _20949_, _21311_);
  and (_21695_, _21651_, _20730_);
  nor (_21706_, _21695_, _21684_);
  and (_21717_, _21706_, _21673_);
  and (_21728_, _21717_, _21618_);
  and (_21739_, _21728_, _21498_);
  and (_21750_, _21180_, _19475_);
  and (_21761_, _21750_, _20730_);
  and (_21772_, _21443_, _21256_);
  and (_21783_, _21410_, _19179_);
  and (_21794_, _21783_, _20949_);
  or (_21805_, _21794_, _21772_);
  nor (_21816_, _21805_, _21761_);
  and (_21827_, _20840_, _21147_);
  and (_21837_, _21322_, _21256_);
  nor (_21848_, _21837_, _21827_);
  and (_21859_, _21848_, _21816_);
  and (_21870_, _20949_, _19743_);
  and (_21881_, _21750_, _21256_);
  nor (_21892_, _21881_, _21870_);
  and (_21903_, _21783_, _21147_);
  and (_21914_, _21629_, _21147_);
  nor (_21925_, _21914_, _21903_);
  and (_21936_, _21925_, _21892_);
  and (_21947_, _21936_, _21859_);
  nor (_21958_, _21377_, _21190_);
  and (_21969_, _19732_, _21300_);
  and (_21980_, _21432_, _19475_);
  and (_21991_, _19179_, _19464_);
  or (_22002_, _21991_, _21980_);
  nor (_22013_, _22002_, _21969_);
  nand (_22024_, _22013_, _21958_);
  and (_22035_, _22024_, _21256_);
  not (_22046_, _22035_);
  and (_22057_, _22046_, _21947_);
  and (_22068_, _22057_, _21739_);
  nor (_22079_, _22068_, _18477_);
  and (_22090_, _21443_, _20949_);
  or (_22101_, _22090_, _21399_);
  and (_22112_, _22101_, _20916_);
  and (_22123_, _21574_, _20905_);
  and (_22134_, _22123_, \oc8051_top_1.oc8051_decoder1.state [0]);
  or (_22145_, _22134_, _20971_);
  or (_22155_, _22145_, _22112_);
  nor (_22166_, _22155_, _22079_);
  nor (_22177_, _22166_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_22188_, _22177_, _21125_);
  and (_22199_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_22210_, _21004_, _19464_);
  and (_22221_, _22210_, _21519_);
  and (_22232_, _22221_, _21180_);
  and (_22243_, _21530_, _21377_);
  or (_22254_, _22243_, _22232_);
  not (_22265_, _22254_);
  and (_22276_, _20949_, _21322_);
  and (_22287_, _21530_, _20993_);
  nor (_22298_, _22287_, _22276_);
  and (_22309_, _21530_, _21432_);
  and (_22320_, _21783_, _21530_);
  nor (_22331_, _22320_, _22309_);
  not (_22342_, _22331_);
  and (_22353_, _21651_, _21530_);
  nor (_22364_, _22353_, _22342_);
  and (_22375_, _22364_, _22298_);
  and (_22386_, _22375_, _22265_);
  and (_22397_, _21530_, _21311_);
  and (_22408_, _21530_, _20796_);
  nor (_22419_, _22408_, _22397_);
  and (_22430_, _20818_, _19157_);
  or (_22441_, _22430_, _21180_);
  and (_22451_, _22441_, _21541_);
  nor (_22462_, _22451_, _21574_);
  and (_22473_, _22462_, _22419_);
  and (_22484_, _22473_, _20872_);
  and (_22495_, _22484_, _22386_);
  nor (_22506_, _22495_, _18477_);
  and (_22517_, _20916_, _20949_);
  and (_22528_, _22517_, _20829_);
  or (_22539_, _22528_, _22134_);
  nor (_22550_, _22539_, _22506_);
  nor (_22561_, _22550_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_22572_, _22561_, _22199_);
  nor (_22583_, _22572_, _22188_);
  and (_22594_, _22583_, _21114_);
  and (_24117_, _22594_, _25964_);
  not (_22615_, _17151_);
  not (_22626_, _16031_);
  nor (_22637_, _16205_, _22626_);
  and (_22648_, _16564_, _15889_);
  and (_22659_, _22648_, _22637_);
  and (_22670_, _22659_, _16390_);
  nand (_22681_, _22670_, _17388_);
  nor (_22692_, _22681_, _22615_);
  and (_22703_, _22692_, ABINPUT[10]);
  nor (_22714_, _22692_, _16052_);
  nor (_22725_, _22714_, _22703_);
  not (_22736_, _22725_);
  not (_22747_, _22692_);
  and (_22758_, _22747_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_22767_, _22692_, ABINPUT[9]);
  nor (_22774_, _22767_, _22758_);
  and (_22782_, _22747_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_22790_, _22692_, ABINPUT[8]);
  nor (_22797_, _22790_, _22782_);
  and (_22805_, _22747_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_22813_, _22692_, ABINPUT[7]);
  nor (_22820_, _22813_, _22805_);
  and (_22827_, _22747_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_22828_, _22692_, ABINPUT[6]);
  nor (_22829_, _22828_, _22827_);
  and (_22831_, _22747_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_22842_, _22692_, ABINPUT[5]);
  nor (_22853_, _22842_, _22831_);
  and (_22864_, _22747_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_22875_, _22692_, ABINPUT[4]);
  nor (_22886_, _22875_, _22864_);
  nor (_22897_, _22692_, _16738_);
  and (_22907_, _22692_, ABINPUT[3]);
  nor (_22918_, _22907_, _22897_);
  and (_22929_, _22918_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_22940_, _22929_, _22886_);
  and (_22951_, _22940_, _22853_);
  and (_22962_, _22951_, _22829_);
  and (_22973_, _22962_, _22820_);
  and (_22984_, _22973_, _22797_);
  and (_22995_, _22984_, _22774_);
  and (_23006_, _22995_, _22736_);
  nor (_23017_, _22995_, _22736_);
  nor (_23028_, _23017_, _23006_);
  and (_23039_, _23028_, _15694_);
  nor (_23050_, _23039_, _16096_);
  nor (_23061_, _23050_, _22692_);
  nor (_23072_, _23061_, _22703_);
  nor (_24137_, _23072_, rst);
  not (_23093_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_23097_, _22918_, _23093_);
  nor (_23098_, _22918_, _23093_);
  nor (_23099_, _23098_, _23097_);
  and (_23100_, _23099_, _15694_);
  nor (_23101_, _23100_, _16748_);
  nor (_23102_, _23101_, _22692_);
  nor (_23103_, _23102_, _22907_);
  nand (_25125_, _23103_, _25964_);
  nor (_23104_, _22929_, _22886_);
  nor (_23105_, _23104_, _22940_);
  nor (_23106_, _23105_, _15683_);
  nor (_23107_, _23106_, _16879_);
  nor (_23108_, _23107_, _22692_);
  nor (_23109_, _23108_, _22875_);
  nand (_25133_, _23109_, _25964_);
  nor (_23110_, _22940_, _22853_);
  nor (_23111_, _23110_, _22951_);
  nor (_23112_, _23111_, _15683_);
  nor (_23113_, _23112_, _16629_);
  nor (_23114_, _23113_, _22692_);
  nor (_23115_, _23114_, _22842_);
  nand (_25141_, _23115_, _25964_);
  nor (_23116_, _22951_, _22829_);
  nor (_23117_, _23116_, _22962_);
  nor (_23118_, _23117_, _15683_);
  nor (_23119_, _23118_, _16292_);
  nor (_23120_, _23119_, _22692_);
  nor (_23121_, _23120_, _22828_);
  nor (_25149_, _23121_, rst);
  nor (_23122_, _22962_, _22820_);
  nor (_23123_, _23122_, _22973_);
  nor (_23124_, _23123_, _15683_);
  nor (_23125_, _23124_, _16498_);
  nor (_23126_, _23125_, _22692_);
  nor (_23127_, _23126_, _22813_);
  nor (_25156_, _23127_, rst);
  nor (_23128_, _22973_, _22797_);
  nor (_23129_, _23128_, _22984_);
  nor (_23130_, _23129_, _15683_);
  nor (_23131_, _23130_, _15726_);
  nor (_23132_, _23131_, _22692_);
  nor (_23133_, _23132_, _22790_);
  nor (_25164_, _23133_, rst);
  nor (_23134_, _22984_, _22774_);
  nor (_23135_, _23134_, _22995_);
  nor (_23136_, _23135_, _15683_);
  nor (_23137_, _23136_, _15944_);
  nor (_23138_, _23137_, _22692_);
  nor (_23139_, _23138_, _22767_);
  nor (_25175_, _23139_, rst);
  and (_23140_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _15520_);
  and (_23141_, _23140_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_23142_, _17757_, _16390_);
  nand (_23143_, _23142_, _22659_);
  nor (_23144_, _23143_, _22615_);
  or (_23145_, _23144_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nand (_23146_, _23144_, _17086_);
  and (_23147_, _23146_, _23145_);
  or (_23148_, _23147_, _23141_);
  not (_23149_, ABINPUT[18]);
  nand (_23150_, _23141_, _23149_);
  and (_23151_, _23150_, _25964_);
  and (_27135_, _23151_, _23148_);
  and (_23152_, _22670_, _17583_);
  and (_23153_, _23152_, _17151_);
  nor (_23154_, _23153_, _23141_);
  and (_23155_, _23154_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nor (_23156_, _23154_, _17086_);
  or (_23157_, _23156_, _23155_);
  and (_27155_, _23157_, _25964_);
  and (_23158_, _17151_, _16390_);
  and (_23159_, _22659_, _17757_);
  and (_23160_, _23159_, _23158_);
  or (_23161_, _23160_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_23162_, ABINPUT[19]);
  nand (_23163_, _23160_, _23162_);
  and (_23164_, _23163_, _23161_);
  or (_23165_, _23164_, _23141_);
  not (_23166_, ABINPUT[11]);
  nand (_23167_, _23141_, _23166_);
  and (_23168_, _23167_, _25964_);
  and (_28332_, _23168_, _23165_);
  or (_23169_, _23144_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nand (_23170_, _23144_, _17475_);
  and (_23171_, _23170_, _23169_);
  or (_23172_, _23171_, _23141_);
  not (_23173_, ABINPUT[12]);
  nand (_23174_, _23141_, _23173_);
  and (_23175_, _23174_, _25964_);
  and (_28341_, _23175_, _23172_);
  or (_23176_, _23144_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nand (_23177_, _23144_, _17670_);
  and (_23178_, _23177_, _23176_);
  or (_23179_, _23178_, _23141_);
  not (_23180_, ABINPUT[13]);
  nand (_23181_, _23141_, _23180_);
  and (_23182_, _23181_, _25964_);
  and (_28349_, _23182_, _23179_);
  or (_23183_, _23160_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nand (_23184_, _23160_, _17845_);
  and (_23185_, _23184_, _23183_);
  or (_23186_, _23185_, _23141_);
  not (_23187_, ABINPUT[14]);
  nand (_23188_, _23141_, _23187_);
  and (_23189_, _23188_, _25964_);
  and (_28358_, _23189_, _23186_);
  or (_23190_, _23144_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand (_23191_, _23144_, _18019_);
  and (_23192_, _23191_, _23190_);
  or (_23193_, _23192_, _23141_);
  not (_23194_, ABINPUT[15]);
  nand (_23195_, _23141_, _23194_);
  and (_23196_, _23195_, _25964_);
  and (_28367_, _23196_, _23193_);
  or (_23197_, _23144_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nand (_23198_, _23144_, _18194_);
  and (_23199_, _23198_, _23197_);
  or (_23200_, _23199_, _23141_);
  not (_23201_, ABINPUT[16]);
  nand (_23202_, _23141_, _23201_);
  and (_23203_, _23202_, _25964_);
  and (_28376_, _23203_, _23200_);
  or (_23204_, _23160_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nand (_23205_, _23160_, _18368_);
  and (_23206_, _23205_, _23204_);
  or (_23207_, _23206_, _23141_);
  not (_23208_, ABINPUT[17]);
  nand (_23209_, _23141_, _23208_);
  and (_23210_, _23209_, _25964_);
  and (_28384_, _23210_, _23207_);
  and (_23211_, _23154_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nor (_23212_, _23154_, _23162_);
  or (_23213_, _23212_, _23211_);
  and (_28393_, _23213_, _25964_);
  and (_23214_, _23154_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nor (_23215_, _23154_, _17475_);
  or (_23216_, _23215_, _23214_);
  and (_28401_, _23216_, _25964_);
  and (_23217_, _23154_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nor (_23218_, _23154_, _17670_);
  or (_23219_, _23218_, _23217_);
  and (_28410_, _23219_, _25964_);
  and (_23220_, _23154_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nor (_23221_, _23154_, _17845_);
  or (_23222_, _23221_, _23220_);
  and (_28418_, _23222_, _25964_);
  and (_23223_, _23154_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nor (_23224_, _23154_, _18019_);
  or (_23225_, _23224_, _23223_);
  and (_28427_, _23225_, _25964_);
  and (_23226_, _23154_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nor (_23227_, _23154_, _18194_);
  or (_23228_, _23227_, _23226_);
  and (_28435_, _23228_, _25964_);
  and (_23229_, _23154_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nor (_23230_, _23154_, _18368_);
  or (_23231_, _23230_, _23229_);
  and (_28444_, _23231_, _25964_);
  nor (_23232_, _16205_, _16031_);
  and (_23233_, _16574_, _15889_);
  and (_23234_, _23233_, _23232_);
  and (_23235_, _23234_, _15585_);
  and (_23236_, _16988_, ABINPUT[0]);
  not (_23237_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_23238_, _16988_, _23237_);
  nor (_23239_, _23238_, _23236_);
  nand (_23240_, _23239_, _23235_);
  nor (_23241_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_23242_, _23241_, ABINPUT[0]);
  nand (_23243_, _23241_, _23237_);
  and (_23244_, _23243_, _23242_);
  or (_23245_, _23244_, _23235_);
  and (_23246_, _23245_, _23240_);
  and (_23247_, _17151_, _17107_);
  and (_23248_, _23247_, _23234_);
  not (_23249_, _23248_);
  and (_23250_, _23249_, _23246_);
  and (_23251_, _23248_, ABINPUT[10]);
  or (_23252_, _23251_, _23250_);
  and (_01600_, _23252_, _25964_);
  nand (_23253_, _23235_, _17388_);
  and (_23254_, _23253_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_23255_, _23235_, _17421_);
  or (_23256_, _23255_, _23248_);
  or (_23257_, _23256_, _23254_);
  not (_23258_, ABINPUT[4]);
  nand (_23259_, _23248_, _23258_);
  and (_23260_, _23259_, _23257_);
  and (_06381_, _23260_, _25964_);
  not (_23261_, _17583_);
  and (_23262_, _23261_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_23263_, _23262_, _17625_);
  nand (_23264_, _23263_, _23235_);
  and (_23265_, ABINPUT[2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_23266_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_23267_, _23266_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_23268_, _23267_, _23265_);
  or (_23269_, _23268_, _23235_);
  and (_23270_, _23269_, _23264_);
  and (_23271_, _23270_, _23249_);
  and (_23272_, _23248_, ABINPUT[5]);
  or (_23273_, _23272_, _23271_);
  and (_06392_, _23273_, _25964_);
  nand (_23274_, _23235_, _17757_);
  and (_23275_, _23274_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_23276_, _23235_, _17790_);
  or (_23277_, _23276_, _23275_);
  and (_23278_, _23277_, _23249_);
  and (_23279_, _23248_, ABINPUT[6]);
  or (_23280_, _23279_, _23278_);
  and (_06403_, _23280_, _25964_);
  nand (_23281_, _23235_, _17931_);
  and (_23282_, _23281_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_23283_, _23235_, _17964_);
  or (_23284_, _23283_, _23282_);
  and (_23285_, _23284_, _23249_);
  and (_23286_, _23248_, ABINPUT[7]);
  or (_23287_, _23286_, _23285_);
  and (_06414_, _23287_, _25964_);
  nand (_23288_, _23235_, _18106_);
  and (_23289_, _23288_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_23290_, _23235_, _18139_);
  or (_23291_, _23290_, _23248_);
  or (_23292_, _23291_, _23289_);
  not (_23293_, ABINPUT[8]);
  nand (_23294_, _23248_, _23293_);
  and (_23295_, _23294_, _23292_);
  and (_06425_, _23295_, _25964_);
  not (_23296_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_23297_, _18281_, _23296_);
  nor (_23298_, _23297_, _18313_);
  nand (_23299_, _23298_, _23235_);
  and (_23300_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_23301_, _23300_, ABINPUT[1]);
  nor (_23302_, _23300_, _23296_);
  or (_23303_, _23302_, _23301_);
  or (_23304_, _23303_, _23235_);
  and (_23305_, _23304_, _23299_);
  and (_23306_, _23305_, _23249_);
  and (_23307_, _23248_, ABINPUT[9]);
  or (_23308_, _23307_, _23306_);
  and (_06436_, _23308_, _25964_);
  not (_23309_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_23310_, _23140_, _23309_);
  and (_23311_, _23310_, ABINPUT[18]);
  nor (_23312_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_23313_, _23312_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_23314_, _17107_, _16390_);
  not (_23315_, _15889_);
  and (_23316_, _16564_, _23315_);
  and (_23317_, _23316_, _23232_);
  and (_23318_, _23317_, _23314_);
  and (_23319_, _23318_, _17151_);
  nor (_23320_, _23319_, _23313_);
  nor (_23321_, _23320_, _17086_);
  not (_23322_, _23320_);
  and (_23323_, _16564_, _16390_);
  and (_23324_, _23323_, _16042_);
  and (_23325_, _23324_, _16216_);
  and (_23326_, _23325_, _15585_);
  nand (_23327_, _23326_, _16988_);
  and (_23328_, _23327_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_23329_, _23326_, _23236_);
  nor (_23330_, _23329_, _23328_);
  nor (_23331_, _23330_, _23322_);
  nor (_23332_, _23331_, _23321_);
  nor (_23333_, _23332_, _23310_);
  nor (_23334_, _23333_, _23311_);
  nor (_07142_, _23334_, rst);
  not (_23335_, _23310_);
  and (_23336_, _23320_, _23335_);
  not (_23337_, _23336_);
  nand (_23338_, _23326_, _17107_);
  and (_23339_, _23338_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_23340_, _23326_, _17248_);
  nor (_23341_, _23340_, _23339_);
  nor (_23342_, _23341_, _23337_);
  not (_23343_, _23342_);
  and (_23344_, _23310_, ABINPUT[11]);
  or (_23345_, _23310_, _23162_);
  nor (_23346_, _23345_, _23320_);
  nor (_23347_, _23346_, _23344_);
  and (_23348_, _23347_, _23343_);
  nor (_08851_, _23348_, rst);
  and (_23349_, _23310_, ABINPUT[12]);
  nor (_23350_, _23320_, _17475_);
  or (_23351_, _23310_, _17388_);
  nand (_23352_, _23351_, _23326_);
  and (_23353_, _23352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_23354_, _23326_, _17421_);
  or (_23355_, _23354_, _23353_);
  and (_23356_, _23355_, _23320_);
  or (_23357_, _23356_, _23350_);
  and (_23358_, _23357_, _23335_);
  nor (_23359_, _23358_, _23349_);
  nor (_08862_, _23359_, rst);
  and (_23360_, _23310_, ABINPUT[13]);
  nand (_23361_, _23326_, _17583_);
  and (_23362_, _23361_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_23363_, _23326_, _17625_);
  nor (_23364_, _23363_, _23362_);
  nor (_23365_, _23364_, _23337_);
  nor (_23366_, _23320_, _17670_);
  or (_23367_, _23366_, _23365_);
  and (_23368_, _23367_, _23335_);
  nor (_23369_, _23368_, _23360_);
  nor (_08873_, _23369_, rst);
  and (_23370_, _23310_, ABINPUT[14]);
  nor (_23371_, _23320_, _17845_);
  nand (_23372_, _23326_, _17757_);
  and (_23373_, _23372_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_23374_, _23326_, _17790_);
  nor (_23375_, _23374_, _23373_);
  nor (_23376_, _23375_, _23322_);
  nor (_23377_, _23376_, _23371_);
  nor (_23378_, _23377_, _23310_);
  nor (_23379_, _23378_, _23370_);
  nor (_08884_, _23379_, rst);
  and (_23380_, _23310_, ABINPUT[15]);
  nand (_23381_, _23326_, _17931_);
  and (_23382_, _23381_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not (_23383_, _23382_);
  not (_23384_, _15585_);
  nor (_23385_, _23384_, _16205_);
  and (_23386_, _23385_, _16042_);
  and (_23387_, _23386_, _23323_);
  nand (_23388_, _23387_, _17964_);
  and (_23389_, _23388_, _23320_);
  and (_23390_, _23389_, _23383_);
  nor (_23391_, _23310_, _18019_);
  nor (_23392_, _23391_, _23336_);
  nor (_23393_, _23392_, _23390_);
  nor (_23394_, _23393_, _23380_);
  nor (_08895_, _23394_, rst);
  and (_23395_, _23310_, ABINPUT[16]);
  nor (_23396_, _23320_, _18194_);
  nand (_23397_, _23326_, _18106_);
  and (_23398_, _23397_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_23399_, _23326_, _18139_);
  nor (_23400_, _23399_, _23398_);
  nor (_23401_, _23400_, _23322_);
  nor (_23402_, _23401_, _23396_);
  nor (_23403_, _23402_, _23310_);
  nor (_23404_, _23403_, _23395_);
  nor (_08906_, _23404_, rst);
  nand (_23405_, _23326_, _18281_);
  and (_23406_, _23405_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_23407_, _23326_, _18313_);
  nor (_23408_, _23407_, _23406_);
  nor (_23409_, _23408_, _23337_);
  not (_23410_, _23409_);
  and (_23411_, _23310_, ABINPUT[17]);
  or (_23412_, _23310_, _18368_);
  nor (_23413_, _23412_, _23320_);
  nor (_23414_, _23413_, _23411_);
  and (_23415_, _23414_, _23410_);
  nor (_08917_, _23415_, rst);
  and (_23416_, _22670_, _16988_);
  or (_23417_, _23416_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nand (_23418_, _23416_, _17020_);
  and (_23419_, _23418_, _15585_);
  and (_23420_, _23419_, _23417_);
  not (_23421_, ABINPUT[10]);
  and (_23422_, _22659_, _23314_);
  nand (_23423_, _23422_, _23421_);
  or (_23424_, _23422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_23425_, _23424_, _17151_);
  and (_23426_, _23425_, _23423_);
  and (_23427_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_23428_, _23427_, rst);
  or (_23429_, _23428_, _23426_);
  or (_19486_, _23429_, _23420_);
  and (_23430_, _23233_, _22637_);
  and (_23431_, _23430_, _17107_);
  and (_23432_, _23431_, ABINPUT[10]);
  not (_23433_, _23431_);
  and (_23434_, _23433_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_23435_, _23434_, _23432_);
  and (_23436_, _23435_, _17151_);
  and (_23437_, _23430_, _16988_);
  nor (_23438_, _23437_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_23439_, _23437_, _17020_);
  or (_23440_, _23439_, _23384_);
  nor (_23441_, _23440_, _23438_);
  and (_23442_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_23443_, _23442_, rst);
  or (_23444_, _23443_, _23441_);
  or (_19509_, _23444_, _23436_);
  and (_23445_, _23316_, _22637_);
  and (_23446_, _23445_, _23314_);
  and (_23447_, _23446_, ABINPUT[10]);
  not (_23448_, _23446_);
  and (_23449_, _23448_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_23450_, _23449_, _23447_);
  and (_23451_, _23450_, _17151_);
  and (_23452_, _23445_, _16390_);
  not (_23453_, _16988_);
  and (_23454_, _23453_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_23455_, _23454_, _23236_);
  and (_23456_, _23455_, _23452_);
  not (_23457_, _23452_);
  and (_23458_, _23457_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_23459_, _23458_, _23456_);
  and (_23460_, _23459_, _15585_);
  and (_23461_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_23462_, _23461_, rst);
  or (_23463_, _23462_, _23460_);
  or (_19532_, _23463_, _23451_);
  nor (_23464_, _16564_, _15889_);
  and (_23465_, _22637_, _23464_);
  and (_23466_, _23465_, _23314_);
  and (_23467_, _23466_, ABINPUT[10]);
  not (_23468_, _23466_);
  and (_23469_, _23468_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_23470_, _23469_, _23467_);
  and (_23471_, _23470_, _17151_);
  and (_23472_, _23453_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_23473_, _23472_, _23236_);
  and (_23474_, _16031_, _23315_);
  and (_23475_, _23474_, _16585_);
  and (_23476_, _23475_, _23473_);
  not (_23477_, _23475_);
  and (_23478_, _23477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_23479_, _23478_, _23476_);
  and (_23480_, _23479_, _15585_);
  and (_23481_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_23482_, _23481_, rst);
  or (_23483_, _23482_, _23480_);
  or (_19555_, _23483_, _23471_);
  not (_23484_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_23485_, _23422_, _23484_);
  and (_23486_, _22670_, _17248_);
  or (_23487_, _23486_, _23485_);
  and (_23488_, _23487_, _15585_);
  and (_23489_, _23422_, ABINPUT[3]);
  or (_23490_, _23489_, _23485_);
  and (_23491_, _23490_, _17151_);
  nor (_23492_, _15574_, _23484_);
  or (_23493_, _23492_, rst);
  or (_23494_, _23493_, _23491_);
  or (_25391_, _23494_, _23488_);
  and (_23495_, _22681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_23496_, _22670_, _17421_);
  or (_23497_, _23496_, _23495_);
  and (_23498_, _23497_, _15585_);
  nand (_23499_, _23422_, _23258_);
  or (_23500_, _23422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_23501_, _23500_, _17151_);
  and (_23502_, _23501_, _23499_);
  and (_23503_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_23504_, _23503_, _23502_);
  or (_23505_, _23504_, _23498_);
  or (_25393_, _23505_, rst);
  not (_23506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_23507_, _23152_, _23506_);
  and (_23508_, _22670_, _17625_);
  or (_23509_, _23508_, _23507_);
  and (_23510_, _23509_, _15585_);
  or (_23511_, _23422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_23512_, _23511_, _17151_);
  not (_23513_, ABINPUT[5]);
  nand (_23514_, _23422_, _23513_);
  and (_23515_, _23514_, _23512_);
  nor (_23516_, _15574_, _23506_);
  or (_23517_, _23516_, rst);
  or (_23518_, _23517_, _23515_);
  or (_25395_, _23518_, _23510_);
  not (_23519_, ABINPUT[6]);
  nand (_23520_, _23422_, _23519_);
  or (_23521_, _23422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_23522_, _23521_, _17151_);
  and (_23523_, _23522_, _23520_);
  and (_23524_, _23143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_23525_, _22670_, _17790_);
  or (_23526_, _23525_, _23524_);
  and (_23527_, _23526_, _15585_);
  and (_23528_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_23529_, _23528_, rst);
  or (_23530_, _23529_, _23527_);
  or (_25397_, _23530_, _23523_);
  nand (_23531_, _22670_, _17931_);
  and (_23532_, _23531_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_23533_, _22670_, _17964_);
  or (_23534_, _23533_, _23532_);
  and (_23535_, _23534_, _15585_);
  not (_23536_, ABINPUT[7]);
  nand (_23537_, _23422_, _23536_);
  or (_23538_, _23422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_23539_, _23538_, _17151_);
  and (_23540_, _23539_, _23537_);
  and (_23541_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_23542_, _23541_, rst);
  or (_23543_, _23542_, _23540_);
  or (_25399_, _23543_, _23535_);
  nand (_23544_, _22670_, _18106_);
  and (_23545_, _23544_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_23546_, _22670_, _18139_);
  or (_23547_, _23546_, _23545_);
  and (_23548_, _23547_, _15585_);
  nand (_23549_, _23422_, _23293_);
  or (_23550_, _23422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_23551_, _23550_, _17151_);
  and (_23552_, _23551_, _23549_);
  and (_23553_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_23554_, _23553_, rst);
  or (_23555_, _23554_, _23552_);
  or (_25401_, _23555_, _23548_);
  nand (_23556_, _22670_, _18281_);
  and (_23557_, _23556_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_23558_, _22670_, _18313_);
  or (_23559_, _23558_, _23557_);
  and (_23560_, _23559_, _15585_);
  not (_23561_, ABINPUT[9]);
  nand (_23562_, _23422_, _23561_);
  or (_23563_, _23422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_23564_, _23563_, _17151_);
  and (_23565_, _23564_, _23562_);
  and (_23566_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_23567_, _23566_, rst);
  or (_23568_, _23567_, _23565_);
  or (_25403_, _23568_, _23560_);
  and (_23569_, _23433_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_23570_, _23431_, ABINPUT[3]);
  or (_23571_, _23570_, _23569_);
  and (_23572_, _23571_, _17151_);
  and (_23573_, _23430_, _17248_);
  or (_23574_, _23573_, _23569_);
  and (_23575_, _23574_, _15585_);
  and (_23576_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_23577_, _23576_, rst);
  or (_23578_, _23577_, _23575_);
  or (_25405_, _23578_, _23572_);
  and (_23579_, _23431_, ABINPUT[4]);
  and (_23580_, _23433_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_23581_, _23580_, _23579_);
  and (_23582_, _23581_, _17151_);
  nand (_23583_, _23430_, _17388_);
  and (_23584_, _23583_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_23585_, _23430_, _17421_);
  or (_23587_, _23585_, _23584_);
  and (_23588_, _23587_, _15585_);
  and (_23589_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_23590_, _23589_, rst);
  or (_23591_, _23590_, _23588_);
  or (_25407_, _23591_, _23582_);
  and (_23592_, _23431_, ABINPUT[5]);
  and (_23593_, _23433_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_23594_, _23593_, _23592_);
  and (_23595_, _23594_, _17151_);
  nand (_23597_, _23430_, _17583_);
  and (_23598_, _23597_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_23599_, _23430_, _17625_);
  or (_23600_, _23599_, _23598_);
  and (_23601_, _23600_, _15585_);
  and (_23602_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_23603_, _23602_, rst);
  or (_23604_, _23603_, _23601_);
  or (_25409_, _23604_, _23595_);
  and (_23605_, _23431_, ABINPUT[6]);
  and (_23607_, _23433_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_23608_, _23607_, _23605_);
  and (_23609_, _23608_, _17151_);
  and (_23610_, _23430_, _17757_);
  nor (_23611_, _23610_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_23612_, _23610_, _17020_);
  or (_23613_, _23612_, _23384_);
  nor (_23614_, _23613_, _23611_);
  and (_23615_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_23616_, _23615_, rst);
  or (_23618_, _23616_, _23614_);
  or (_25411_, _23618_, _23609_);
  and (_23619_, _23431_, ABINPUT[7]);
  and (_23620_, _23433_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_23621_, _23620_, _23619_);
  and (_23622_, _23621_, _17151_);
  nand (_23623_, _23430_, _17931_);
  and (_23624_, _23623_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_23625_, _23430_, _17964_);
  or (_23626_, _23625_, _23624_);
  and (_23628_, _23626_, _15585_);
  and (_23629_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_23630_, _23629_, rst);
  or (_23631_, _23630_, _23628_);
  or (_25413_, _23631_, _23622_);
  and (_23632_, _23431_, ABINPUT[8]);
  and (_23633_, _23433_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_23634_, _23633_, _23632_);
  and (_23635_, _23634_, _17151_);
  and (_23636_, _23430_, _18106_);
  nor (_23638_, _23636_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_23639_, _23636_, _17020_);
  or (_23640_, _23639_, _23384_);
  nor (_23641_, _23640_, _23638_);
  and (_23642_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_23643_, _23642_, rst);
  or (_23644_, _23643_, _23641_);
  or (_25415_, _23644_, _23635_);
  and (_23645_, _23431_, ABINPUT[9]);
  and (_23646_, _23433_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_23648_, _23646_, _23645_);
  and (_23649_, _23648_, _17151_);
  and (_23650_, _23430_, _18281_);
  nor (_23651_, _23650_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_23652_, _23650_, _17020_);
  or (_23653_, _23652_, _23384_);
  nor (_23654_, _23653_, _23651_);
  and (_23655_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_23656_, _23655_, rst);
  or (_23657_, _23656_, _23654_);
  or (_25417_, _23657_, _23649_);
  and (_23658_, _23446_, ABINPUT[3]);
  and (_23659_, _23448_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_23660_, _23659_, _23658_);
  and (_23661_, _23660_, _17151_);
  and (_23662_, _23457_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  not (_23663_, _17107_);
  and (_23664_, _23663_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_23665_, _23664_, _17248_);
  and (_23666_, _23665_, _23452_);
  or (_23667_, _23666_, _23662_);
  and (_23668_, _23667_, _15585_);
  and (_23669_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_23670_, _23669_, rst);
  or (_23671_, _23670_, _23668_);
  or (_25419_, _23671_, _23661_);
  and (_23672_, _23446_, ABINPUT[4]);
  and (_23673_, _23448_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_23674_, _23673_, _23672_);
  and (_23675_, _23674_, _17151_);
  not (_23676_, _17388_);
  and (_23677_, _23676_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_23678_, _23677_, _17421_);
  and (_23679_, _23678_, _23452_);
  and (_23680_, _23457_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_23681_, _23680_, _23679_);
  and (_23682_, _23681_, _15585_);
  and (_23683_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_23684_, _23683_, rst);
  or (_23685_, _23684_, _23682_);
  or (_25421_, _23685_, _23675_);
  and (_23686_, _23446_, ABINPUT[5]);
  and (_23687_, _23448_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_23688_, _23687_, _23686_);
  and (_23689_, _23688_, _17151_);
  and (_23690_, _23261_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_23691_, _23690_, _17625_);
  and (_23692_, _23691_, _23452_);
  and (_23693_, _23457_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_23694_, _23693_, _23692_);
  and (_23695_, _23694_, _15585_);
  and (_23696_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_23697_, _23696_, rst);
  or (_23698_, _23697_, _23695_);
  or (_25423_, _23698_, _23689_);
  and (_23699_, _23446_, ABINPUT[6]);
  and (_23700_, _23448_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_23701_, _23700_, _23699_);
  and (_23702_, _23701_, _17151_);
  not (_23703_, _17757_);
  and (_23704_, _23703_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_23705_, _23704_, _17790_);
  and (_23706_, _23705_, _23452_);
  and (_23707_, _23457_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_23708_, _23707_, _23706_);
  and (_23709_, _23708_, _15585_);
  and (_23710_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_23711_, _23710_, rst);
  or (_23712_, _23711_, _23709_);
  or (_25425_, _23712_, _23702_);
  and (_23713_, _23446_, ABINPUT[7]);
  and (_23714_, _23448_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_23715_, _23714_, _23713_);
  and (_23716_, _23715_, _17151_);
  not (_23717_, _17931_);
  and (_23718_, _23717_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_23719_, _23718_, _17964_);
  and (_23720_, _23719_, _23452_);
  and (_23721_, _23457_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_23722_, _23721_, _23720_);
  and (_23723_, _23722_, _15585_);
  and (_23724_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_23725_, _23724_, rst);
  or (_23726_, _23725_, _23723_);
  or (_25427_, _23726_, _23716_);
  and (_23727_, _23446_, ABINPUT[8]);
  and (_23728_, _23448_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_23729_, _23728_, _23727_);
  and (_23730_, _23729_, _17151_);
  not (_23731_, _18106_);
  and (_23732_, _23731_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_23733_, _23732_, _18139_);
  and (_23734_, _23733_, _23452_);
  and (_23735_, _23457_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_23736_, _23735_, _23734_);
  and (_23737_, _23736_, _15585_);
  and (_23738_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_23739_, _23738_, rst);
  or (_23740_, _23739_, _23737_);
  or (_25429_, _23740_, _23730_);
  and (_23741_, _23446_, ABINPUT[9]);
  and (_23742_, _23448_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_23743_, _23742_, _23741_);
  and (_23744_, _23743_, _17151_);
  not (_23745_, _18281_);
  and (_23746_, _23745_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_23747_, _23746_, _18313_);
  and (_23748_, _23747_, _23452_);
  and (_23749_, _23457_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_23750_, _23749_, _23748_);
  and (_23751_, _23750_, _15585_);
  and (_23752_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_23753_, _23752_, rst);
  or (_23754_, _23753_, _23751_);
  or (_25431_, _23754_, _23744_);
  and (_23755_, _23466_, ABINPUT[3]);
  and (_23756_, _23468_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_23757_, _23756_, _23755_);
  and (_23758_, _23757_, _17151_);
  and (_23759_, _23663_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_23760_, _23759_, _17248_);
  and (_23761_, _23760_, _23475_);
  and (_23762_, _23477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_23763_, _23762_, _23761_);
  and (_23764_, _23763_, _15585_);
  and (_23765_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_23766_, _23765_, rst);
  or (_23767_, _23766_, _23764_);
  or (_25433_, _23767_, _23758_);
  and (_23768_, _23466_, ABINPUT[4]);
  and (_23769_, _23468_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_23770_, _23769_, _23768_);
  and (_23771_, _23770_, _17151_);
  and (_23772_, _23676_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_23773_, _23772_, _17421_);
  and (_23774_, _23773_, _23475_);
  and (_23775_, _23477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_23776_, _23775_, _23774_);
  and (_23777_, _23776_, _15585_);
  and (_23778_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_23779_, _23778_, rst);
  or (_23780_, _23779_, _23777_);
  or (_25435_, _23780_, _23771_);
  and (_23781_, _23466_, ABINPUT[5]);
  and (_23782_, _23468_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_23783_, _23782_, _23781_);
  and (_23784_, _23783_, _17151_);
  and (_23785_, _23261_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_23786_, _23785_, _17625_);
  and (_23787_, _23786_, _23475_);
  and (_23788_, _23477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_23789_, _23788_, _23787_);
  and (_23790_, _23789_, _15585_);
  and (_23791_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_23792_, _23791_, rst);
  or (_23793_, _23792_, _23790_);
  or (_25437_, _23793_, _23784_);
  and (_23794_, _23466_, ABINPUT[6]);
  and (_23795_, _23468_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_23796_, _23795_, _23794_);
  and (_23797_, _23796_, _17151_);
  and (_23798_, _23703_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_23799_, _23798_, _17790_);
  and (_23800_, _23799_, _23475_);
  and (_23801_, _23477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_23802_, _23801_, _23800_);
  and (_23803_, _23802_, _15585_);
  and (_23804_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_23805_, _23804_, rst);
  or (_23806_, _23805_, _23803_);
  or (_25439_, _23806_, _23797_);
  and (_23807_, _23466_, ABINPUT[7]);
  and (_23808_, _23468_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_23809_, _23808_, _23807_);
  and (_23810_, _23809_, _17151_);
  and (_23811_, _23717_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_23812_, _23811_, _17964_);
  and (_23813_, _23812_, _23475_);
  and (_23814_, _23477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_23815_, _23814_, _23813_);
  and (_23816_, _23815_, _15585_);
  and (_23817_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_23818_, _23817_, rst);
  or (_23819_, _23818_, _23816_);
  or (_25441_, _23819_, _23810_);
  and (_23820_, _23466_, ABINPUT[8]);
  and (_23821_, _23468_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_23822_, _23821_, _23820_);
  and (_23823_, _23822_, _17151_);
  and (_23824_, _23731_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_23825_, _23824_, _18139_);
  and (_23826_, _23825_, _23475_);
  and (_23827_, _23477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_23828_, _23827_, _23826_);
  and (_23829_, _23828_, _15585_);
  and (_23830_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_23831_, _23830_, rst);
  or (_23832_, _23831_, _23829_);
  or (_25443_, _23832_, _23823_);
  and (_23833_, _23466_, ABINPUT[9]);
  and (_23834_, _23468_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_23835_, _23834_, _23833_);
  and (_23836_, _23835_, _17151_);
  and (_23837_, _23745_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_23838_, _23837_, _18313_);
  and (_23839_, _23838_, _23475_);
  and (_23840_, _23477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_23841_, _23840_, _23839_);
  and (_23842_, _23841_, _15585_);
  and (_23843_, _17064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_23844_, _23843_, rst);
  or (_23845_, _23844_, _23842_);
  or (_25445_, _23845_, _23836_);
  and (_23846_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_23847_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _25964_);
  and (_25967_, _23847_, _23846_);
  and (_23848_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_23849_, _23848_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_23850_, _23849_);
  and (_23851_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_23852_, _23851_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_23853_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_23854_, _23853_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor (_23855_, _23854_, _23852_);
  and (_23856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_23857_, _23856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  not (_23858_, _23857_);
  and (_23859_, _23858_, _23855_);
  and (_23860_, _23859_, _23850_);
  not (_23861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_23862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_23863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_23864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_23865_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _23864_);
  or (_23866_, _23865_, _23863_);
  nor (_23867_, _23866_, _23862_);
  nor (_23868_, _23867_, _23861_);
  nor (_23869_, _23868_, _23860_);
  and (_23870_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _23861_);
  not (_23871_, _23870_);
  not (_23872_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_23873_, _23851_, _23872_);
  not (_23874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_23875_, _23853_, _23874_);
  nor (_23876_, _23875_, _23873_);
  not (_23877_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_23878_, _23848_, _23877_);
  not (_23879_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_23880_, _23856_, _23879_);
  nor (_23881_, _23880_, _23878_);
  and (_23882_, _23881_, _23876_);
  nor (_23883_, _23882_, _23871_);
  nor (_23884_, _23883_, _23869_);
  and (_23885_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  not (_23886_, _23869_);
  nor (_23887_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _23864_);
  and (_23888_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _23864_);
  nor (_23889_, _23888_, _23887_);
  nor (_23890_, _23889_, _23886_);
  or (_23891_, _23890_, _23885_);
  or (_23892_, _23891_, _23846_);
  not (_23893_, _23846_);
  or (_23894_, _23889_, _23893_);
  and (_23895_, _23894_, _25964_);
  and (_25969_, _23895_, _23892_);
  nand (_23896_, _23860_, _23861_);
  or (_23897_, _23896_, _23883_);
  nand (_23898_, _23887_, _23846_);
  and (_23899_, _23898_, _25964_);
  and (_25972_, _23899_, _23897_);
  and (_23900_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_23901_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_23902_, _23901_, _23859_);
  and (_23903_, _23849_, _23864_);
  not (_23904_, _23855_);
  or (_23905_, _23904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_23906_, _23905_, _23903_);
  and (_23907_, _23906_, _23902_);
  and (_23908_, _23907_, _23869_);
  or (_23909_, _23908_, _23900_);
  and (_23910_, _23883_, _23886_);
  and (_23911_, _23878_, _23864_);
  or (_23912_, _23911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  not (_23913_, _23876_);
  and (_23914_, _23880_, _23864_);
  nor (_23915_, _23914_, _23913_);
  and (_23916_, _23915_, _23912_);
  and (_23917_, _23901_, _23913_);
  or (_23918_, _23917_, _23916_);
  and (_23919_, _23918_, _23910_);
  or (_23920_, _23919_, _23846_);
  or (_23921_, _23920_, _23909_);
  or (_23922_, _23893_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_23923_, _23922_, _25964_);
  and (_25975_, _23923_, _23921_);
  and (_23924_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_23925_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _23864_);
  or (_23926_, _23925_, _23859_);
  and (_23927_, _23849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_23928_, _23904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_23929_, _23928_, _23927_);
  and (_23930_, _23929_, _23926_);
  and (_23931_, _23930_, _23869_);
  or (_23932_, _23931_, _23924_);
  and (_23933_, _23878_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_23934_, _23933_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_23935_, _23880_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_23936_, _23935_, _23913_);
  and (_23937_, _23936_, _23934_);
  and (_23938_, _23925_, _23913_);
  or (_23939_, _23938_, _23937_);
  and (_23940_, _23939_, _23910_);
  or (_23941_, _23940_, _23846_);
  or (_23942_, _23941_, _23932_);
  or (_23943_, _23893_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_23944_, _23943_, _25964_);
  and (_25978_, _23944_, _23942_);
  nor (_23945_, _23846_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_23946_, _23945_, _23869_);
  nand (_23947_, _23945_, _23883_);
  and (_23948_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _25964_);
  nand (_23949_, _23948_, _23947_);
  nor (_25979_, _23949_, _23946_);
  nor (_23950_, _23846_, _23864_);
  and (_23951_, _23950_, _23869_);
  nand (_23952_, _23950_, _23883_);
  and (_23953_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _25964_);
  nand (_23954_, _23953_, _23952_);
  nor (_25981_, _23954_, _23951_);
  nor (_23955_, _23384_, _16390_);
  and (_23956_, _23955_, _22659_);
  and (_23957_, _23956_, _17757_);
  nand (_23958_, _23957_, _17020_);
  and (_23959_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_23960_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _23864_);
  and (_23961_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_23962_, _23961_, _23960_);
  nor (_23963_, _23962_, _23861_);
  nand (_23964_, _23963_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and (_23965_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _23864_);
  and (_23966_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_23967_, _23966_, _23965_);
  nor (_23968_, _23967_, _23861_);
  nor (_23969_, _23925_, _23901_);
  nand (_23970_, _23969_, _23968_);
  or (_23971_, _23970_, _23964_);
  and (_23972_, _23971_, _23959_);
  or (_23973_, _23972_, _23957_);
  and (_23974_, _23973_, _23958_);
  and (_23975_, _23247_, _16400_);
  and (_23976_, _23975_, _22659_);
  or (_23977_, _23976_, _23974_);
  nand (_23978_, _23976_, _23519_);
  and (_23979_, _23978_, _25964_);
  and (_26016_, _23979_, _23977_);
  not (_23980_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_23981_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _23980_);
  nor (_23982_, _23969_, _23861_);
  or (_23983_, _23982_, _23968_);
  or (_23984_, _23983_, _23964_);
  and (_23985_, _23984_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_23986_, _23985_, _23981_);
  nand (_23987_, _23956_, _17388_);
  and (_23988_, _23987_, _23986_);
  nor (_23989_, _23987_, _17020_);
  or (_23990_, _23989_, _23976_);
  or (_23991_, _23990_, _23988_);
  nand (_23992_, _23976_, _23258_);
  and (_23993_, _23992_, _25964_);
  and (_26018_, _23993_, _23991_);
  not (_23994_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_23995_, _23963_, _23994_);
  or (_23996_, _23995_, _23970_);
  nand (_23997_, _23996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_23998_, _23956_, _18106_);
  nor (_23999_, _23998_, _23997_);
  and (_24000_, _23998_, ABINPUT[0]);
  or (_24001_, _24000_, _23976_);
  or (_24002_, _24001_, _23999_);
  nand (_24003_, _23976_, _23293_);
  and (_24004_, _24003_, _25964_);
  and (_26020_, _24004_, _24002_);
  nand (_24005_, _23982_, _23967_);
  or (_24006_, _24005_, _23995_);
  nand (_24007_, _24006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_24008_, _23956_, _16988_);
  nor (_24009_, _24008_, _24007_);
  and (_24010_, _24008_, ABINPUT[0]);
  or (_24011_, _24010_, _23976_);
  or (_24012_, _24011_, _24009_);
  nand (_24013_, _23976_, _23421_);
  and (_24014_, _24013_, _25964_);
  and (_26022_, _24014_, _24012_);
  nand (_24015_, _23956_, _18281_);
  and (_24016_, _24015_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_24017_, _23956_, _18313_);
  or (_24018_, _24017_, _23976_);
  or (_24019_, _24018_, _24016_);
  nand (_24020_, _23976_, _23561_);
  and (_24021_, _24020_, _25964_);
  and (_26024_, _24021_, _24019_);
  and (_24022_, _23975_, _23445_);
  and (_24023_, _23955_, _23445_);
  and (_24024_, _24023_, _16988_);
  nand (_24025_, _24024_, _17020_);
  or (_24026_, _24024_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_24027_, _24026_, _24025_);
  or (_24028_, _24027_, _24022_);
  nand (_24029_, _24022_, _23421_);
  and (_24030_, _24029_, _25964_);
  and (_26027_, _24030_, _24028_);
  and (_24031_, _23975_, _23465_);
  not (_24032_, _16564_);
  and (_24033_, _23955_, _24032_);
  and (_24034_, _24033_, _16216_);
  and (_24035_, _24034_, _23474_);
  and (_24036_, _24035_, _16988_);
  nand (_24037_, _24036_, _17020_);
  or (_24038_, _24036_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_24039_, _24038_, _24037_);
  or (_24040_, _24039_, _24031_);
  nand (_24041_, _24031_, _23421_);
  and (_24042_, _24041_, _25964_);
  and (_26028_, _24042_, _24040_);
  nor (_24043_, _23884_, _23846_);
  and (_24044_, _23846_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_24045_, _24044_, _24043_);
  and (_26952_, _24045_, _25964_);
  and (_24046_, _23846_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_24047_, _24046_, _24043_);
  and (_26954_, _24047_, _25964_);
  and (_24048_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _25964_);
  and (_26956_, _24048_, _23846_);
  not (_24049_, _23875_);
  nor (_24050_, _23878_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_24051_, _24050_, _23880_);
  or (_24052_, _24051_, _23873_);
  and (_24053_, _24052_, _24049_);
  and (_24054_, _24053_, _23910_);
  not (_24055_, _23854_);
  or (_24056_, _23849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_24057_, _24056_, _23858_);
  or (_24058_, _24057_, _23852_);
  and (_24059_, _24058_, _24055_);
  and (_24060_, _24059_, _23869_);
  or (_24061_, _24060_, _23846_);
  or (_24062_, _24061_, _24054_);
  or (_24063_, _23893_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_24064_, _24063_, _25964_);
  and (_26958_, _24064_, _24062_);
  nand (_24065_, _23876_, _23870_);
  nor (_24066_, _24065_, _23881_);
  or (_24067_, _24066_, _23869_);
  nand (_24068_, _23869_, _23904_);
  and (_24069_, _24068_, _24067_);
  or (_24070_, _24069_, _23846_);
  or (_24071_, _23893_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_24072_, _24071_, _25964_);
  and (_26960_, _24072_, _24070_);
  and (_24073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _25964_);
  and (_26962_, _24073_, _23846_);
  and (_24074_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _25964_);
  and (_26964_, _24074_, _23846_);
  nand (_24075_, _23945_, _23884_);
  nor (_24076_, _23869_, _23846_);
  or (_24077_, _24076_, _23864_);
  and (_24078_, _24077_, _25964_);
  and (_26966_, _24078_, _24075_);
  not (_24079_, _24043_);
  and (_24080_, _24079_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_24081_, _23903_);
  and (_24082_, _24081_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_24083_, _23857_, _23864_);
  or (_24084_, _24083_, _23852_);
  or (_24085_, _24084_, _24082_);
  not (_24086_, _23852_);
  or (_24087_, _23961_, _24086_);
  and (_24088_, _24087_, _24085_);
  or (_24089_, _24088_, _23854_);
  or (_24090_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _23864_);
  or (_24091_, _24090_, _24055_);
  and (_24092_, _24091_, _23869_);
  and (_24093_, _24092_, _24089_);
  not (_24094_, _23911_);
  and (_24095_, _24094_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_24096_, _23914_, _23873_);
  or (_24097_, _24096_, _24095_);
  not (_24098_, _23873_);
  or (_24099_, _23961_, _24098_);
  and (_24100_, _24099_, _24049_);
  and (_24101_, _24100_, _24097_);
  and (_24102_, _24090_, _23875_);
  or (_24103_, _24102_, _24101_);
  and (_24104_, _24103_, _23910_);
  or (_24105_, _24104_, _24093_);
  and (_24106_, _24105_, _23893_);
  or (_24107_, _24106_, _24080_);
  and (_26968_, _24107_, _25964_);
  and (_24108_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_24109_, _24108_, _23846_);
  and (_24110_, _24081_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_24111_, _24110_, _24084_);
  or (_24112_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _23864_);
  or (_24113_, _24112_, _24086_);
  and (_24114_, _24113_, _24111_);
  or (_24115_, _24114_, _23854_);
  or (_24116_, _23966_, _24055_);
  and (_24118_, _24116_, _23869_);
  and (_24119_, _24118_, _24115_);
  and (_24120_, _24094_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_24121_, _24120_, _24096_);
  or (_24122_, _24112_, _24098_);
  and (_24123_, _24122_, _24049_);
  and (_24124_, _24123_, _24121_);
  and (_24125_, _23966_, _23875_);
  or (_24126_, _24125_, _24124_);
  and (_24127_, _24126_, _23910_);
  or (_24128_, _24127_, _24119_);
  or (_24129_, _24128_, _24109_);
  or (_24130_, _23893_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_24131_, _24130_, _25964_);
  and (_26970_, _24131_, _24129_);
  and (_24132_, _24079_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not (_24133_, _23927_);
  and (_24134_, _24133_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_24135_, _23857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_24136_, _24135_, _23852_);
  or (_24138_, _24136_, _24134_);
  or (_24139_, _23960_, _24086_);
  and (_24140_, _24139_, _24138_);
  or (_24141_, _24140_, _23854_);
  or (_24142_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_24143_, _24142_, _24055_);
  and (_24144_, _24143_, _23869_);
  and (_24145_, _24144_, _24141_);
  not (_24146_, _23933_);
  and (_24147_, _24146_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_24148_, _23935_, _23873_);
  or (_24149_, _24148_, _24147_);
  or (_24150_, _23960_, _24098_);
  and (_24151_, _24150_, _24049_);
  and (_24152_, _24151_, _24149_);
  and (_24153_, _24142_, _23875_);
  or (_24154_, _24153_, _24152_);
  and (_24155_, _24154_, _23910_);
  or (_24156_, _24155_, _24145_);
  and (_24157_, _24156_, _23893_);
  or (_24158_, _24157_, _24132_);
  and (_26972_, _24158_, _25964_);
  and (_24159_, _23884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_24160_, _24159_, _23846_);
  and (_24161_, _24133_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_24162_, _24161_, _24136_);
  or (_24163_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_24164_, _24163_, _24086_);
  and (_24165_, _24164_, _24162_);
  or (_24166_, _24165_, _23854_);
  or (_24167_, _23965_, _24055_);
  and (_24168_, _24167_, _23869_);
  and (_24169_, _24168_, _24166_);
  and (_24170_, _24146_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_24171_, _24170_, _24148_);
  or (_24172_, _24163_, _24098_);
  and (_24173_, _24172_, _24049_);
  and (_24174_, _24173_, _24171_);
  and (_24175_, _23965_, _23875_);
  or (_24176_, _24175_, _24174_);
  and (_24177_, _24176_, _23910_);
  or (_24178_, _24177_, _24169_);
  or (_24179_, _24178_, _24160_);
  or (_24180_, _23893_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_24181_, _24180_, _25964_);
  and (_26974_, _24181_, _24179_);
  and (_24182_, _23947_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_24183_, _24182_, _23946_);
  and (_26976_, _24183_, _25964_);
  and (_24184_, _23952_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_24185_, _24184_, _23951_);
  and (_26978_, _24185_, _25964_);
  and (_24186_, _23956_, _17107_);
  nand (_24187_, _24186_, _17020_);
  or (_24188_, _24186_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_24189_, _24188_, _24187_);
  or (_24190_, _24189_, _23976_);
  not (_24191_, ABINPUT[3]);
  nand (_24192_, _23976_, _24191_);
  and (_24193_, _24192_, _25964_);
  and (_26980_, _24193_, _24190_);
  nand (_24194_, _23956_, _17583_);
  and (_24195_, _24194_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_24196_, _23956_, _17625_);
  or (_24197_, _24196_, _23976_);
  or (_24198_, _24197_, _24195_);
  nand (_24199_, _23976_, _23513_);
  and (_24200_, _24199_, _25964_);
  and (_26982_, _24200_, _24198_);
  nand (_24201_, _23956_, _17931_);
  and (_24202_, _24201_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_24203_, _23956_, _17964_);
  or (_24204_, _24203_, _23976_);
  or (_24205_, _24204_, _24202_);
  nand (_24206_, _23976_, _23536_);
  and (_24207_, _24206_, _25964_);
  and (_26984_, _24207_, _24205_);
  nand (_24208_, _24023_, _17107_);
  and (_24209_, _24208_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_24210_, _24023_, _17248_);
  or (_24211_, _24210_, _24022_);
  or (_24212_, _24211_, _24209_);
  nand (_24213_, _24022_, _24191_);
  and (_24214_, _24213_, _25964_);
  and (_26986_, _24214_, _24212_);
  nand (_24215_, _24023_, _17388_);
  and (_24216_, _24215_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_24217_, _24023_, _17421_);
  or (_24218_, _24217_, _24022_);
  or (_24219_, _24218_, _24216_);
  nand (_24220_, _24022_, _23258_);
  and (_24221_, _24220_, _25964_);
  and (_26988_, _24221_, _24219_);
  and (_24222_, _24023_, _17583_);
  or (_24223_, _24222_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nand (_24224_, _24222_, _17020_);
  and (_24225_, _24224_, _24223_);
  or (_24226_, _24225_, _24022_);
  nand (_24227_, _24022_, _23513_);
  and (_24228_, _24227_, _25964_);
  and (_26990_, _24228_, _24226_);
  nand (_24229_, _24023_, _17757_);
  and (_24230_, _24229_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_24231_, _24023_, _17790_);
  or (_24232_, _24231_, _24022_);
  or (_24233_, _24232_, _24230_);
  nand (_24234_, _24022_, _23519_);
  and (_24235_, _24234_, _25964_);
  and (_26991_, _24235_, _24233_);
  nand (_24236_, _24023_, _17931_);
  and (_24237_, _24236_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_24238_, _24023_, _17964_);
  or (_24239_, _24238_, _24022_);
  or (_24240_, _24239_, _24237_);
  nand (_24241_, _24022_, _23536_);
  and (_24242_, _24241_, _25964_);
  and (_26993_, _24242_, _24240_);
  nand (_24243_, _24023_, _18106_);
  and (_24244_, _24243_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_24245_, _24023_, _18139_);
  or (_24246_, _24245_, _24022_);
  or (_24247_, _24246_, _24244_);
  nand (_24248_, _24022_, _23293_);
  and (_24249_, _24248_, _25964_);
  and (_26995_, _24249_, _24247_);
  nand (_24250_, _24023_, _18281_);
  and (_24251_, _24250_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_24252_, _24023_, _18313_);
  or (_24253_, _24252_, _24022_);
  or (_24254_, _24253_, _24251_);
  nand (_24255_, _24022_, _23561_);
  and (_24256_, _24255_, _25964_);
  and (_26997_, _24256_, _24254_);
  and (_24257_, _24035_, _17107_);
  nand (_24258_, _24257_, _17020_);
  or (_24259_, _24257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_24260_, _24259_, _24258_);
  or (_24261_, _24260_, _24031_);
  nand (_24262_, _24031_, _24191_);
  and (_24263_, _24262_, _25964_);
  and (_26999_, _24263_, _24261_);
  nand (_24264_, _24035_, _17388_);
  and (_24265_, _24264_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_24266_, _24035_, _17421_);
  or (_24267_, _24266_, _24031_);
  or (_24268_, _24267_, _24265_);
  nand (_24269_, _24031_, _23258_);
  and (_24270_, _24269_, _25964_);
  and (_27001_, _24270_, _24268_);
  and (_24271_, _24035_, _17583_);
  or (_24272_, _24271_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nand (_24273_, _24271_, _17020_);
  and (_24274_, _24273_, _24272_);
  or (_24275_, _24274_, _24031_);
  nand (_24276_, _24031_, _23513_);
  and (_24277_, _24276_, _25964_);
  and (_27003_, _24277_, _24275_);
  nand (_24278_, _24035_, _17757_);
  and (_24279_, _24278_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_24280_, _24035_, _17790_);
  or (_24281_, _24280_, _24031_);
  or (_24282_, _24281_, _24279_);
  nand (_24283_, _24031_, _23519_);
  and (_24284_, _24283_, _25964_);
  and (_27005_, _24284_, _24282_);
  nand (_24285_, _24035_, _17931_);
  and (_24296_, _24285_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_24298_, _24035_, _17964_);
  or (_24299_, _24298_, _24031_);
  or (_24300_, _24299_, _24296_);
  nand (_24301_, _24031_, _23536_);
  and (_24302_, _24301_, _25964_);
  and (_27007_, _24302_, _24300_);
  nand (_24303_, _24035_, _18106_);
  and (_24304_, _24303_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_24305_, _24035_, _18139_);
  or (_24306_, _24305_, _24031_);
  or (_24307_, _24306_, _24304_);
  nand (_24308_, _24031_, _23293_);
  and (_24309_, _24308_, _25964_);
  and (_27009_, _24309_, _24307_);
  nand (_24310_, _24035_, _18281_);
  and (_24311_, _24310_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_24312_, _24035_, _18313_);
  or (_24313_, _24312_, _24031_);
  or (_24314_, _24313_, _24311_);
  nand (_24315_, _24031_, _23561_);
  and (_24316_, _24315_, _25964_);
  and (_27011_, _24316_, _24314_);
  not (_24317_, _22572_);
  nor (_24318_, _24317_, _22188_);
  not (_24319_, _18521_);
  and (_24320_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_24321_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_24322_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_24323_, _24322_, _24321_);
  and (_24324_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_24325_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_24326_, _24325_, _24324_);
  and (_24327_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_24328_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_24329_, _24328_, _24327_);
  and (_24330_, _24329_, _24326_);
  and (_24331_, _24330_, _24323_);
  nor (_24332_, _18850_, _24319_);
  not (_24333_, _24332_);
  nor (_24334_, _24333_, _24331_);
  nor (_24335_, _24334_, _24320_);
  not (_24336_, _24335_);
  and (_24337_, _24336_, _24318_);
  not (_24338_, _24337_);
  and (_24339_, _24317_, _22188_);
  and (_24340_, _24339_, _21114_);
  and (_24341_, _15552_, _16183_);
  nor (_24342_, _16727_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_24343_, _24342_, _16966_);
  and (_24344_, _24343_, _24341_);
  and (_24345_, _19984_, _16846_);
  nor (_24346_, _19984_, _16846_);
  nor (_24347_, _24346_, _24345_);
  and (_24348_, _24347_, _24344_);
  and (_24349_, _23249_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_24350_, _24349_, _23279_);
  and (_24351_, _24350_, _16400_);
  nor (_24352_, _24350_, _16400_);
  nor (_24353_, _24352_, _24351_);
  and (_24354_, _24353_, _24348_);
  nor (_24355_, _24350_, _19984_);
  and (_24356_, _24355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_24357_, _24350_, _19984_);
  and (_24358_, _24357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_24359_, _24358_, _24356_);
  nor (_24360_, _24350_, _21136_);
  and (_24361_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_24362_, _24350_, _21136_);
  and (_24363_, _24362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_24364_, _24363_, _24361_);
  and (_24365_, _24364_, _24359_);
  nor (_24366_, _24365_, _24354_);
  and (_24367_, _24354_, ABINPUT[10]);
  nor (_24368_, _24367_, _24366_);
  not (_24369_, _24368_);
  and (_24370_, _24369_, _24340_);
  not (_24371_, _24370_);
  not (_24372_, _21114_);
  not (_24373_, _22583_);
  nor (_24374_, _23072_, _24373_);
  nor (_24375_, _24374_, _24372_);
  and (_24376_, _24375_, _24371_);
  and (_24377_, _24376_, _24338_);
  not (_24378_, _18477_);
  or (_24379_, _21870_, _21827_);
  or (_24380_, _21794_, _21158_);
  or (_24381_, _24380_, _24379_);
  not (_24382_, _21925_);
  nor (_24383_, _24382_, _21223_);
  nand (_24384_, _24383_, _21487_);
  or (_24385_, _24384_, _24381_);
  and (_24386_, _24385_, _24378_);
  and (_24387_, _21421_, _20949_);
  nor (_24388_, _22090_, _24387_);
  not (_24389_, _20916_);
  nor (_24390_, _24389_, _24388_);
  nor (_24391_, _24390_, _24386_);
  not (_24392_, _24391_);
  and (_24393_, _24392_, _24377_);
  and (_24394_, _24357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_24395_, _24355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_24396_, _24395_, _24394_);
  and (_24397_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_24398_, _24362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_24399_, _24398_, _24397_);
  and (_24400_, _24399_, _24396_);
  nor (_24401_, _24400_, _24354_);
  and (_24402_, _24354_, ABINPUT[8]);
  nor (_24403_, _24402_, _24401_);
  not (_24404_, _24403_);
  and (_24405_, _24404_, _24340_);
  and (_24406_, _24318_, _21114_);
  and (_24407_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_24408_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_24409_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_24410_, _24409_, _24408_);
  and (_24411_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_24412_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_24413_, _24412_, _24411_);
  and (_24414_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_24415_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_24416_, _24415_, _24414_);
  and (_24417_, _24416_, _24413_);
  and (_24418_, _24417_, _24410_);
  nor (_24419_, _24418_, _24333_);
  nor (_24420_, _24419_, _24407_);
  not (_24421_, _24420_);
  and (_24422_, _24421_, _24406_);
  nor (_24423_, _24422_, _24405_);
  and (_24424_, _22572_, _22188_);
  and (_24425_, _24424_, _24372_);
  and (_24426_, _23133_, _21114_);
  nor (_24427_, _24426_, _24373_);
  or (_24428_, _24427_, _24425_);
  not (_24429_, _24428_);
  and (_24430_, _24429_, _24423_);
  not (_24431_, _24430_);
  and (_24432_, _24431_, _24393_);
  and (_24433_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_24434_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_24435_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_24436_, _24435_, _24434_);
  and (_24437_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_24438_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_24439_, _24438_, _24437_);
  and (_24440_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_24441_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_24442_, _24441_, _24440_);
  and (_24443_, _24442_, _24439_);
  and (_24444_, _24443_, _24436_);
  nor (_24445_, _24444_, _24333_);
  nor (_24446_, _24445_, _24433_);
  not (_24447_, _24446_);
  and (_24448_, _24447_, _24406_);
  and (_24449_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_24450_, _24357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_24451_, _24450_, _24449_);
  and (_24452_, _24362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_24453_, _24355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_24454_, _24453_, _24452_);
  and (_24455_, _24454_, _24451_);
  nor (_24456_, _24455_, _24354_);
  and (_24457_, _24354_, ABINPUT[5]);
  nor (_24458_, _24457_, _24456_);
  not (_24459_, _24458_);
  and (_24460_, _24459_, _24340_);
  nor (_24461_, _24460_, _24448_);
  not (_24462_, _23115_);
  and (_24463_, _24462_, _22594_);
  and (_24464_, _24424_, _21114_);
  and (_24465_, _24464_, _20467_);
  nor (_24466_, _24465_, _24463_);
  and (_24467_, _24466_, _24461_);
  nor (_24468_, _24467_, _24392_);
  nor (_24469_, _24468_, _24432_);
  and (_24470_, _16205_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_24471_, _24470_, _23315_);
  nor (_24472_, _16716_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_24473_, _24472_, _24471_);
  not (_24474_, _24473_);
  and (_24475_, _24474_, _24469_);
  not (_24476_, _24350_);
  and (_24477_, _24464_, _24476_);
  and (_24478_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_24479_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_24480_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_24481_, _24480_, _24479_);
  and (_24482_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_24483_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_24484_, _24483_, _24482_);
  and (_24485_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_24486_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_24487_, _24486_, _24485_);
  and (_24488_, _24487_, _24484_);
  and (_24489_, _24488_, _24481_);
  nor (_24490_, _24489_, _24333_);
  nor (_24491_, _24490_, _24478_);
  not (_24492_, _24491_);
  and (_24493_, _24492_, _24406_);
  nor (_24494_, _24493_, _24477_);
  not (_24495_, _23121_);
  and (_24496_, _24495_, _22594_);
  and (_24497_, _24357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_24498_, _24355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_24499_, _24498_, _24497_);
  and (_24500_, _24362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  not (_24501_, _24500_);
  and (_24502_, _24501_, _24499_);
  and (_24503_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_24504_, _24503_, _24354_);
  and (_24505_, _24504_, _24502_);
  and (_24506_, _24354_, _23519_);
  or (_24507_, _24506_, _24505_);
  not (_24508_, _24507_);
  and (_24509_, _24508_, _24340_);
  nor (_24510_, _24509_, _24496_);
  and (_24511_, _24510_, _24494_);
  not (_24512_, _24511_);
  and (_24513_, _24512_, _24393_);
  and (_24514_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_24515_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_24516_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_24517_, _24516_, _24515_);
  and (_24518_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_24519_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_24520_, _24519_, _24518_);
  and (_24521_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_24522_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_24523_, _24522_, _24521_);
  and (_24524_, _24523_, _24520_);
  and (_24525_, _24524_, _24517_);
  nor (_24526_, _24525_, _24333_);
  nor (_24527_, _24526_, _24514_);
  not (_24528_, _24527_);
  and (_24529_, _24528_, _24406_);
  and (_24530_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_24531_, _24357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_24532_, _24531_, _24530_);
  and (_24533_, _24362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_24534_, _24355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_24535_, _24534_, _24533_);
  and (_24536_, _24535_, _24532_);
  nor (_24537_, _24536_, _24354_);
  and (_24538_, _24354_, ABINPUT[3]);
  nor (_24539_, _24538_, _24537_);
  not (_24540_, _24539_);
  and (_24541_, _24540_, _24340_);
  nor (_24542_, _24541_, _24529_);
  not (_24543_, _23103_);
  and (_24544_, _24543_, _22594_);
  and (_24545_, _24464_, _19984_);
  nor (_24546_, _24545_, _24544_);
  and (_24547_, _24546_, _24542_);
  nor (_24548_, _24547_, _24392_);
  nor (_24549_, _24548_, _24513_);
  and (_24550_, _24470_, _16400_);
  nor (_24551_, _16846_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_24552_, _24551_, _24550_);
  not (_24553_, _24552_);
  nor (_24554_, _24553_, _24549_);
  nor (_24555_, _24554_, _24475_);
  nor (_24556_, _24474_, _24469_);
  not (_24557_, _24556_);
  and (_24558_, _24357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_24559_, _24355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_24560_, _24559_, _24558_);
  and (_24561_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_24562_, _24362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_24563_, _24562_, _24561_);
  and (_24564_, _24563_, _24560_);
  nor (_24565_, _24564_, _24354_);
  and (_24566_, _24354_, ABINPUT[9]);
  nor (_24567_, _24566_, _24565_);
  not (_24568_, _24567_);
  and (_24569_, _24568_, _24340_);
  not (_24570_, _23139_);
  and (_24571_, _24570_, _22594_);
  nor (_24572_, _24571_, _24569_);
  and (_24573_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_24574_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_24575_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_24576_, _24575_, _24574_);
  and (_24577_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_24578_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_24579_, _24578_, _24577_);
  and (_24580_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_24581_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_24582_, _24581_, _24580_);
  and (_24583_, _24582_, _24579_);
  and (_24584_, _24583_, _24576_);
  nor (_24585_, _24584_, _24333_);
  nor (_24586_, _24585_, _24573_);
  not (_24587_, _24586_);
  and (_24588_, _24587_, _24406_);
  nor (_24589_, _24339_, _21114_);
  nor (_24590_, _24589_, _24588_);
  and (_24591_, _24590_, _24572_);
  and (_24592_, _24591_, _24393_);
  nor (_24593_, _24512_, _24393_);
  nor (_24594_, _24593_, _24592_);
  nor (_24595_, _24470_, _16400_);
  and (_24596_, _24470_, _16031_);
  nor (_24597_, _24596_, _24595_);
  not (_24598_, _24597_);
  and (_24599_, _24598_, _24594_);
  nor (_24600_, _24598_, _24594_);
  nor (_24601_, _24600_, _24599_);
  and (_24602_, _24601_, _24557_);
  and (_24603_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_24604_, _24357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_24605_, _24604_, _24603_);
  and (_24606_, _24362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_24607_, _24355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_24608_, _24607_, _24606_);
  and (_24609_, _24608_, _24605_);
  nor (_24610_, _24609_, _24354_);
  and (_24611_, _24354_, ABINPUT[7]);
  nor (_24612_, _24611_, _24610_);
  not (_24613_, _24612_);
  and (_24614_, _24613_, _24340_);
  not (_24615_, _24614_);
  and (_24616_, _24372_, _22572_);
  not (_24617_, _23127_);
  and (_24618_, _24617_, _22594_);
  nor (_24619_, _24618_, _24616_);
  and (_24620_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_24621_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_24622_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_24623_, _24622_, _24621_);
  and (_24624_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_24625_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_24626_, _24625_, _24624_);
  and (_24627_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_24628_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_24629_, _24628_, _24627_);
  and (_24630_, _24629_, _24626_);
  and (_24631_, _24630_, _24623_);
  nor (_24632_, _24631_, _24333_);
  nor (_24633_, _24632_, _24620_);
  not (_24634_, _24633_);
  and (_24635_, _24634_, _24406_);
  and (_24636_, _23249_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_24637_, _24636_, _23286_);
  not (_24638_, _24637_);
  and (_24639_, _24638_, _24464_);
  nor (_24640_, _24639_, _24635_);
  and (_24641_, _24640_, _24619_);
  and (_24642_, _24641_, _24615_);
  not (_24643_, _24642_);
  and (_24644_, _24643_, _24393_);
  and (_24645_, _24339_, _24372_);
  not (_24646_, _23109_);
  and (_24647_, _24646_, _22594_);
  nor (_24648_, _24647_, _24645_);
  and (_24649_, _24464_, _20236_);
  and (_24650_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_24651_, _24357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_24652_, _24651_, _24650_);
  and (_24653_, _24362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_24654_, _24355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_24655_, _24654_, _24653_);
  and (_24656_, _24655_, _24652_);
  nor (_24657_, _24656_, _24354_);
  and (_24658_, _24354_, ABINPUT[4]);
  nor (_24659_, _24658_, _24657_);
  not (_24660_, _24659_);
  and (_24661_, _24660_, _24340_);
  and (_24662_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_24663_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_24664_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_24665_, _24664_, _24663_);
  and (_24666_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_24667_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_24668_, _24667_, _24666_);
  and (_24669_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_24670_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_24671_, _24670_, _24669_);
  and (_24672_, _24671_, _24668_);
  and (_24673_, _24672_, _24665_);
  nor (_24674_, _24673_, _24333_);
  nor (_24675_, _24674_, _24662_);
  not (_24676_, _24675_);
  and (_24677_, _24676_, _24406_);
  or (_24678_, _24677_, _24661_);
  nor (_24679_, _24678_, _24649_);
  and (_24680_, _24679_, _24648_);
  nor (_24681_, _24680_, _24392_);
  nor (_24682_, _24681_, _24644_);
  and (_24683_, _24470_, _24032_);
  nor (_24684_, _16966_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_24685_, _24684_, _24683_);
  nand (_24686_, _24685_, _24682_);
  or (_24687_, _24685_, _24682_);
  and (_24688_, _24687_, _24686_);
  not (_24689_, _24688_);
  not (_24690_, _24341_);
  and (_24691_, _24553_, _24549_);
  nor (_24692_, _24691_, _24690_);
  and (_24693_, _24692_, _24689_);
  and (_24694_, _24693_, _24602_);
  and (_24695_, _24694_, _24555_);
  not (_24696_, _24469_);
  and (_24697_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_24698_, _24549_);
  and (_24699_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_24700_, _24699_, _24697_);
  and (_24701_, _24700_, _24682_);
  not (_24702_, _24682_);
  and (_24703_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_24704_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_24705_, _24704_, _24703_);
  and (_24706_, _24705_, _24702_);
  or (_24707_, _24706_, _24701_);
  or (_24708_, _24707_, _24696_);
  not (_24709_, _24594_);
  and (_24710_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_24711_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_24712_, _24711_, _24710_);
  and (_24713_, _24712_, _24682_);
  and (_24714_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_24715_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_24716_, _24715_, _24714_);
  and (_24717_, _24716_, _24702_);
  or (_24718_, _24717_, _24713_);
  or (_24719_, _24718_, _24469_);
  and (_24720_, _24719_, _24709_);
  and (_24721_, _24720_, _24708_);
  or (_24722_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_24723_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_24724_, _24723_, _24722_);
  and (_24725_, _24724_, _24682_);
  or (_24726_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_24727_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_24728_, _24727_, _24726_);
  and (_24729_, _24728_, _24702_);
  or (_24730_, _24729_, _24725_);
  or (_24731_, _24730_, _24696_);
  or (_24732_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_24733_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_24734_, _24733_, _24732_);
  and (_24735_, _24734_, _24682_);
  or (_24736_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_24737_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_24738_, _24737_, _24736_);
  and (_24739_, _24738_, _24702_);
  or (_24740_, _24739_, _24735_);
  or (_24741_, _24740_, _24469_);
  and (_24742_, _24741_, _24594_);
  and (_24743_, _24742_, _24731_);
  or (_24744_, _24743_, _24721_);
  or (_24745_, _24744_, _24695_);
  not (_24746_, _24695_);
  or (_24747_, _24746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_24748_, _24747_, _25964_);
  and (_27093_, _24748_, _24745_);
  nor (_24749_, _24552_, _24690_);
  nor (_24750_, _24685_, _24690_);
  and (_24751_, _24750_, _24749_);
  and (_24752_, _24597_, _24341_);
  nor (_24753_, _24473_, _24690_);
  and (_24754_, _24753_, _24752_);
  and (_24755_, _24754_, _24751_);
  or (_24756_, _24755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_24757_, _24755_);
  and (_24758_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_24759_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_24760_, _24759_, _24758_);
  and (_24761_, _24760_, ABINPUT[0]);
  not (_24762_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_24763_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not (_24764_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_24765_, _24764_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_24766_, _24765_, _24763_);
  and (_24767_, _24758_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_24768_, _24767_);
  and (_24769_, _24768_, _24766_);
  or (_24770_, _24769_, _24762_);
  or (_24771_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , ABINPUT[10]);
  and (_24772_, _24771_, _24770_);
  or (_24773_, _24772_, _24761_);
  and (_24774_, _24773_, _24341_);
  or (_24775_, _24774_, _24757_);
  and (_27105_, _24775_, _24756_);
  nor (_24776_, _24753_, _24752_);
  nor (_24777_, _24750_, _24749_);
  and (_24778_, _24777_, _24341_);
  and (_24779_, _24778_, _24776_);
  not (_24780_, _24779_);
  and (_24781_, _24780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  not (_24782_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_24783_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _24782_);
  nor (_24784_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_24785_, _24784_, _24783_);
  and (_24786_, _24785_, ABINPUT[0]);
  and (_24787_, _24762_, ABINPUT[3]);
  or (_24788_, _24787_, _24786_);
  and (_24789_, _24784_, _24782_);
  nor (_24790_, _24789_, _24762_);
  nor (_24791_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_24792_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _24764_);
  nor (_24793_, _24792_, _24791_);
  and (_24794_, _24793_, _24790_);
  or (_24795_, _24794_, _24788_);
  and (_24796_, _24795_, _24341_);
  and (_24797_, _24796_, _24779_);
  or (_27382_, _24797_, _24781_);
  and (_24798_, _24780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_24799_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_24800_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _24764_);
  nor (_24801_, _24800_, _24799_);
  not (_24802_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  nor (_24803_, _24802_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_24804_, _24803_, _24782_);
  nor (_24805_, _24804_, _24762_);
  and (_24806_, _24805_, _24801_);
  and (_24807_, _24803_, _24783_);
  and (_24808_, _24807_, ABINPUT[0]);
  and (_24809_, _24762_, ABINPUT[4]);
  or (_24810_, _24809_, _24808_);
  or (_24811_, _24810_, _24806_);
  and (_24812_, _24811_, _24341_);
  and (_24813_, _24812_, _24779_);
  or (_27388_, _24813_, _24798_);
  and (_24814_, _24780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_24815_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  nor (_24816_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _24764_);
  nor (_24817_, _24816_, _24815_);
  and (_24818_, _24802_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_24819_, _24818_, _24782_);
  nor (_24820_, _24819_, _24762_);
  and (_24821_, _24820_, _24817_);
  and (_24822_, _24783_, _24818_);
  and (_24823_, _24822_, ABINPUT[0]);
  and (_24824_, _24762_, ABINPUT[5]);
  or (_24825_, _24824_, _24823_);
  or (_24826_, _24825_, _24821_);
  and (_24827_, _24826_, _24341_);
  and (_24828_, _24827_, _24779_);
  or (_27394_, _24828_, _24814_);
  and (_24829_, _24780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_24830_, _24783_, _24758_);
  and (_24831_, _24830_, ABINPUT[0]);
  nor (_24832_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_24833_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _24764_);
  nor (_24834_, _24833_, _24832_);
  and (_24835_, _24758_, _24782_);
  not (_24836_, _24835_);
  and (_24837_, _24836_, _24834_);
  or (_24838_, _24837_, _24762_);
  or (_24839_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , ABINPUT[6]);
  and (_24840_, _24839_, _24838_);
  or (_24841_, _24840_, _24831_);
  and (_24842_, _24841_, _24341_);
  and (_24843_, _24842_, _24779_);
  or (_27400_, _24843_, _24829_);
  and (_24844_, _24780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_24845_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_24846_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _24764_);
  nor (_24847_, _24846_, _24845_);
  and (_24848_, _24784_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_24849_, _24848_, _24762_);
  and (_24850_, _24849_, _24847_);
  and (_24851_, _24784_, _24759_);
  and (_24852_, _24851_, ABINPUT[0]);
  and (_24853_, _24762_, ABINPUT[7]);
  or (_24854_, _24853_, _24852_);
  or (_24855_, _24854_, _24850_);
  and (_24856_, _24855_, _24341_);
  and (_24857_, _24856_, _24779_);
  or (_27406_, _24857_, _24844_);
  and (_24858_, _24780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_24859_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_24860_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _24764_);
  nor (_24861_, _24860_, _24859_);
  and (_24862_, _24803_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_24863_, _24862_, _24762_);
  and (_24864_, _24863_, _24861_);
  and (_24865_, _24803_, _24759_);
  and (_24866_, _24865_, ABINPUT[0]);
  and (_24867_, _24762_, ABINPUT[8]);
  or (_24868_, _24867_, _24866_);
  or (_24869_, _24868_, _24864_);
  and (_24870_, _24869_, _24341_);
  and (_24871_, _24870_, _24779_);
  or (_27412_, _24871_, _24858_);
  and (_24872_, _24780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_24873_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_24874_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _24764_);
  nor (_24875_, _24874_, _24873_);
  and (_24876_, _24818_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_24877_, _24876_, _24762_);
  and (_24878_, _24877_, _24875_);
  and (_24879_, _24818_, _24759_);
  and (_24880_, _24879_, ABINPUT[0]);
  and (_24881_, _24762_, ABINPUT[9]);
  or (_24882_, _24881_, _24880_);
  or (_24883_, _24882_, _24878_);
  and (_24884_, _24883_, _24341_);
  and (_24885_, _24884_, _24779_);
  or (_27418_, _24885_, _24872_);
  and (_24886_, _24780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_24887_, _24779_, _24774_);
  or (_27421_, _24887_, _24886_);
  and (_24888_, _24749_, _24685_);
  and (_24889_, _24888_, _24776_);
  or (_24890_, _24889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  not (_24891_, _24889_);
  or (_24892_, _24891_, _24796_);
  and (_27429_, _24892_, _24890_);
  or (_24893_, _24889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_24894_, _24891_, _24812_);
  and (_27433_, _24894_, _24893_);
  or (_24895_, _24889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_24896_, _24891_, _24827_);
  and (_27437_, _24896_, _24895_);
  or (_24897_, _24889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_24898_, _24891_, _24842_);
  and (_27441_, _24898_, _24897_);
  or (_24899_, _24889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_24900_, _24891_, _24856_);
  and (_27445_, _24900_, _24899_);
  or (_24901_, _24889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_24902_, _24891_, _24870_);
  and (_27449_, _24902_, _24901_);
  or (_24903_, _24889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_24904_, _24891_, _24884_);
  and (_27453_, _24904_, _24903_);
  or (_24905_, _24889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_24906_, _24891_, _24774_);
  and (_27456_, _24906_, _24905_);
  and (_24907_, _24750_, _24552_);
  and (_24908_, _24907_, _24776_);
  or (_24909_, _24908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  not (_24910_, _24908_);
  or (_24911_, _24910_, _24796_);
  and (_27464_, _24911_, _24909_);
  or (_24912_, _24908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_24913_, _24910_, _24812_);
  and (_27468_, _24913_, _24912_);
  or (_24914_, _24908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_24915_, _24910_, _24827_);
  and (_27472_, _24915_, _24914_);
  or (_24916_, _24908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_24917_, _24910_, _24842_);
  and (_27476_, _24917_, _24916_);
  or (_24918_, _24908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_24919_, _24910_, _24856_);
  and (_27480_, _24919_, _24918_);
  or (_24920_, _24908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_24921_, _24910_, _24870_);
  and (_27484_, _24921_, _24920_);
  or (_24922_, _24908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_24923_, _24910_, _24884_);
  and (_27488_, _24923_, _24922_);
  or (_24924_, _24908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_24925_, _24910_, _24774_);
  and (_27491_, _24925_, _24924_);
  and (_24926_, _24776_, _24751_);
  or (_24927_, _24926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  not (_24928_, _24926_);
  or (_24929_, _24928_, _24796_);
  and (_27497_, _24929_, _24927_);
  or (_24930_, _24926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_24931_, _24928_, _24812_);
  and (_27501_, _24931_, _24930_);
  or (_24932_, _24926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_24933_, _24928_, _24827_);
  and (_27505_, _24933_, _24932_);
  or (_24934_, _24926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_24935_, _24928_, _24842_);
  and (_27509_, _24935_, _24934_);
  or (_24936_, _24926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_24937_, _24928_, _24856_);
  and (_27513_, _24937_, _24936_);
  or (_24938_, _24926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_24939_, _24928_, _24870_);
  and (_27517_, _24939_, _24938_);
  or (_24940_, _24926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_24941_, _24928_, _24884_);
  and (_27521_, _24941_, _24940_);
  or (_24942_, _24926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_24943_, _24928_, _24774_);
  and (_27524_, _24943_, _24942_);
  and (_24944_, _24753_, _24598_);
  and (_24945_, _24944_, _24777_);
  or (_24946_, _24945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  not (_24947_, _24945_);
  or (_24948_, _24947_, _24796_);
  and (_27532_, _24948_, _24946_);
  or (_24949_, _24945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_24950_, _24947_, _24812_);
  and (_27536_, _24950_, _24949_);
  or (_24951_, _24945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_24952_, _24947_, _24827_);
  and (_27540_, _24952_, _24951_);
  or (_24953_, _24945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_24954_, _24947_, _24842_);
  and (_27544_, _24954_, _24953_);
  or (_24955_, _24945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_24956_, _24947_, _24856_);
  and (_27548_, _24956_, _24955_);
  or (_24957_, _24945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_24958_, _24947_, _24870_);
  and (_27552_, _24958_, _24957_);
  or (_24959_, _24945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_24960_, _24947_, _24884_);
  and (_27556_, _24960_, _24959_);
  or (_24961_, _24945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_24962_, _24947_, _24774_);
  and (_27559_, _24962_, _24961_);
  and (_24963_, _24944_, _24888_);
  or (_24964_, _24963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  not (_24965_, _24963_);
  or (_24966_, _24965_, _24796_);
  and (_27564_, _24966_, _24964_);
  or (_24967_, _24963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_24968_, _24965_, _24812_);
  and (_27568_, _24968_, _24967_);
  or (_24969_, _24963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_24970_, _24965_, _24827_);
  and (_27572_, _24970_, _24969_);
  or (_24971_, _24963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_24972_, _24965_, _24842_);
  and (_27576_, _24972_, _24971_);
  or (_24973_, _24963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_24974_, _24965_, _24856_);
  and (_27580_, _24974_, _24973_);
  or (_24975_, _24963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_24976_, _24965_, _24870_);
  and (_27584_, _24976_, _24975_);
  or (_24977_, _24963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_24978_, _24965_, _24884_);
  and (_27588_, _24978_, _24977_);
  or (_24979_, _24963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_24980_, _24965_, _24774_);
  and (_27591_, _24980_, _24979_);
  and (_24981_, _24944_, _24907_);
  or (_24982_, _24981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  not (_24983_, _24981_);
  or (_24984_, _24983_, _24796_);
  and (_27596_, _24984_, _24982_);
  or (_24985_, _24981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_24986_, _24983_, _24812_);
  and (_27600_, _24986_, _24985_);
  or (_24987_, _24981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_24988_, _24983_, _24827_);
  and (_27604_, _24988_, _24987_);
  or (_24989_, _24981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_24990_, _24983_, _24842_);
  and (_27608_, _24990_, _24989_);
  or (_24991_, _24981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_24992_, _24983_, _24856_);
  and (_27612_, _24992_, _24991_);
  or (_24993_, _24981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_24994_, _24983_, _24870_);
  and (_27616_, _24994_, _24993_);
  or (_24995_, _24981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_24996_, _24983_, _24884_);
  and (_27619_, _24996_, _24995_);
  or (_24997_, _24981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_24998_, _24983_, _24774_);
  and (_27622_, _24998_, _24997_);
  and (_24999_, _24944_, _24751_);
  or (_25000_, _24999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  not (_25001_, _24999_);
  or (_25002_, _25001_, _24796_);
  and (_27627_, _25002_, _25000_);
  or (_25003_, _24999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_25004_, _25001_, _24812_);
  and (_27631_, _25004_, _25003_);
  or (_25005_, _24999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_25006_, _25001_, _24827_);
  and (_27635_, _25006_, _25005_);
  or (_25007_, _24999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_25008_, _25001_, _24842_);
  and (_27639_, _25008_, _25007_);
  or (_25009_, _24999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_25010_, _25001_, _24856_);
  and (_27643_, _25010_, _25009_);
  or (_25011_, _24999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_25012_, _25001_, _24870_);
  and (_27647_, _25012_, _25011_);
  or (_25013_, _24999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_25014_, _25001_, _24884_);
  and (_27651_, _25014_, _25013_);
  or (_25015_, _24999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_25016_, _25001_, _24774_);
  and (_27654_, _25016_, _25015_);
  and (_25017_, _24752_, _24473_);
  and (_25018_, _25017_, _24777_);
  or (_25019_, _25018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  not (_25020_, _25018_);
  or (_25021_, _25020_, _24796_);
  and (_27662_, _25021_, _25019_);
  or (_25022_, _25018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_25023_, _25020_, _24812_);
  and (_27666_, _25023_, _25022_);
  or (_25024_, _25018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_25025_, _25020_, _24827_);
  and (_27670_, _25025_, _25024_);
  or (_25026_, _25018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_25027_, _25020_, _24842_);
  and (_27674_, _25027_, _25026_);
  or (_25028_, _25018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_25029_, _25020_, _24856_);
  and (_27678_, _25029_, _25028_);
  or (_25030_, _25018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_25031_, _25020_, _24870_);
  and (_27682_, _25031_, _25030_);
  or (_25032_, _25018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_25033_, _25020_, _24884_);
  and (_27686_, _25033_, _25032_);
  or (_25034_, _25018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_25035_, _25020_, _24774_);
  and (_27689_, _25035_, _25034_);
  and (_25036_, _25017_, _24888_);
  or (_25037_, _25036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  not (_25038_, _25036_);
  or (_25039_, _25038_, _24796_);
  and (_27694_, _25039_, _25037_);
  or (_25040_, _25036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_25041_, _25038_, _24812_);
  and (_27698_, _25041_, _25040_);
  or (_25042_, _25036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_25043_, _25038_, _24827_);
  and (_27702_, _25043_, _25042_);
  or (_25044_, _25036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_25045_, _25038_, _24842_);
  and (_27706_, _25045_, _25044_);
  or (_25046_, _25036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_25047_, _25038_, _24856_);
  and (_27710_, _25047_, _25046_);
  or (_25048_, _25036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_25049_, _25038_, _24870_);
  and (_27714_, _25049_, _25048_);
  or (_25050_, _25036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_25051_, _25038_, _24884_);
  and (_27718_, _25051_, _25050_);
  or (_25052_, _25036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_25053_, _25038_, _24774_);
  and (_27728_, _25053_, _25052_);
  and (_25054_, _25017_, _24907_);
  or (_25055_, _25054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  not (_25056_, _25054_);
  or (_25057_, _25056_, _24796_);
  and (_27747_, _25057_, _25055_);
  or (_25058_, _25054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_25059_, _25056_, _24812_);
  and (_27763_, _25059_, _25058_);
  or (_25060_, _25054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_25061_, _25056_, _24827_);
  and (_27776_, _25061_, _25060_);
  or (_25062_, _25054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_25063_, _25056_, _24842_);
  and (_27794_, _25063_, _25062_);
  or (_25064_, _25054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_25065_, _25056_, _24856_);
  and (_27805_, _25065_, _25064_);
  or (_25066_, _25054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_25067_, _25056_, _24870_);
  and (_27822_, _25067_, _25066_);
  or (_25068_, _25054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_25069_, _25056_, _24884_);
  and (_27841_, _25069_, _25068_);
  or (_25070_, _25054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_25071_, _25056_, _24774_);
  and (_27851_, _25071_, _25070_);
  and (_25072_, _25017_, _24751_);
  or (_25073_, _25072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  not (_25074_, _25072_);
  or (_25075_, _25074_, _24796_);
  and (_27877_, _25075_, _25073_);
  or (_25076_, _25072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_25077_, _25074_, _24812_);
  and (_27895_, _25077_, _25076_);
  or (_25078_, _25072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_25079_, _25074_, _24827_);
  and (_27913_, _25079_, _25078_);
  or (_25080_, _25072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_25081_, _25074_, _24842_);
  and (_27934_, _25081_, _25080_);
  or (_25082_, _25072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_25083_, _25074_, _24856_);
  and (_27954_, _25083_, _25082_);
  or (_25084_, _25072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_25085_, _25074_, _24870_);
  and (_27968_, _25085_, _25084_);
  or (_25086_, _25072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_25087_, _25074_, _24884_);
  and (_27972_, _25087_, _25086_);
  or (_25088_, _25072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_25089_, _25074_, _24774_);
  and (_27975_, _25089_, _25088_);
  and (_25090_, _24777_, _24754_);
  or (_25091_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  not (_25092_, _25090_);
  or (_25093_, _25092_, _24796_);
  and (_27981_, _25093_, _25091_);
  or (_25094_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_25095_, _25092_, _24812_);
  and (_27985_, _25095_, _25094_);
  or (_25096_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_25097_, _25092_, _24827_);
  and (_27989_, _25097_, _25096_);
  or (_25098_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_25099_, _25092_, _24842_);
  and (_27993_, _25099_, _25098_);
  or (_25100_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_25101_, _25092_, _24856_);
  and (_27997_, _25101_, _25100_);
  or (_25102_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_25103_, _25092_, _24870_);
  and (_28001_, _25103_, _25102_);
  or (_25104_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_25105_, _25092_, _24884_);
  and (_28005_, _25105_, _25104_);
  or (_25106_, _25090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_25107_, _25092_, _24774_);
  and (_28008_, _25107_, _25106_);
  and (_25108_, _24888_, _24754_);
  or (_25109_, _25108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  not (_25110_, _25108_);
  or (_25111_, _25110_, _24796_);
  and (_28013_, _25111_, _25109_);
  or (_25112_, _25108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_25113_, _25110_, _24812_);
  and (_28017_, _25113_, _25112_);
  or (_25114_, _25108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_25115_, _25110_, _24827_);
  and (_28021_, _25115_, _25114_);
  or (_25116_, _25108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_25117_, _25110_, _24842_);
  and (_28025_, _25117_, _25116_);
  or (_25118_, _25108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_25119_, _25110_, _24856_);
  and (_28029_, _25119_, _25118_);
  or (_25120_, _25108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_25121_, _25110_, _24870_);
  and (_28033_, _25121_, _25120_);
  or (_25122_, _25108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_25123_, _25110_, _24884_);
  and (_28037_, _25123_, _25122_);
  or (_25124_, _25108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_25126_, _25110_, _24774_);
  and (_28040_, _25126_, _25124_);
  and (_25127_, _24907_, _24754_);
  or (_25128_, _25127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  not (_25129_, _25127_);
  or (_25130_, _25129_, _24796_);
  and (_28045_, _25130_, _25128_);
  or (_25131_, _25127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_25132_, _25129_, _24812_);
  and (_28049_, _25132_, _25131_);
  or (_25134_, _25127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_25135_, _25129_, _24827_);
  and (_28053_, _25135_, _25134_);
  or (_25136_, _25127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_25137_, _25129_, _24842_);
  and (_28057_, _25137_, _25136_);
  or (_25138_, _25127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_25139_, _25129_, _24856_);
  and (_28061_, _25139_, _25138_);
  or (_25140_, _25127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_25142_, _25129_, _24870_);
  and (_28065_, _25142_, _25140_);
  or (_25143_, _25127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_25144_, _25129_, _24884_);
  and (_28069_, _25144_, _25143_);
  or (_25145_, _25127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_25146_, _25129_, _24774_);
  and (_28072_, _25146_, _25145_);
  or (_25147_, _24755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_25148_, _24796_, _24757_);
  and (_28077_, _25148_, _25147_);
  or (_25150_, _24755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_25151_, _24812_, _24757_);
  and (_28081_, _25151_, _25150_);
  or (_25152_, _24755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_25153_, _24827_, _24757_);
  and (_28085_, _25153_, _25152_);
  or (_25154_, _24755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_25155_, _24842_, _24757_);
  and (_28089_, _25155_, _25154_);
  or (_25157_, _24755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_25158_, _24856_, _24757_);
  and (_28093_, _25158_, _25157_);
  or (_25159_, _24755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_25160_, _24870_, _24757_);
  and (_28097_, _25160_, _25159_);
  or (_25161_, _24755_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_25162_, _24884_, _24757_);
  and (_28101_, _25162_, _25161_);
  and (_25163_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_25165_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_25166_, _25165_, _25163_);
  and (_25167_, _25166_, _24682_);
  and (_25168_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_25169_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_25170_, _25169_, _25168_);
  and (_25171_, _25170_, _24702_);
  or (_25172_, _25171_, _25167_);
  or (_25173_, _25172_, _24696_);
  and (_25174_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_25176_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_25177_, _25176_, _25174_);
  and (_25178_, _25177_, _24682_);
  and (_25179_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_25180_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_25181_, _25180_, _25179_);
  and (_25182_, _25181_, _24702_);
  or (_25183_, _25182_, _25178_);
  or (_25184_, _25183_, _24469_);
  and (_25185_, _25184_, _24709_);
  and (_25186_, _25185_, _25173_);
  or (_25187_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_25188_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_25189_, _25188_, _25187_);
  and (_25190_, _25189_, _24682_);
  or (_25191_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_25192_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_25193_, _25192_, _25191_);
  and (_25194_, _25193_, _24702_);
  or (_25195_, _25194_, _25190_);
  or (_25196_, _25195_, _24696_);
  or (_25197_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_25198_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_25199_, _25198_, _25197_);
  and (_25200_, _25199_, _24682_);
  or (_25201_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_25202_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_25203_, _25202_, _25201_);
  and (_25204_, _25203_, _24702_);
  or (_25205_, _25204_, _25200_);
  or (_25206_, _25205_, _24469_);
  and (_25207_, _25206_, _24594_);
  and (_25208_, _25207_, _25196_);
  or (_25209_, _25208_, _25186_);
  or (_25210_, _25209_, _24695_);
  or (_25211_, _24746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_25212_, _25211_, _25964_);
  and (_00046_, _25212_, _25210_);
  and (_25213_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_25214_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_25215_, _25214_, _25213_);
  and (_25216_, _25215_, _24682_);
  and (_25217_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_25218_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_25219_, _25218_, _25217_);
  and (_25220_, _25219_, _24702_);
  or (_25221_, _25220_, _25216_);
  or (_25222_, _25221_, _24696_);
  and (_25223_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_25224_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_25225_, _25224_, _25223_);
  and (_25226_, _25225_, _24682_);
  and (_25227_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_25228_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_25229_, _25228_, _25227_);
  and (_25230_, _25229_, _24702_);
  or (_25231_, _25230_, _25226_);
  or (_25232_, _25231_, _24469_);
  and (_25233_, _25232_, _24709_);
  and (_25234_, _25233_, _25222_);
  or (_25235_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_25236_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_25237_, _25236_, _25235_);
  and (_25238_, _25237_, _24682_);
  or (_25239_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_25240_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_25241_, _25240_, _25239_);
  and (_25242_, _25241_, _24702_);
  or (_25243_, _25242_, _25238_);
  or (_25244_, _25243_, _24696_);
  or (_25245_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_25246_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_25247_, _25246_, _25245_);
  and (_25248_, _25247_, _24682_);
  or (_25249_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_25250_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_25251_, _25250_, _25249_);
  and (_25252_, _25251_, _24702_);
  or (_25253_, _25252_, _25248_);
  or (_25254_, _25253_, _24469_);
  and (_25255_, _25254_, _24594_);
  and (_25256_, _25255_, _25244_);
  or (_25257_, _25256_, _25234_);
  or (_25258_, _25257_, _24695_);
  or (_25259_, _24746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_25260_, _25259_, _25964_);
  and (_00048_, _25260_, _25258_);
  and (_25261_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_25262_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_25263_, _25262_, _25261_);
  and (_25264_, _25263_, _24682_);
  and (_25265_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  and (_25266_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_25267_, _25266_, _25265_);
  and (_25268_, _25267_, _24702_);
  or (_25269_, _25268_, _25264_);
  or (_25270_, _25269_, _24696_);
  and (_25271_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_25272_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_25273_, _25272_, _25271_);
  and (_25274_, _25273_, _24682_);
  and (_25275_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_25276_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_25277_, _25276_, _25275_);
  and (_25278_, _25277_, _24702_);
  or (_25279_, _25278_, _25274_);
  or (_25280_, _25279_, _24469_);
  and (_25281_, _25280_, _24709_);
  and (_25282_, _25281_, _25270_);
  or (_25283_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_25284_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_25285_, _25284_, _25283_);
  and (_25286_, _25285_, _24682_);
  or (_25287_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_25288_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_25289_, _25288_, _25287_);
  and (_25290_, _25289_, _24702_);
  or (_25291_, _25290_, _25286_);
  or (_25292_, _25291_, _24696_);
  or (_25293_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_25294_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_25295_, _25294_, _25293_);
  and (_25296_, _25295_, _24682_);
  or (_25297_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_25298_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_25299_, _25298_, _25297_);
  and (_25300_, _25299_, _24702_);
  or (_25301_, _25300_, _25296_);
  or (_25302_, _25301_, _24469_);
  and (_25305_, _25302_, _24594_);
  and (_25308_, _25305_, _25292_);
  or (_25311_, _25308_, _25282_);
  or (_25316_, _25311_, _24695_);
  or (_25319_, _24746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_25321_, _25319_, _25964_);
  and (_00050_, _25321_, _25316_);
  and (_25327_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_25329_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_25332_, _25329_, _25327_);
  and (_25337_, _25332_, _24682_);
  and (_25339_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_25340_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_25341_, _25340_, _25339_);
  and (_25342_, _25341_, _24702_);
  or (_25343_, _25342_, _25337_);
  or (_25344_, _25343_, _24696_);
  and (_25345_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_25346_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_25347_, _25346_, _25345_);
  and (_25348_, _25347_, _24682_);
  and (_25349_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_25350_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_25351_, _25350_, _25349_);
  and (_25352_, _25351_, _24702_);
  or (_25353_, _25352_, _25348_);
  or (_25354_, _25353_, _24469_);
  and (_25355_, _25354_, _24709_);
  and (_25356_, _25355_, _25344_);
  or (_25357_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_25358_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_25359_, _25358_, _25357_);
  and (_25360_, _25359_, _24682_);
  or (_25361_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_25362_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_25363_, _25362_, _25361_);
  and (_25364_, _25363_, _24702_);
  or (_25365_, _25364_, _25360_);
  or (_25366_, _25365_, _24696_);
  or (_25367_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_25368_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_25369_, _25368_, _25367_);
  and (_25370_, _25369_, _24682_);
  or (_25371_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_25372_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_25373_, _25372_, _25371_);
  and (_25374_, _25373_, _24702_);
  or (_25375_, _25374_, _25370_);
  or (_25376_, _25375_, _24469_);
  and (_25377_, _25376_, _24594_);
  and (_25378_, _25377_, _25366_);
  or (_25379_, _25378_, _25356_);
  or (_25380_, _25379_, _24695_);
  or (_25381_, _24746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_25382_, _25381_, _25964_);
  and (_00052_, _25382_, _25380_);
  and (_25383_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_25384_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_25385_, _25384_, _25383_);
  and (_25386_, _25385_, _24682_);
  and (_25387_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_25388_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_25389_, _25388_, _25387_);
  and (_25390_, _25389_, _24702_);
  or (_25392_, _25390_, _25386_);
  or (_25394_, _25392_, _24696_);
  and (_25396_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_25398_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_25400_, _25398_, _25396_);
  and (_25402_, _25400_, _24682_);
  and (_25404_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_25406_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_25408_, _25406_, _25404_);
  and (_25410_, _25408_, _24702_);
  or (_25412_, _25410_, _25402_);
  or (_25414_, _25412_, _24469_);
  and (_25416_, _25414_, _24709_);
  and (_25418_, _25416_, _25394_);
  or (_25420_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_25422_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_25424_, _25422_, _25420_);
  and (_25426_, _25424_, _24682_);
  or (_25428_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_25430_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_25432_, _25430_, _25428_);
  and (_25434_, _25432_, _24702_);
  or (_25436_, _25434_, _25426_);
  or (_25438_, _25436_, _24696_);
  or (_25440_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_25442_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_25444_, _25442_, _25440_);
  and (_25446_, _25444_, _24682_);
  or (_25447_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_25448_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_25449_, _25448_, _25447_);
  and (_25450_, _25449_, _24702_);
  or (_25451_, _25450_, _25446_);
  or (_25452_, _25451_, _24469_);
  and (_25453_, _25452_, _24594_);
  and (_25454_, _25453_, _25438_);
  or (_25455_, _25454_, _25418_);
  or (_25456_, _25455_, _24695_);
  or (_25457_, _24746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_25458_, _25457_, _25964_);
  and (_00054_, _25458_, _25456_);
  and (_25459_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_25460_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_25461_, _25460_, _25459_);
  and (_25462_, _25461_, _24682_);
  and (_25463_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_25464_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_25465_, _25464_, _25463_);
  and (_25466_, _25465_, _24702_);
  or (_25467_, _25466_, _25462_);
  or (_25468_, _25467_, _24696_);
  and (_25469_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_25470_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_25471_, _25470_, _25469_);
  and (_25472_, _25471_, _24682_);
  and (_25473_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_25474_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_25475_, _25474_, _25473_);
  and (_25476_, _25475_, _24702_);
  or (_25477_, _25476_, _25472_);
  or (_25478_, _25477_, _24469_);
  and (_25479_, _25478_, _24709_);
  and (_25480_, _25479_, _25468_);
  or (_25481_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_25482_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_25483_, _25482_, _25481_);
  and (_25484_, _25483_, _24682_);
  or (_25485_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_25486_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_25487_, _25486_, _25485_);
  and (_25488_, _25487_, _24702_);
  or (_25489_, _25488_, _25484_);
  or (_25490_, _25489_, _24696_);
  or (_25491_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_25492_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_25493_, _25492_, _25491_);
  and (_25494_, _25493_, _24682_);
  or (_25495_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_25496_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_25497_, _25496_, _25495_);
  and (_25498_, _25497_, _24702_);
  or (_25499_, _25498_, _25494_);
  or (_25500_, _25499_, _24469_);
  and (_25501_, _25500_, _24594_);
  and (_25502_, _25501_, _25490_);
  or (_25503_, _25502_, _25480_);
  or (_25504_, _25503_, _24695_);
  or (_25505_, _24746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_25506_, _25505_, _25964_);
  and (_00056_, _25506_, _25504_);
  and (_25507_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_25508_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_25509_, _25508_, _25507_);
  and (_25510_, _25509_, _24682_);
  and (_25511_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_25512_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_25513_, _25512_, _25511_);
  and (_25514_, _25513_, _24702_);
  or (_25515_, _25514_, _25510_);
  or (_25516_, _25515_, _24696_);
  and (_25517_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_25518_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_25519_, _25518_, _25517_);
  and (_25520_, _25519_, _24682_);
  and (_25521_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_25522_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_25523_, _25522_, _25521_);
  and (_25524_, _25523_, _24702_);
  or (_25525_, _25524_, _25520_);
  or (_25526_, _25525_, _24469_);
  and (_25527_, _25526_, _24709_);
  and (_25528_, _25527_, _25516_);
  or (_25529_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_25530_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_25531_, _25530_, _25529_);
  and (_25532_, _25531_, _24682_);
  or (_25533_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_25534_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_25535_, _25534_, _25533_);
  and (_25536_, _25535_, _24702_);
  or (_25537_, _25536_, _25532_);
  or (_25538_, _25537_, _24696_);
  or (_25539_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_25540_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_25541_, _25540_, _25539_);
  and (_25542_, _25541_, _24682_);
  or (_25543_, _24549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_25544_, _24698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_25545_, _25544_, _25543_);
  and (_25546_, _25545_, _24702_);
  or (_25547_, _25546_, _25542_);
  or (_25548_, _25547_, _24469_);
  and (_25549_, _25548_, _24594_);
  and (_25550_, _25549_, _25538_);
  or (_25551_, _25550_, _25528_);
  or (_25552_, _25551_, _24695_);
  or (_25553_, _24746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_25554_, _25553_, _25964_);
  and (_00058_, _25554_, _25552_);
  or (_25555_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_25556_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_25557_, _25556_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_25558_, _25557_, _25555_);
  nand (_25559_, _25558_, _25964_);
  or (_25560_, \oc8051_gm_cxrom_1.cell0.data [7], _25964_);
  and (_00066_, _25560_, _25559_);
  or (_25561_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_25562_, \oc8051_gm_cxrom_1.cell0.data [0], _25556_);
  nand (_25563_, _25562_, _25561_);
  nand (_25564_, _25563_, _25964_);
  or (_25565_, \oc8051_gm_cxrom_1.cell0.data [0], _25964_);
  and (_00098_, _25565_, _25564_);
  or (_25566_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_25567_, \oc8051_gm_cxrom_1.cell0.data [1], _25556_);
  nand (_25568_, _25567_, _25566_);
  nand (_25569_, _25568_, _25964_);
  or (_25570_, \oc8051_gm_cxrom_1.cell0.data [1], _25964_);
  and (_00100_, _25570_, _25569_);
  or (_25571_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_25572_, \oc8051_gm_cxrom_1.cell0.data [2], _25556_);
  nand (_25575_, _25572_, _25571_);
  nand (_25576_, _25575_, _25964_);
  or (_25577_, \oc8051_gm_cxrom_1.cell0.data [2], _25964_);
  and (_00102_, _25577_, _25576_);
  or (_25578_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_25579_, \oc8051_gm_cxrom_1.cell0.data [3], _25556_);
  nand (_25580_, _25579_, _25578_);
  nand (_25581_, _25580_, _25964_);
  or (_25582_, \oc8051_gm_cxrom_1.cell0.data [3], _25964_);
  and (_00104_, _25582_, _25581_);
  or (_25583_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_25584_, \oc8051_gm_cxrom_1.cell0.data [4], _25556_);
  nand (_25585_, _25584_, _25583_);
  nand (_25586_, _25585_, _25964_);
  or (_25587_, \oc8051_gm_cxrom_1.cell0.data [4], _25964_);
  and (_00106_, _25587_, _25586_);
  or (_25588_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_25589_, \oc8051_gm_cxrom_1.cell0.data [5], _25556_);
  nand (_25590_, _25589_, _25588_);
  nand (_25591_, _25590_, _25964_);
  or (_25592_, \oc8051_gm_cxrom_1.cell0.data [5], _25964_);
  and (_00108_, _25592_, _25591_);
  or (_25593_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_25594_, \oc8051_gm_cxrom_1.cell0.data [6], _25556_);
  nand (_25595_, _25594_, _25593_);
  nand (_25596_, _25595_, _25964_);
  or (_25597_, \oc8051_gm_cxrom_1.cell0.data [6], _25964_);
  and (_00110_, _25597_, _25596_);
  or (_25598_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_25599_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_25600_, _25599_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_25601_, _25600_, _25598_);
  nand (_25602_, _25601_, _25964_);
  or (_25603_, \oc8051_gm_cxrom_1.cell1.data [7], _25964_);
  and (_00117_, _25603_, _25602_);
  or (_25604_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_25605_, \oc8051_gm_cxrom_1.cell1.data [0], _25599_);
  nand (_25606_, _25605_, _25604_);
  nand (_25607_, _25606_, _25964_);
  or (_25608_, \oc8051_gm_cxrom_1.cell1.data [0], _25964_);
  and (_00149_, _25608_, _25607_);
  or (_25609_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_25610_, \oc8051_gm_cxrom_1.cell1.data [1], _25599_);
  nand (_25611_, _25610_, _25609_);
  nand (_25612_, _25611_, _25964_);
  or (_25613_, \oc8051_gm_cxrom_1.cell1.data [1], _25964_);
  and (_00151_, _25613_, _25612_);
  or (_25614_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_25615_, \oc8051_gm_cxrom_1.cell1.data [2], _25599_);
  nand (_25616_, _25615_, _25614_);
  nand (_25617_, _25616_, _25964_);
  or (_25618_, \oc8051_gm_cxrom_1.cell1.data [2], _25964_);
  and (_00153_, _25618_, _25617_);
  or (_25619_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_25620_, \oc8051_gm_cxrom_1.cell1.data [3], _25599_);
  nand (_25621_, _25620_, _25619_);
  nand (_25622_, _25621_, _25964_);
  or (_25623_, \oc8051_gm_cxrom_1.cell1.data [3], _25964_);
  and (_00155_, _25623_, _25622_);
  or (_25624_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_25625_, \oc8051_gm_cxrom_1.cell1.data [4], _25599_);
  nand (_25626_, _25625_, _25624_);
  nand (_25627_, _25626_, _25964_);
  or (_25628_, \oc8051_gm_cxrom_1.cell1.data [4], _25964_);
  and (_00157_, _25628_, _25627_);
  or (_25629_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_25630_, \oc8051_gm_cxrom_1.cell1.data [5], _25599_);
  nand (_25631_, _25630_, _25629_);
  nand (_25632_, _25631_, _25964_);
  or (_25633_, \oc8051_gm_cxrom_1.cell1.data [5], _25964_);
  and (_00159_, _25633_, _25632_);
  or (_25634_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_25635_, \oc8051_gm_cxrom_1.cell1.data [6], _25599_);
  nand (_25636_, _25635_, _25634_);
  nand (_25637_, _25636_, _25964_);
  or (_25638_, \oc8051_gm_cxrom_1.cell1.data [6], _25964_);
  and (_00161_, _25638_, _25637_);
  or (_25639_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_25640_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_25641_, _25640_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_25642_, _25641_, _25639_);
  nand (_25643_, _25642_, _25964_);
  or (_25644_, \oc8051_gm_cxrom_1.cell2.data [7], _25964_);
  and (_00169_, _25644_, _25643_);
  or (_25645_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_25646_, \oc8051_gm_cxrom_1.cell2.data [0], _25640_);
  nand (_25647_, _25646_, _25645_);
  nand (_25648_, _25647_, _25964_);
  or (_25649_, \oc8051_gm_cxrom_1.cell2.data [0], _25964_);
  and (_00201_, _25649_, _25648_);
  or (_25650_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_25651_, \oc8051_gm_cxrom_1.cell2.data [1], _25640_);
  nand (_25652_, _25651_, _25650_);
  nand (_25653_, _25652_, _25964_);
  or (_25654_, \oc8051_gm_cxrom_1.cell2.data [1], _25964_);
  and (_00203_, _25654_, _25653_);
  or (_25655_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_25656_, \oc8051_gm_cxrom_1.cell2.data [2], _25640_);
  nand (_25657_, _25656_, _25655_);
  nand (_25658_, _25657_, _25964_);
  or (_25659_, \oc8051_gm_cxrom_1.cell2.data [2], _25964_);
  and (_00205_, _25659_, _25658_);
  or (_25660_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_25661_, \oc8051_gm_cxrom_1.cell2.data [3], _25640_);
  nand (_25662_, _25661_, _25660_);
  nand (_25663_, _25662_, _25964_);
  or (_25664_, \oc8051_gm_cxrom_1.cell2.data [3], _25964_);
  and (_00207_, _25664_, _25663_);
  or (_25665_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_25666_, \oc8051_gm_cxrom_1.cell2.data [4], _25640_);
  nand (_25667_, _25666_, _25665_);
  nand (_25668_, _25667_, _25964_);
  or (_25669_, \oc8051_gm_cxrom_1.cell2.data [4], _25964_);
  and (_00209_, _25669_, _25668_);
  or (_25670_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_25671_, \oc8051_gm_cxrom_1.cell2.data [5], _25640_);
  nand (_25672_, _25671_, _25670_);
  nand (_25673_, _25672_, _25964_);
  or (_25674_, \oc8051_gm_cxrom_1.cell2.data [5], _25964_);
  and (_00211_, _25674_, _25673_);
  or (_25675_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_25676_, \oc8051_gm_cxrom_1.cell2.data [6], _25640_);
  nand (_25677_, _25676_, _25675_);
  nand (_25678_, _25677_, _25964_);
  or (_25679_, \oc8051_gm_cxrom_1.cell2.data [6], _25964_);
  and (_00213_, _25679_, _25678_);
  or (_25680_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_25681_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_25682_, _25681_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_25683_, _25682_, _25680_);
  nand (_25684_, _25683_, _25964_);
  or (_25685_, \oc8051_gm_cxrom_1.cell3.data [7], _25964_);
  and (_00221_, _25685_, _25684_);
  or (_25686_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_25687_, \oc8051_gm_cxrom_1.cell3.data [0], _25681_);
  nand (_25688_, _25687_, _25686_);
  nand (_25689_, _25688_, _25964_);
  or (_25690_, \oc8051_gm_cxrom_1.cell3.data [0], _25964_);
  and (_00253_, _25690_, _25689_);
  or (_25691_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_25692_, \oc8051_gm_cxrom_1.cell3.data [1], _25681_);
  nand (_25693_, _25692_, _25691_);
  nand (_25694_, _25693_, _25964_);
  or (_25695_, \oc8051_gm_cxrom_1.cell3.data [1], _25964_);
  and (_00255_, _25695_, _25694_);
  or (_25696_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_25697_, \oc8051_gm_cxrom_1.cell3.data [2], _25681_);
  nand (_25698_, _25697_, _25696_);
  nand (_25699_, _25698_, _25964_);
  or (_25700_, \oc8051_gm_cxrom_1.cell3.data [2], _25964_);
  and (_00257_, _25700_, _25699_);
  or (_25701_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_25702_, \oc8051_gm_cxrom_1.cell3.data [3], _25681_);
  nand (_25703_, _25702_, _25701_);
  nand (_25704_, _25703_, _25964_);
  or (_25705_, \oc8051_gm_cxrom_1.cell3.data [3], _25964_);
  and (_00259_, _25705_, _25704_);
  or (_25706_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_25707_, \oc8051_gm_cxrom_1.cell3.data [4], _25681_);
  nand (_25708_, _25707_, _25706_);
  nand (_25709_, _25708_, _25964_);
  or (_25710_, \oc8051_gm_cxrom_1.cell3.data [4], _25964_);
  and (_00261_, _25710_, _25709_);
  or (_25711_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_25712_, \oc8051_gm_cxrom_1.cell3.data [5], _25681_);
  nand (_25713_, _25712_, _25711_);
  nand (_25714_, _25713_, _25964_);
  or (_25715_, \oc8051_gm_cxrom_1.cell3.data [5], _25964_);
  and (_00263_, _25715_, _25714_);
  or (_25716_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_25717_, \oc8051_gm_cxrom_1.cell3.data [6], _25681_);
  nand (_25718_, _25717_, _25716_);
  nand (_25719_, _25718_, _25964_);
  or (_25720_, \oc8051_gm_cxrom_1.cell3.data [6], _25964_);
  and (_00265_, _25720_, _25719_);
  or (_25721_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_25722_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_25723_, _25722_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_25724_, _25723_, _25721_);
  nand (_25725_, _25724_, _25964_);
  or (_25726_, \oc8051_gm_cxrom_1.cell4.data [7], _25964_);
  and (_00273_, _25726_, _25725_);
  or (_25727_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_25728_, \oc8051_gm_cxrom_1.cell4.data [0], _25722_);
  nand (_25729_, _25728_, _25727_);
  nand (_25730_, _25729_, _25964_);
  or (_25731_, \oc8051_gm_cxrom_1.cell4.data [0], _25964_);
  and (_00305_, _25731_, _25730_);
  or (_25732_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_25733_, \oc8051_gm_cxrom_1.cell4.data [1], _25722_);
  nand (_25734_, _25733_, _25732_);
  nand (_25735_, _25734_, _25964_);
  or (_25736_, \oc8051_gm_cxrom_1.cell4.data [1], _25964_);
  and (_00307_, _25736_, _25735_);
  or (_25737_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_25738_, \oc8051_gm_cxrom_1.cell4.data [2], _25722_);
  nand (_25739_, _25738_, _25737_);
  nand (_25740_, _25739_, _25964_);
  or (_25741_, \oc8051_gm_cxrom_1.cell4.data [2], _25964_);
  and (_00309_, _25741_, _25740_);
  or (_25742_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_25743_, \oc8051_gm_cxrom_1.cell4.data [3], _25722_);
  nand (_25744_, _25743_, _25742_);
  nand (_25745_, _25744_, _25964_);
  or (_25746_, \oc8051_gm_cxrom_1.cell4.data [3], _25964_);
  and (_00311_, _25746_, _25745_);
  or (_25747_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_25748_, \oc8051_gm_cxrom_1.cell4.data [4], _25722_);
  nand (_25749_, _25748_, _25747_);
  nand (_25750_, _25749_, _25964_);
  or (_25751_, \oc8051_gm_cxrom_1.cell4.data [4], _25964_);
  and (_00313_, _25751_, _25750_);
  or (_25752_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_25753_, \oc8051_gm_cxrom_1.cell4.data [5], _25722_);
  nand (_25754_, _25753_, _25752_);
  nand (_25755_, _25754_, _25964_);
  or (_25756_, \oc8051_gm_cxrom_1.cell4.data [5], _25964_);
  and (_00315_, _25756_, _25755_);
  or (_25757_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_25758_, \oc8051_gm_cxrom_1.cell4.data [6], _25722_);
  nand (_25759_, _25758_, _25757_);
  nand (_25760_, _25759_, _25964_);
  or (_25761_, \oc8051_gm_cxrom_1.cell4.data [6], _25964_);
  and (_00317_, _25761_, _25760_);
  or (_25762_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_25763_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_25764_, _25763_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_25765_, _25764_, _25762_);
  nand (_25766_, _25765_, _25964_);
  or (_25767_, \oc8051_gm_cxrom_1.cell5.data [7], _25964_);
  and (_00325_, _25767_, _25766_);
  or (_25768_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_25769_, \oc8051_gm_cxrom_1.cell5.data [0], _25763_);
  nand (_25770_, _25769_, _25768_);
  nand (_25771_, _25770_, _25964_);
  or (_25772_, \oc8051_gm_cxrom_1.cell5.data [0], _25964_);
  and (_00357_, _25772_, _25771_);
  or (_25773_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_25774_, \oc8051_gm_cxrom_1.cell5.data [1], _25763_);
  nand (_25775_, _25774_, _25773_);
  nand (_25776_, _25775_, _25964_);
  or (_25777_, \oc8051_gm_cxrom_1.cell5.data [1], _25964_);
  and (_00359_, _25777_, _25776_);
  or (_25778_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_25779_, \oc8051_gm_cxrom_1.cell5.data [2], _25763_);
  nand (_25780_, _25779_, _25778_);
  nand (_25781_, _25780_, _25964_);
  or (_25782_, \oc8051_gm_cxrom_1.cell5.data [2], _25964_);
  and (_00361_, _25782_, _25781_);
  or (_25783_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_25784_, \oc8051_gm_cxrom_1.cell5.data [3], _25763_);
  nand (_25785_, _25784_, _25783_);
  nand (_25786_, _25785_, _25964_);
  or (_25787_, \oc8051_gm_cxrom_1.cell5.data [3], _25964_);
  and (_00363_, _25787_, _25786_);
  or (_25788_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_25789_, \oc8051_gm_cxrom_1.cell5.data [4], _25763_);
  nand (_25790_, _25789_, _25788_);
  nand (_25791_, _25790_, _25964_);
  or (_25792_, \oc8051_gm_cxrom_1.cell5.data [4], _25964_);
  and (_00365_, _25792_, _25791_);
  or (_25793_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_25794_, \oc8051_gm_cxrom_1.cell5.data [5], _25763_);
  nand (_25795_, _25794_, _25793_);
  nand (_25796_, _25795_, _25964_);
  or (_25797_, \oc8051_gm_cxrom_1.cell5.data [5], _25964_);
  and (_00367_, _25797_, _25796_);
  or (_25798_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_25799_, \oc8051_gm_cxrom_1.cell5.data [6], _25763_);
  nand (_25800_, _25799_, _25798_);
  nand (_25801_, _25800_, _25964_);
  or (_25802_, \oc8051_gm_cxrom_1.cell5.data [6], _25964_);
  and (_00369_, _25802_, _25801_);
  or (_25803_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_25804_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_25805_, _25804_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_25806_, _25805_, _25803_);
  nand (_25807_, _25806_, _25964_);
  or (_25808_, \oc8051_gm_cxrom_1.cell6.data [7], _25964_);
  and (_00377_, _25808_, _25807_);
  or (_25809_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_25810_, \oc8051_gm_cxrom_1.cell6.data [0], _25804_);
  nand (_25811_, _25810_, _25809_);
  nand (_25812_, _25811_, _25964_);
  or (_25813_, \oc8051_gm_cxrom_1.cell6.data [0], _25964_);
  and (_00409_, _25813_, _25812_);
  or (_25814_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_25815_, \oc8051_gm_cxrom_1.cell6.data [1], _25804_);
  nand (_25816_, _25815_, _25814_);
  nand (_25817_, _25816_, _25964_);
  or (_25818_, \oc8051_gm_cxrom_1.cell6.data [1], _25964_);
  and (_00411_, _25818_, _25817_);
  or (_25819_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_25820_, \oc8051_gm_cxrom_1.cell6.data [2], _25804_);
  nand (_25821_, _25820_, _25819_);
  nand (_25822_, _25821_, _25964_);
  or (_25823_, \oc8051_gm_cxrom_1.cell6.data [2], _25964_);
  and (_00413_, _25823_, _25822_);
  or (_25824_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_25825_, \oc8051_gm_cxrom_1.cell6.data [3], _25804_);
  nand (_25826_, _25825_, _25824_);
  nand (_25827_, _25826_, _25964_);
  or (_25828_, \oc8051_gm_cxrom_1.cell6.data [3], _25964_);
  and (_00415_, _25828_, _25827_);
  or (_25829_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_25830_, \oc8051_gm_cxrom_1.cell6.data [4], _25804_);
  nand (_25831_, _25830_, _25829_);
  nand (_25832_, _25831_, _25964_);
  or (_25833_, \oc8051_gm_cxrom_1.cell6.data [4], _25964_);
  and (_00417_, _25833_, _25832_);
  or (_25834_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_25835_, \oc8051_gm_cxrom_1.cell6.data [5], _25804_);
  nand (_25836_, _25835_, _25834_);
  nand (_25837_, _25836_, _25964_);
  or (_25838_, \oc8051_gm_cxrom_1.cell6.data [5], _25964_);
  and (_00419_, _25838_, _25837_);
  or (_25839_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_25840_, \oc8051_gm_cxrom_1.cell6.data [6], _25804_);
  nand (_25841_, _25840_, _25839_);
  nand (_25842_, _25841_, _25964_);
  or (_25843_, \oc8051_gm_cxrom_1.cell6.data [6], _25964_);
  and (_00421_, _25843_, _25842_);
  or (_25844_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_25845_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_25846_, _25845_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_25847_, _25846_, _25844_);
  nand (_25848_, _25847_, _25964_);
  or (_25849_, \oc8051_gm_cxrom_1.cell7.data [7], _25964_);
  and (_00429_, _25849_, _25848_);
  or (_25850_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_25851_, \oc8051_gm_cxrom_1.cell7.data [0], _25845_);
  nand (_25852_, _25851_, _25850_);
  nand (_25853_, _25852_, _25964_);
  or (_25854_, \oc8051_gm_cxrom_1.cell7.data [0], _25964_);
  and (_00461_, _25854_, _25853_);
  or (_25855_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_25856_, \oc8051_gm_cxrom_1.cell7.data [1], _25845_);
  nand (_25857_, _25856_, _25855_);
  nand (_25858_, _25857_, _25964_);
  or (_25859_, \oc8051_gm_cxrom_1.cell7.data [1], _25964_);
  and (_00463_, _25859_, _25858_);
  or (_25860_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_25861_, \oc8051_gm_cxrom_1.cell7.data [2], _25845_);
  nand (_25862_, _25861_, _25860_);
  nand (_25863_, _25862_, _25964_);
  or (_25864_, \oc8051_gm_cxrom_1.cell7.data [2], _25964_);
  and (_00465_, _25864_, _25863_);
  or (_25865_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_25866_, \oc8051_gm_cxrom_1.cell7.data [3], _25845_);
  nand (_25867_, _25866_, _25865_);
  nand (_25868_, _25867_, _25964_);
  or (_25869_, \oc8051_gm_cxrom_1.cell7.data [3], _25964_);
  and (_00467_, _25869_, _25868_);
  or (_25870_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_25871_, \oc8051_gm_cxrom_1.cell7.data [4], _25845_);
  nand (_25872_, _25871_, _25870_);
  nand (_25873_, _25872_, _25964_);
  or (_25874_, \oc8051_gm_cxrom_1.cell7.data [4], _25964_);
  and (_00469_, _25874_, _25873_);
  or (_25875_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_25876_, \oc8051_gm_cxrom_1.cell7.data [5], _25845_);
  nand (_25877_, _25876_, _25875_);
  nand (_25878_, _25877_, _25964_);
  or (_25879_, \oc8051_gm_cxrom_1.cell7.data [5], _25964_);
  and (_00471_, _25879_, _25878_);
  or (_25880_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_25881_, \oc8051_gm_cxrom_1.cell7.data [6], _25845_);
  nand (_25882_, _25881_, _25880_);
  nand (_25883_, _25882_, _25964_);
  or (_25884_, \oc8051_gm_cxrom_1.cell7.data [6], _25964_);
  and (_00473_, _25884_, _25883_);
  or (_25885_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_25886_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_25887_, _25886_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_25888_, _25887_, _25885_);
  nand (_25889_, _25888_, _25964_);
  or (_25890_, \oc8051_gm_cxrom_1.cell8.data [7], _25964_);
  and (_00481_, _25890_, _25889_);
  or (_25891_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_25892_, \oc8051_gm_cxrom_1.cell8.data [0], _25886_);
  nand (_25893_, _25892_, _25891_);
  nand (_25894_, _25893_, _25964_);
  or (_25895_, \oc8051_gm_cxrom_1.cell8.data [0], _25964_);
  and (_00514_, _25895_, _25894_);
  or (_25896_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_25897_, \oc8051_gm_cxrom_1.cell8.data [1], _25886_);
  nand (_25898_, _25897_, _25896_);
  nand (_25899_, _25898_, _25964_);
  or (_25900_, \oc8051_gm_cxrom_1.cell8.data [1], _25964_);
  and (_00516_, _25900_, _25899_);
  or (_25901_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_25902_, \oc8051_gm_cxrom_1.cell8.data [2], _25886_);
  nand (_25903_, _25902_, _25901_);
  nand (_25904_, _25903_, _25964_);
  or (_25905_, \oc8051_gm_cxrom_1.cell8.data [2], _25964_);
  and (_00517_, _25905_, _25904_);
  or (_25906_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_25907_, \oc8051_gm_cxrom_1.cell8.data [3], _25886_);
  nand (_25908_, _25907_, _25906_);
  nand (_25909_, _25908_, _25964_);
  or (_25910_, \oc8051_gm_cxrom_1.cell8.data [3], _25964_);
  and (_00519_, _25910_, _25909_);
  or (_25911_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_25912_, \oc8051_gm_cxrom_1.cell8.data [4], _25886_);
  nand (_25913_, _25912_, _25911_);
  nand (_25914_, _25913_, _25964_);
  or (_25915_, \oc8051_gm_cxrom_1.cell8.data [4], _25964_);
  and (_00521_, _25915_, _25914_);
  or (_25916_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_25917_, \oc8051_gm_cxrom_1.cell8.data [5], _25886_);
  nand (_25918_, _25917_, _25916_);
  nand (_25919_, _25918_, _25964_);
  or (_25920_, \oc8051_gm_cxrom_1.cell8.data [5], _25964_);
  and (_00523_, _25920_, _25919_);
  or (_25921_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_25922_, \oc8051_gm_cxrom_1.cell8.data [6], _25886_);
  nand (_25923_, _25922_, _25921_);
  nand (_25924_, _25923_, _25964_);
  or (_25925_, \oc8051_gm_cxrom_1.cell8.data [6], _25964_);
  and (_00525_, _25925_, _25924_);
  or (_25926_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_25927_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_25928_, _25927_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_25929_, _25928_, _25926_);
  nand (_25930_, _25929_, _25964_);
  or (_25931_, \oc8051_gm_cxrom_1.cell9.data [7], _25964_);
  and (_00533_, _25931_, _25930_);
  or (_25932_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_25933_, \oc8051_gm_cxrom_1.cell9.data [0], _25927_);
  nand (_25934_, _25933_, _25932_);
  nand (_25935_, _25934_, _25964_);
  or (_25936_, \oc8051_gm_cxrom_1.cell9.data [0], _25964_);
  and (_00566_, _25936_, _25935_);
  or (_25937_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_25938_, \oc8051_gm_cxrom_1.cell9.data [1], _25927_);
  nand (_25939_, _25938_, _25937_);
  nand (_25940_, _25939_, _25964_);
  or (_25941_, \oc8051_gm_cxrom_1.cell9.data [1], _25964_);
  and (_00568_, _25941_, _25940_);
  or (_25942_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_25943_, \oc8051_gm_cxrom_1.cell9.data [2], _25927_);
  nand (_25944_, _25943_, _25942_);
  nand (_25945_, _25944_, _25964_);
  or (_25946_, \oc8051_gm_cxrom_1.cell9.data [2], _25964_);
  and (_00570_, _25946_, _25945_);
  or (_25947_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_25948_, \oc8051_gm_cxrom_1.cell9.data [3], _25927_);
  nand (_25949_, _25948_, _25947_);
  nand (_25950_, _25949_, _25964_);
  or (_25951_, \oc8051_gm_cxrom_1.cell9.data [3], _25964_);
  and (_00572_, _25951_, _25950_);
  or (_25952_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_25953_, \oc8051_gm_cxrom_1.cell9.data [4], _25927_);
  nand (_25954_, _25953_, _25952_);
  nand (_25955_, _25954_, _25964_);
  or (_25956_, \oc8051_gm_cxrom_1.cell9.data [4], _25964_);
  and (_00574_, _25956_, _25955_);
  or (_25957_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_25958_, \oc8051_gm_cxrom_1.cell9.data [5], _25927_);
  nand (_25959_, _25958_, _25957_);
  nand (_25960_, _25959_, _25964_);
  or (_25961_, \oc8051_gm_cxrom_1.cell9.data [5], _25964_);
  and (_00575_, _25961_, _25960_);
  or (_25962_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_25963_, \oc8051_gm_cxrom_1.cell9.data [6], _25927_);
  nand (_25965_, _25963_, _25962_);
  nand (_25966_, _25965_, _25964_);
  or (_25968_, \oc8051_gm_cxrom_1.cell9.data [6], _25964_);
  and (_00577_, _25968_, _25966_);
  or (_25970_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_25971_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_25973_, _25971_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_25974_, _25973_, _25970_);
  nand (_25976_, _25974_, _25964_);
  or (_25977_, \oc8051_gm_cxrom_1.cell10.data [7], _25964_);
  and (_00585_, _25977_, _25976_);
  or (_25980_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_25982_, \oc8051_gm_cxrom_1.cell10.data [0], _25971_);
  nand (_25983_, _25982_, _25980_);
  nand (_25984_, _25983_, _25964_);
  or (_25985_, \oc8051_gm_cxrom_1.cell10.data [0], _25964_);
  and (_00617_, _25985_, _25984_);
  or (_25986_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_25987_, \oc8051_gm_cxrom_1.cell10.data [1], _25971_);
  nand (_25988_, _25987_, _25986_);
  nand (_25989_, _25988_, _25964_);
  or (_25990_, \oc8051_gm_cxrom_1.cell10.data [1], _25964_);
  and (_00619_, _25990_, _25989_);
  or (_25991_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_25992_, \oc8051_gm_cxrom_1.cell10.data [2], _25971_);
  nand (_25993_, _25992_, _25991_);
  nand (_25994_, _25993_, _25964_);
  or (_25995_, \oc8051_gm_cxrom_1.cell10.data [2], _25964_);
  and (_00621_, _25995_, _25994_);
  or (_25996_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_25997_, \oc8051_gm_cxrom_1.cell10.data [3], _25971_);
  nand (_25998_, _25997_, _25996_);
  nand (_25999_, _25998_, _25964_);
  or (_26000_, \oc8051_gm_cxrom_1.cell10.data [3], _25964_);
  and (_00623_, _26000_, _25999_);
  or (_26001_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_26002_, \oc8051_gm_cxrom_1.cell10.data [4], _25971_);
  nand (_26003_, _26002_, _26001_);
  nand (_26004_, _26003_, _25964_);
  or (_26005_, \oc8051_gm_cxrom_1.cell10.data [4], _25964_);
  and (_00625_, _26005_, _26004_);
  or (_26006_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_26007_, \oc8051_gm_cxrom_1.cell10.data [5], _25971_);
  nand (_26008_, _26007_, _26006_);
  nand (_26009_, _26008_, _25964_);
  or (_26010_, \oc8051_gm_cxrom_1.cell10.data [5], _25964_);
  and (_00627_, _26010_, _26009_);
  or (_26011_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_26012_, \oc8051_gm_cxrom_1.cell10.data [6], _25971_);
  nand (_26013_, _26012_, _26011_);
  nand (_26014_, _26013_, _25964_);
  or (_26015_, \oc8051_gm_cxrom_1.cell10.data [6], _25964_);
  and (_00629_, _26015_, _26014_);
  or (_26017_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_26019_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_26021_, _26019_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_26023_, _26021_, _26017_);
  nand (_26025_, _26023_, _25964_);
  or (_26026_, \oc8051_gm_cxrom_1.cell11.data [7], _25964_);
  and (_00637_, _26026_, _26025_);
  or (_26029_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_26030_, \oc8051_gm_cxrom_1.cell11.data [0], _26019_);
  nand (_26031_, _26030_, _26029_);
  nand (_26032_, _26031_, _25964_);
  or (_26033_, \oc8051_gm_cxrom_1.cell11.data [0], _25964_);
  and (_00669_, _26033_, _26032_);
  or (_26034_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_26035_, \oc8051_gm_cxrom_1.cell11.data [1], _26019_);
  nand (_26036_, _26035_, _26034_);
  nand (_26037_, _26036_, _25964_);
  or (_26038_, \oc8051_gm_cxrom_1.cell11.data [1], _25964_);
  and (_00671_, _26038_, _26037_);
  or (_26039_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_26040_, \oc8051_gm_cxrom_1.cell11.data [2], _26019_);
  nand (_26041_, _26040_, _26039_);
  nand (_26042_, _26041_, _25964_);
  or (_26043_, \oc8051_gm_cxrom_1.cell11.data [2], _25964_);
  and (_00673_, _26043_, _26042_);
  or (_26044_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_26045_, \oc8051_gm_cxrom_1.cell11.data [3], _26019_);
  nand (_26046_, _26045_, _26044_);
  nand (_26047_, _26046_, _25964_);
  or (_26048_, \oc8051_gm_cxrom_1.cell11.data [3], _25964_);
  and (_00675_, _26048_, _26047_);
  or (_26049_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_26050_, \oc8051_gm_cxrom_1.cell11.data [4], _26019_);
  nand (_26051_, _26050_, _26049_);
  nand (_26052_, _26051_, _25964_);
  or (_26053_, \oc8051_gm_cxrom_1.cell11.data [4], _25964_);
  and (_00677_, _26053_, _26052_);
  or (_26054_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_26055_, \oc8051_gm_cxrom_1.cell11.data [5], _26019_);
  nand (_26056_, _26055_, _26054_);
  nand (_26057_, _26056_, _25964_);
  or (_26058_, \oc8051_gm_cxrom_1.cell11.data [5], _25964_);
  and (_00679_, _26058_, _26057_);
  or (_26059_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_26060_, \oc8051_gm_cxrom_1.cell11.data [6], _26019_);
  nand (_26061_, _26060_, _26059_);
  nand (_26062_, _26061_, _25964_);
  or (_26063_, \oc8051_gm_cxrom_1.cell11.data [6], _25964_);
  and (_00681_, _26063_, _26062_);
  or (_26064_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_26065_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_26066_, _26065_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_26067_, _26066_, _26064_);
  nand (_26068_, _26067_, _25964_);
  or (_26069_, \oc8051_gm_cxrom_1.cell12.data [7], _25964_);
  and (_00688_, _26069_, _26068_);
  or (_26070_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_26071_, \oc8051_gm_cxrom_1.cell12.data [0], _26065_);
  nand (_26072_, _26071_, _26070_);
  nand (_26073_, _26072_, _25964_);
  or (_26074_, \oc8051_gm_cxrom_1.cell12.data [0], _25964_);
  and (_00720_, _26074_, _26073_);
  or (_26075_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_26076_, \oc8051_gm_cxrom_1.cell12.data [1], _26065_);
  nand (_26077_, _26076_, _26075_);
  nand (_26078_, _26077_, _25964_);
  or (_26079_, \oc8051_gm_cxrom_1.cell12.data [1], _25964_);
  and (_00722_, _26079_, _26078_);
  or (_26080_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_26081_, \oc8051_gm_cxrom_1.cell12.data [2], _26065_);
  nand (_26082_, _26081_, _26080_);
  nand (_26083_, _26082_, _25964_);
  or (_26084_, \oc8051_gm_cxrom_1.cell12.data [2], _25964_);
  and (_00724_, _26084_, _26083_);
  or (_26085_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_26086_, \oc8051_gm_cxrom_1.cell12.data [3], _26065_);
  nand (_26087_, _26086_, _26085_);
  nand (_26088_, _26087_, _25964_);
  or (_26089_, \oc8051_gm_cxrom_1.cell12.data [3], _25964_);
  and (_00726_, _26089_, _26088_);
  or (_26090_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_26091_, \oc8051_gm_cxrom_1.cell12.data [4], _26065_);
  nand (_26092_, _26091_, _26090_);
  nand (_26093_, _26092_, _25964_);
  or (_26094_, \oc8051_gm_cxrom_1.cell12.data [4], _25964_);
  and (_00728_, _26094_, _26093_);
  or (_26095_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_26096_, \oc8051_gm_cxrom_1.cell12.data [5], _26065_);
  nand (_26097_, _26096_, _26095_);
  nand (_26098_, _26097_, _25964_);
  or (_26099_, \oc8051_gm_cxrom_1.cell12.data [5], _25964_);
  and (_00730_, _26099_, _26098_);
  or (_26100_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_26101_, \oc8051_gm_cxrom_1.cell12.data [6], _26065_);
  nand (_26102_, _26101_, _26100_);
  nand (_26103_, _26102_, _25964_);
  or (_26104_, \oc8051_gm_cxrom_1.cell12.data [6], _25964_);
  and (_00732_, _26104_, _26103_);
  or (_26105_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_26106_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_26107_, _26106_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_26108_, _26107_, _26105_);
  nand (_26109_, _26108_, _25964_);
  or (_26110_, \oc8051_gm_cxrom_1.cell13.data [7], _25964_);
  and (_00740_, _26110_, _26109_);
  or (_26111_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_26112_, \oc8051_gm_cxrom_1.cell13.data [0], _26106_);
  nand (_26113_, _26112_, _26111_);
  nand (_26114_, _26113_, _25964_);
  or (_26115_, \oc8051_gm_cxrom_1.cell13.data [0], _25964_);
  and (_00772_, _26115_, _26114_);
  or (_26116_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_26117_, \oc8051_gm_cxrom_1.cell13.data [1], _26106_);
  nand (_26118_, _26117_, _26116_);
  nand (_26119_, _26118_, _25964_);
  or (_26120_, \oc8051_gm_cxrom_1.cell13.data [1], _25964_);
  and (_00774_, _26120_, _26119_);
  or (_26121_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_26122_, \oc8051_gm_cxrom_1.cell13.data [2], _26106_);
  nand (_26123_, _26122_, _26121_);
  nand (_26124_, _26123_, _25964_);
  or (_26125_, \oc8051_gm_cxrom_1.cell13.data [2], _25964_);
  and (_00776_, _26125_, _26124_);
  or (_26126_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_26127_, \oc8051_gm_cxrom_1.cell13.data [3], _26106_);
  nand (_26128_, _26127_, _26126_);
  nand (_26129_, _26128_, _25964_);
  or (_26130_, \oc8051_gm_cxrom_1.cell13.data [3], _25964_);
  and (_00778_, _26130_, _26129_);
  or (_26131_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_26132_, \oc8051_gm_cxrom_1.cell13.data [4], _26106_);
  nand (_26133_, _26132_, _26131_);
  nand (_26134_, _26133_, _25964_);
  or (_26135_, \oc8051_gm_cxrom_1.cell13.data [4], _25964_);
  and (_00780_, _26135_, _26134_);
  or (_26136_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_26137_, \oc8051_gm_cxrom_1.cell13.data [5], _26106_);
  nand (_26138_, _26137_, _26136_);
  nand (_26139_, _26138_, _25964_);
  or (_26140_, \oc8051_gm_cxrom_1.cell13.data [5], _25964_);
  and (_00782_, _26140_, _26139_);
  or (_26141_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_26142_, \oc8051_gm_cxrom_1.cell13.data [6], _26106_);
  nand (_26143_, _26142_, _26141_);
  nand (_26144_, _26143_, _25964_);
  or (_26145_, \oc8051_gm_cxrom_1.cell13.data [6], _25964_);
  and (_00784_, _26145_, _26144_);
  or (_26146_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_26147_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_26148_, _26147_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_26149_, _26148_, _26146_);
  nand (_26150_, _26149_, _25964_);
  or (_26151_, \oc8051_gm_cxrom_1.cell14.data [7], _25964_);
  and (_00792_, _26151_, _26150_);
  or (_26152_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_26153_, \oc8051_gm_cxrom_1.cell14.data [0], _26147_);
  nand (_26154_, _26153_, _26152_);
  nand (_26155_, _26154_, _25964_);
  or (_26156_, \oc8051_gm_cxrom_1.cell14.data [0], _25964_);
  and (_00824_, _26156_, _26155_);
  or (_26157_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_26158_, \oc8051_gm_cxrom_1.cell14.data [1], _26147_);
  nand (_26159_, _26158_, _26157_);
  nand (_26160_, _26159_, _25964_);
  or (_26161_, \oc8051_gm_cxrom_1.cell14.data [1], _25964_);
  and (_00826_, _26161_, _26160_);
  or (_26162_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_26163_, \oc8051_gm_cxrom_1.cell14.data [2], _26147_);
  nand (_26164_, _26163_, _26162_);
  nand (_26165_, _26164_, _25964_);
  or (_26166_, \oc8051_gm_cxrom_1.cell14.data [2], _25964_);
  and (_00827_, _26166_, _26165_);
  or (_26167_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_26168_, \oc8051_gm_cxrom_1.cell14.data [3], _26147_);
  nand (_26169_, _26168_, _26167_);
  nand (_26170_, _26169_, _25964_);
  or (_26171_, \oc8051_gm_cxrom_1.cell14.data [3], _25964_);
  and (_00829_, _26171_, _26170_);
  or (_26172_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_26173_, \oc8051_gm_cxrom_1.cell14.data [4], _26147_);
  nand (_26174_, _26173_, _26172_);
  nand (_26175_, _26174_, _25964_);
  or (_26176_, \oc8051_gm_cxrom_1.cell14.data [4], _25964_);
  and (_00831_, _26176_, _26175_);
  or (_26177_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_26178_, \oc8051_gm_cxrom_1.cell14.data [5], _26147_);
  nand (_26179_, _26178_, _26177_);
  nand (_26180_, _26179_, _25964_);
  or (_26181_, \oc8051_gm_cxrom_1.cell14.data [5], _25964_);
  and (_00833_, _26181_, _26180_);
  or (_26182_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_26183_, \oc8051_gm_cxrom_1.cell14.data [6], _26147_);
  nand (_26184_, _26183_, _26182_);
  nand (_26185_, _26184_, _25964_);
  or (_26186_, \oc8051_gm_cxrom_1.cell14.data [6], _25964_);
  and (_00835_, _26186_, _26185_);
  or (_26187_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_26188_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_26189_, _26188_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_26190_, _26189_, _26187_);
  nand (_26191_, _26190_, _25964_);
  or (_26192_, \oc8051_gm_cxrom_1.cell15.data [7], _25964_);
  and (_00843_, _26192_, _26191_);
  or (_26193_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_26194_, \oc8051_gm_cxrom_1.cell15.data [0], _26188_);
  nand (_26195_, _26194_, _26193_);
  nand (_26196_, _26195_, _25964_);
  or (_26197_, \oc8051_gm_cxrom_1.cell15.data [0], _25964_);
  and (_00875_, _26197_, _26196_);
  or (_26198_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_26199_, \oc8051_gm_cxrom_1.cell15.data [1], _26188_);
  nand (_26200_, _26199_, _26198_);
  nand (_26201_, _26200_, _25964_);
  or (_26202_, \oc8051_gm_cxrom_1.cell15.data [1], _25964_);
  and (_00877_, _26202_, _26201_);
  or (_26203_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_26204_, \oc8051_gm_cxrom_1.cell15.data [2], _26188_);
  nand (_26205_, _26204_, _26203_);
  nand (_26206_, _26205_, _25964_);
  or (_26207_, \oc8051_gm_cxrom_1.cell15.data [2], _25964_);
  and (_00879_, _26207_, _26206_);
  or (_26208_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_26209_, \oc8051_gm_cxrom_1.cell15.data [3], _26188_);
  nand (_26210_, _26209_, _26208_);
  nand (_26211_, _26210_, _25964_);
  or (_26212_, \oc8051_gm_cxrom_1.cell15.data [3], _25964_);
  and (_00881_, _26212_, _26211_);
  or (_26213_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_26214_, \oc8051_gm_cxrom_1.cell15.data [4], _26188_);
  nand (_26215_, _26214_, _26213_);
  nand (_26216_, _26215_, _25964_);
  or (_26217_, \oc8051_gm_cxrom_1.cell15.data [4], _25964_);
  and (_00883_, _26217_, _26216_);
  or (_26218_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_26219_, \oc8051_gm_cxrom_1.cell15.data [5], _26188_);
  nand (_26220_, _26219_, _26218_);
  nand (_26221_, _26220_, _25964_);
  or (_26222_, \oc8051_gm_cxrom_1.cell15.data [5], _25964_);
  and (_00885_, _26222_, _26221_);
  or (_26223_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_26224_, \oc8051_gm_cxrom_1.cell15.data [6], _26188_);
  nand (_26225_, _26224_, _26223_);
  nand (_26226_, _26225_, _25964_);
  or (_26227_, \oc8051_gm_cxrom_1.cell15.data [6], _25964_);
  and (_00887_, _26227_, _26226_);
  nor (_00918_, _19135_, rst);
  nor (_00922_, _24335_, rst);
  and (_26228_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_26229_, _18850_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_26230_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_26231_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_26232_, _26231_, _26230_);
  and (_26233_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_26234_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_26235_, _26234_, _26233_);
  and (_26236_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_26237_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_26238_, _26237_, _26236_);
  and (_26239_, _26238_, _26235_);
  and (_26240_, _26239_, _26232_);
  nor (_26241_, _26240_, _18850_);
  nor (_26242_, _26241_, _26229_);
  nor (_26243_, _26242_, _24319_);
  nor (_26244_, _26243_, _26228_);
  nor (_00926_, _26244_, rst);
  nor (_01047_, _19962_, rst);
  and (_01050_, _20214_, _25964_);
  nor (_01053_, _20445_, rst);
  nor (_01056_, _20686_, rst);
  and (_01058_, _19442_, _25964_);
  nor (_01061_, _19699_, rst);
  nor (_01064_, _18905_, rst);
  nor (_01067_, _24527_, rst);
  nor (_01070_, _24675_, rst);
  nor (_01073_, _24446_, rst);
  nor (_01076_, _24491_, rst);
  nor (_01079_, _24633_, rst);
  nor (_01082_, _24420_, rst);
  nor (_01085_, _24586_, rst);
  and (_26245_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_26246_, _18850_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_26247_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_26248_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_26249_, _26248_, _26247_);
  and (_26250_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_26251_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_26252_, _26251_, _26250_);
  and (_26253_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_26254_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_26255_, _26254_, _26253_);
  and (_26256_, _26255_, _26252_);
  and (_26257_, _26256_, _26249_);
  nor (_26258_, _26257_, _18850_);
  nor (_26259_, _26258_, _26246_);
  nor (_26260_, _26259_, _24319_);
  nor (_26261_, _26260_, _26245_);
  nor (_01088_, _26261_, rst);
  and (_26262_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_26263_, _18850_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_26264_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_26265_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_26266_, _26265_, _26264_);
  and (_26267_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_26268_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_26269_, _26268_, _26267_);
  and (_26270_, _26269_, _26266_);
  and (_26271_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_26272_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_26273_, _26272_, _26271_);
  and (_26274_, _26273_, _26270_);
  nor (_26275_, _26274_, _18850_);
  nor (_26276_, _26275_, _26263_);
  nor (_26277_, _26276_, _24319_);
  nor (_26278_, _26277_, _26262_);
  nor (_01091_, _26278_, rst);
  and (_26279_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_26280_, _18850_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_26281_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_26282_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_26283_, _26282_, _26281_);
  and (_26284_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_26285_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_26286_, _26285_, _26284_);
  and (_26287_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_26288_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_26289_, _26288_, _26287_);
  and (_26290_, _26289_, _26286_);
  and (_26291_, _26290_, _26283_);
  nor (_26292_, _26291_, _18850_);
  nor (_26293_, _26292_, _26280_);
  nor (_26294_, _26293_, _24319_);
  nor (_26295_, _26294_, _26279_);
  nor (_01094_, _26295_, rst);
  and (_26296_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_26297_, _18850_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_26298_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_26299_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_26300_, _26299_, _26298_);
  and (_26301_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_26302_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_26303_, _26302_, _26301_);
  and (_26304_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_26305_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_26306_, _26305_, _26304_);
  and (_26307_, _26306_, _26303_);
  and (_26308_, _26307_, _26300_);
  nor (_26309_, _26308_, _18850_);
  nor (_26310_, _26309_, _26297_);
  nor (_26311_, _26310_, _24319_);
  nor (_26312_, _26311_, _26296_);
  nor (_01097_, _26312_, rst);
  and (_26313_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_26314_, _18850_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_26315_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_26316_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_26317_, _26316_, _26315_);
  and (_26318_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_26319_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_26320_, _26319_, _26318_);
  and (_26321_, _26320_, _26317_);
  and (_26322_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_26323_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_26324_, _26323_, _26322_);
  and (_26325_, _26324_, _26321_);
  nor (_26326_, _26325_, _18850_);
  nor (_26327_, _26326_, _26314_);
  nor (_26328_, _26327_, _24319_);
  nor (_26329_, _26328_, _26313_);
  nor (_01100_, _26329_, rst);
  and (_26330_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_26331_, _18850_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_26332_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_26333_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_26334_, _26333_, _26332_);
  and (_26335_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_26336_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_26337_, _26336_, _26335_);
  and (_26338_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_26339_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_26340_, _26339_, _26338_);
  and (_26341_, _26340_, _26337_);
  and (_26342_, _26341_, _26334_);
  nor (_26343_, _26342_, _18850_);
  nor (_26344_, _26343_, _26331_);
  nor (_26345_, _26344_, _24319_);
  nor (_26346_, _26345_, _26330_);
  nor (_01103_, _26346_, rst);
  and (_26347_, _24319_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_26348_, _18850_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_26349_, _18696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_26350_, _18653_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_26351_, _26350_, _26349_);
  and (_26352_, _18598_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_26353_, _18740_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_26354_, _26353_, _26352_);
  and (_26355_, _26354_, _26351_);
  and (_26356_, _18784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_26357_, _18806_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_26358_, _26357_, _26356_);
  and (_26359_, _26358_, _26355_);
  nor (_26360_, _26359_, _18850_);
  nor (_26361_, _26360_, _26348_);
  nor (_26362_, _26361_, _24319_);
  nor (_26363_, _26362_, _26347_);
  nor (_01105_, _26363_, rst);
  and (_26364_, _24511_, _24642_);
  nor (_26365_, _24591_, _24377_);
  and (_26366_, _26365_, _24431_);
  and (_26367_, _26366_, _26364_);
  and (_26368_, _26367_, _23313_);
  not (_26369_, _26367_);
  and (_26370_, _24643_, _24430_);
  and (_26371_, _26365_, _26370_);
  and (_26372_, _26371_, _24511_);
  and (_26373_, _24591_, _24430_);
  nor (_26374_, _24642_, _24377_);
  and (_26375_, _26374_, _26373_);
  and (_26376_, _26375_, _24512_);
  nor (_26377_, _26376_, _26372_);
  and (_26378_, _26377_, _26369_);
  and (_26379_, _24591_, _24431_);
  nor (_26380_, _24643_, _24377_);
  and (_26381_, _26380_, _26379_);
  and (_26382_, _26381_, _24511_);
  and (_26383_, _26373_, _26380_);
  and (_26384_, _26383_, _24511_);
  nor (_26385_, _26384_, _26382_);
  and (_26386_, _26374_, _26379_);
  and (_26387_, _26386_, _24511_);
  and (_26388_, _26375_, _24511_);
  nor (_26389_, _26388_, _26387_);
  and (_26390_, _26389_, _26385_);
  and (_26391_, _26386_, _24512_);
  not (_26392_, _26391_);
  and (_26393_, _26380_, _24512_);
  and (_26394_, _26393_, _24591_);
  nor (_26395_, _24512_, _24642_);
  and (_26396_, _26366_, _26395_);
  nor (_26397_, _26396_, _26394_);
  and (_26398_, _26397_, _26392_);
  and (_26399_, _26398_, _26390_);
  and (_26400_, _26399_, _26378_);
  and (_26401_, _24642_, _24032_);
  nor (_26402_, _24642_, _24032_);
  or (_26403_, _26402_, _26401_);
  not (_26404_, _26403_);
  nor (_26405_, _24430_, _23315_);
  and (_26406_, _24430_, _23315_);
  nor (_26407_, _26406_, _26405_);
  and (_26408_, _24591_, _22626_);
  nor (_26409_, _24591_, _22626_);
  nor (_26410_, _26409_, _26408_);
  and (_26411_, _26410_, _26407_);
  nor (_26412_, _24377_, _16216_);
  and (_26413_, _24377_, _16216_);
  nor (_26414_, _26413_, _26412_);
  nor (_26415_, _24511_, _16400_);
  and (_26416_, _24511_, _16400_);
  nor (_26417_, _26416_, _26415_);
  and (_26418_, _26417_, _26414_);
  and (_26419_, _26418_, _26411_);
  and (_26420_, _26419_, _26404_);
  nor (_26421_, _24680_, _17561_);
  and (_26422_, _24680_, _17561_);
  nor (_26423_, _26422_, _26421_);
  nor (_26424_, _24547_, _17366_);
  and (_26425_, _24547_, _17366_);
  nor (_26426_, _26425_, _26424_);
  nor (_26427_, _24467_, _16727_);
  and (_26428_, _24467_, _16727_);
  nor (_26429_, _26428_, _26427_);
  and (_26430_, _26429_, _26426_);
  and (_26431_, _26430_, _26423_);
  and (_26432_, _26431_, _26420_);
  nand (_26433_, _26432_, _15585_);
  or (_26434_, _26433_, _26400_);
  or (_26435_, _26434_, ABINPUT[0]);
  not (_26436_, _24467_);
  nor (_26437_, _24547_, _24680_);
  and (_26438_, _26437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  not (_26439_, _24547_);
  and (_26440_, _26439_, _24680_);
  and (_26441_, _26440_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_26442_, _26441_, _26438_);
  nor (_26443_, _26439_, _24680_);
  and (_26444_, _26443_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_26445_, _24547_, _24680_);
  and (_26446_, _26445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_26447_, _26446_, _26444_);
  or (_26448_, _26447_, _26442_);
  and (_26449_, _26448_, _26436_);
  and (_26450_, _26443_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_26451_, _26445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_26452_, _26451_, _26450_);
  and (_26453_, _26440_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_26454_, _26437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_26455_, _26454_, _26453_);
  or (_26456_, _26455_, _26452_);
  and (_26457_, _26456_, _24467_);
  or (_26458_, _26457_, _26449_);
  and (_26459_, _26458_, _26391_);
  and (_26460_, _26443_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_26461_, _26437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_26462_, _26461_, _26460_);
  and (_26463_, _26445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_26464_, _26440_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_26465_, _26464_, _26463_);
  or (_26466_, _26465_, _26462_);
  and (_26467_, _26466_, _26436_);
  and (_26468_, _26443_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_26469_, _26437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_26470_, _26469_, _26468_);
  and (_26471_, _26445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_26472_, _26440_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_26473_, _26472_, _26471_);
  or (_26474_, _26473_, _26470_);
  and (_26475_, _26474_, _24467_);
  or (_26476_, _26475_, _26467_);
  and (_26477_, _26394_, _24431_);
  and (_26478_, _26477_, _26476_);
  or (_26479_, _26478_, _26459_);
  and (_26480_, _20708_, _19464_);
  and (_26481_, _26480_, _21180_);
  nor (_26482_, _26481_, _22232_);
  not (_26483_, _21662_);
  and (_26484_, _21980_, _21256_);
  and (_26485_, _21585_, _20927_);
  nor (_26486_, _26485_, _26484_);
  and (_26487_, _26486_, _26483_);
  and (_26488_, _21541_, _20927_);
  nor (_26489_, _26488_, _21333_);
  and (_26490_, _26489_, _26487_);
  and (_26491_, _26490_, _26482_);
  and (_26492_, _21015_, _21234_);
  and (_26493_, _26492_, _21190_);
  not (_26494_, _26493_);
  and (_26495_, _26494_, _21212_);
  nor (_26496_, _22309_, _21695_);
  nor (_26497_, _21432_, _21322_);
  nor (_26498_, _26497_, _21004_);
  not (_26499_, _26498_);
  and (_26500_, _26499_, _26496_);
  and (_26501_, _26500_, _26495_);
  and (_26502_, _26501_, _26491_);
  and (_26503_, _26502_, _21947_);
  nor (_26504_, _26503_, _18477_);
  and (_26505_, _18532_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_26506_, _26505_);
  and (_26507_, _26506_, p0in_reg[6]);
  and (_26508_, _26505_, p0_in[6]);
  or (_26509_, _26508_, _26507_);
  or (_26510_, _26509_, _26504_);
  not (_26511_, _26504_);
  or (_26512_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_26513_, _26512_, _26510_);
  and (_26514_, _26513_, _26436_);
  and (_26515_, _26506_, p0in_reg[2]);
  and (_26516_, _26505_, p0_in[2]);
  or (_26517_, _26516_, _26515_);
  or (_26518_, _26517_, _26504_);
  nand (_26519_, _26504_, _23506_);
  and (_26520_, _26519_, _26518_);
  and (_26521_, _26520_, _24467_);
  or (_26522_, _26521_, _26514_);
  and (_26523_, _26522_, _26443_);
  and (_26524_, _26506_, p0in_reg[1]);
  and (_26525_, _26505_, p0_in[1]);
  or (_26526_, _26525_, _26524_);
  or (_26527_, _26526_, _26504_);
  or (_26528_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_26529_, _26528_, _26527_);
  or (_26530_, _26529_, _26436_);
  and (_26531_, _26506_, p0in_reg[5]);
  and (_26532_, _26505_, p0_in[5]);
  or (_26533_, _26532_, _26531_);
  or (_26534_, _26533_, _26504_);
  or (_26535_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_26536_, _26535_, _26534_);
  or (_26537_, _26536_, _24467_);
  and (_26538_, _26537_, _26440_);
  and (_26539_, _26538_, _26530_);
  and (_26540_, _26506_, p0in_reg[7]);
  and (_26541_, _26505_, p0_in[7]);
  or (_26542_, _26541_, _26540_);
  or (_26543_, _26542_, _26504_);
  or (_26544_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_26545_, _26544_, _26543_);
  and (_26546_, _26545_, _26436_);
  and (_26547_, _26506_, p0in_reg[3]);
  and (_26548_, _26505_, p0_in[3]);
  or (_26549_, _26548_, _26547_);
  or (_26550_, _26549_, _26504_);
  or (_26551_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_26552_, _26551_, _26550_);
  and (_26553_, _26552_, _24467_);
  or (_26554_, _26553_, _26546_);
  and (_26555_, _26554_, _26437_);
  and (_26556_, _26506_, p0in_reg[0]);
  and (_26557_, _26505_, p0_in[0]);
  or (_26558_, _26557_, _26556_);
  or (_26559_, _26558_, _26504_);
  nand (_26560_, _26504_, _23484_);
  and (_26561_, _26560_, _26559_);
  or (_26562_, _26561_, _26436_);
  and (_26563_, _26506_, p0in_reg[4]);
  and (_26564_, _26505_, p0_in[4]);
  or (_26565_, _26564_, _26563_);
  or (_26566_, _26565_, _26504_);
  or (_26567_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_26568_, _26567_, _26566_);
  or (_26569_, _26568_, _24467_);
  and (_26570_, _26569_, _26445_);
  and (_26571_, _26570_, _26562_);
  or (_26572_, _26571_, _26555_);
  or (_26573_, _26572_, _26539_);
  or (_26574_, _26573_, _26523_);
  and (_26575_, _26574_, _26384_);
  and (_26576_, _26506_, p2in_reg[2]);
  and (_26577_, _26505_, p2_in[2]);
  or (_26578_, _26577_, _26576_);
  or (_26579_, _26578_, _26504_);
  or (_26580_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_26581_, _26580_, _26579_);
  or (_26582_, _26581_, _26436_);
  and (_26583_, _26506_, p2in_reg[6]);
  and (_26584_, _26505_, p2_in[6]);
  or (_26585_, _26584_, _26583_);
  or (_26586_, _26585_, _26504_);
  or (_26587_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_26588_, _26587_, _26586_);
  or (_26589_, _26588_, _24467_);
  and (_26590_, _26589_, _26443_);
  and (_26591_, _26590_, _26582_);
  and (_26592_, _26506_, p2in_reg[5]);
  and (_26593_, _26505_, p2_in[5]);
  or (_26594_, _26593_, _26592_);
  or (_26595_, _26594_, _26504_);
  or (_26596_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_26597_, _26596_, _26595_);
  and (_26598_, _26597_, _26436_);
  and (_26599_, _26506_, p2in_reg[1]);
  and (_26600_, _26505_, p2_in[1]);
  or (_26601_, _26600_, _26599_);
  or (_26602_, _26601_, _26504_);
  or (_26603_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_26604_, _26603_, _26602_);
  and (_26605_, _26604_, _24467_);
  or (_26606_, _26605_, _26598_);
  and (_26607_, _26606_, _26440_);
  and (_26608_, _26506_, p2in_reg[4]);
  and (_26609_, _26505_, p2_in[4]);
  or (_26610_, _26609_, _26608_);
  or (_26611_, _26610_, _26504_);
  or (_26612_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_26613_, _26612_, _26611_);
  and (_26614_, _26613_, _26436_);
  and (_26615_, _26506_, p2in_reg[0]);
  and (_26616_, _26505_, p2_in[0]);
  or (_26617_, _26616_, _26615_);
  or (_26618_, _26617_, _26504_);
  or (_26619_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_26620_, _26619_, _26618_);
  and (_26621_, _26620_, _24467_);
  or (_26622_, _26621_, _26614_);
  and (_26623_, _26622_, _26445_);
  and (_26624_, _26506_, p2in_reg[3]);
  and (_26625_, _26505_, p2_in[3]);
  or (_26626_, _26625_, _26624_);
  or (_26627_, _26626_, _26504_);
  or (_26628_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_26629_, _26628_, _26627_);
  or (_26630_, _26629_, _26436_);
  and (_26631_, _26506_, p2in_reg[7]);
  and (_26632_, _26505_, p2_in[7]);
  or (_26633_, _26632_, _26631_);
  or (_26634_, _26633_, _26504_);
  or (_26635_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_26636_, _26635_, _26634_);
  or (_26637_, _26636_, _24467_);
  and (_26638_, _26637_, _26437_);
  and (_26639_, _26638_, _26630_);
  or (_26640_, _26639_, _26623_);
  or (_26641_, _26640_, _26607_);
  or (_26642_, _26641_, _26591_);
  and (_26643_, _26642_, _26382_);
  or (_26644_, _26643_, _26575_);
  or (_26645_, _26644_, _26479_);
  and (_26646_, _26436_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_26647_, _24467_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_26648_, _26647_, _26646_);
  and (_26649_, _26648_, _26443_);
  or (_26650_, _26436_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_26651_, _24467_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_26652_, _26651_, _26440_);
  and (_26653_, _26652_, _26650_);
  and (_26654_, _26436_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_26655_, _24467_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_26656_, _26655_, _26654_);
  and (_26657_, _26656_, _26437_);
  or (_26658_, _26436_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_26659_, _24467_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_26660_, _26659_, _26445_);
  and (_26661_, _26660_, _26658_);
  or (_26662_, _26661_, _26657_);
  or (_26663_, _26662_, _26653_);
  or (_26664_, _26663_, _26649_);
  and (_26665_, _26664_, _26367_);
  nor (_26666_, _23379_, _23369_);
  and (_26667_, _23379_, _23369_);
  nor (_26668_, _26667_, _26666_);
  and (_26669_, _23359_, _23348_);
  nor (_26670_, _23359_, _23348_);
  or (_26671_, _26670_, _26669_);
  nor (_26672_, _26671_, _26668_);
  and (_26673_, _26671_, _26668_);
  nor (_26674_, _26673_, _26672_);
  and (_26675_, _23394_, _23334_);
  nor (_26676_, _23394_, _23334_);
  or (_26677_, _26676_, _26675_);
  not (_26678_, _26677_);
  not (_26679_, _23415_);
  and (_26680_, _26679_, _23404_);
  nor (_26681_, _26679_, _23404_);
  nor (_26682_, _26681_, _26680_);
  and (_26683_, _26682_, _26678_);
  nor (_26684_, _26682_, _26678_);
  nor (_26685_, _26684_, _26683_);
  or (_26686_, _26685_, _26674_);
  nand (_26687_, _26685_, _26674_);
  and (_26688_, _26687_, _26686_);
  and (_26689_, _26688_, _26445_);
  and (_26690_, _26443_, _23273_);
  or (_26691_, _26690_, _26689_);
  and (_26692_, _26691_, _24467_);
  and (_26693_, _26436_, _23295_);
  and (_26694_, _24467_, _23260_);
  or (_26695_, _26694_, _26693_);
  and (_26696_, _26695_, _26440_);
  and (_26697_, _26436_, _23252_);
  and (_26698_, _24467_, _23280_);
  or (_26699_, _26698_, _26697_);
  and (_26700_, _26699_, _26437_);
  or (_26701_, _26700_, _26696_);
  and (_26702_, _26445_, _23287_);
  and (_26703_, _26443_, _23308_);
  or (_26704_, _26703_, _26702_);
  and (_26705_, _26704_, _26436_);
  or (_26706_, _26705_, _26701_);
  or (_26707_, _26706_, _26692_);
  and (_26708_, _26707_, _26372_);
  or (_26709_, _26708_, _26665_);
  nand (_26710_, _24467_, _17226_);
  or (_26711_, _24467_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_26712_, _26711_, _26445_);
  and (_26713_, _26712_, _26710_);
  and (_26714_, _26436_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_26715_, _24467_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_26716_, _26715_, _26714_);
  and (_26717_, _26716_, _26443_);
  and (_26718_, _26436_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_26719_, _24467_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_26720_, _26719_, _26718_);
  and (_26721_, _26720_, _26440_);
  or (_26722_, _26721_, _26717_);
  or (_26723_, _26436_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_26724_, _24467_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_26725_, _26724_, _26437_);
  and (_26726_, _26725_, _26723_);
  or (_26727_, _26726_, _26722_);
  or (_26728_, _26727_, _26713_);
  and (_26729_, _26728_, _26396_);
  and (_26730_, _26506_, p1in_reg[4]);
  and (_26731_, _26505_, p1_in[4]);
  or (_26732_, _26731_, _26730_);
  or (_26733_, _26732_, _26504_);
  or (_26734_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_26735_, _26734_, _26733_);
  and (_26736_, _26735_, _26445_);
  and (_26737_, _26506_, p1in_reg[6]);
  and (_26738_, _26505_, p1_in[6]);
  or (_26739_, _26738_, _26737_);
  or (_26740_, _26739_, _26504_);
  or (_26741_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_26742_, _26741_, _26740_);
  and (_26743_, _26742_, _26443_);
  or (_26744_, _26743_, _26736_);
  and (_26745_, _26506_, p1in_reg[5]);
  and (_26746_, _26505_, p1_in[5]);
  or (_26747_, _26746_, _26745_);
  or (_26748_, _26747_, _26504_);
  or (_26749_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_26750_, _26749_, _26748_);
  and (_26751_, _26750_, _26440_);
  and (_26752_, _26506_, p1in_reg[7]);
  and (_26753_, _26505_, p1_in[7]);
  or (_26754_, _26753_, _26752_);
  or (_26755_, _26754_, _26504_);
  or (_26756_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_26757_, _26756_, _26755_);
  and (_26758_, _26757_, _26437_);
  or (_26759_, _26758_, _26751_);
  or (_26760_, _26759_, _26744_);
  and (_26761_, _26760_, _26436_);
  and (_26762_, _26506_, p1in_reg[1]);
  and (_26763_, _26505_, p1_in[1]);
  or (_26764_, _26763_, _26762_);
  or (_26765_, _26764_, _26504_);
  or (_26766_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_26767_, _26766_, _26765_);
  and (_26768_, _26767_, _26440_);
  and (_26769_, _26506_, p1in_reg[3]);
  and (_26770_, _26505_, p1_in[3]);
  or (_26771_, _26770_, _26769_);
  or (_26772_, _26771_, _26504_);
  or (_26773_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_26774_, _26773_, _26772_);
  and (_26775_, _26774_, _26437_);
  or (_26776_, _26775_, _26768_);
  and (_26777_, _26506_, p1in_reg[2]);
  and (_26778_, _26505_, p1_in[2]);
  or (_26779_, _26778_, _26777_);
  or (_26780_, _26779_, _26504_);
  or (_26781_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_26782_, _26781_, _26780_);
  and (_26783_, _26782_, _26443_);
  and (_26784_, _26506_, p1in_reg[0]);
  and (_26785_, _26505_, p1_in[0]);
  or (_26786_, _26785_, _26784_);
  or (_26787_, _26786_, _26504_);
  or (_26788_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_26789_, _26788_, _26787_);
  and (_26790_, _26789_, _26445_);
  or (_26791_, _26790_, _26783_);
  or (_26792_, _26791_, _26776_);
  and (_26793_, _26792_, _24467_);
  or (_26794_, _26793_, _26761_);
  and (_26795_, _26794_, _26388_);
  or (_26796_, _26795_, _26729_);
  or (_26797_, _26796_, _26709_);
  and (_26798_, _26393_, _26373_);
  and (_26799_, _26440_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_26800_, _26437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_26801_, _26800_, _26799_);
  and (_26802_, _26445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_26803_, _26443_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_26804_, _26803_, _26802_);
  or (_26805_, _26804_, _26801_);
  and (_26806_, _26805_, _24467_);
  and (_26807_, _26440_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_26808_, _26437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_26809_, _26808_, _26807_);
  and (_26810_, _26445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_26811_, _26443_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_26812_, _26811_, _26810_);
  or (_26813_, _26812_, _26809_);
  and (_26814_, _26813_, _26436_);
  or (_26815_, _26814_, _26806_);
  and (_26816_, _26815_, _26798_);
  and (_26817_, _26506_, p3in_reg[7]);
  and (_26818_, _26505_, p3_in[7]);
  or (_26819_, _26818_, _26817_);
  or (_26820_, _26819_, _26504_);
  or (_26821_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_26822_, _26821_, _26820_);
  and (_26823_, _26822_, _26437_);
  and (_26824_, _26506_, p3in_reg[5]);
  and (_26825_, _26505_, p3_in[5]);
  or (_26826_, _26825_, _26824_);
  or (_26827_, _26826_, _26504_);
  or (_26828_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_26829_, _26828_, _26827_);
  and (_26830_, _26829_, _26440_);
  or (_26831_, _26830_, _26823_);
  and (_26832_, _26831_, _26436_);
  and (_26833_, _26506_, p3in_reg[4]);
  and (_26834_, _26505_, p3_in[4]);
  or (_26835_, _26834_, _26833_);
  or (_26836_, _26835_, _26504_);
  or (_26837_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_26838_, _26837_, _26836_);
  and (_26839_, _26838_, _26436_);
  and (_26840_, _26506_, p3in_reg[0]);
  and (_26841_, _26505_, p3_in[0]);
  or (_26842_, _26841_, _26840_);
  or (_26843_, _26842_, _26504_);
  or (_26844_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_26845_, _26844_, _26843_);
  and (_26846_, _26845_, _24467_);
  or (_26847_, _26846_, _26839_);
  and (_26848_, _26847_, _26445_);
  and (_26849_, _26506_, p3in_reg[6]);
  and (_26850_, _26505_, p3_in[6]);
  or (_26851_, _26850_, _26849_);
  or (_26852_, _26851_, _26504_);
  or (_26853_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_26854_, _26853_, _26852_);
  and (_26855_, _26854_, _26436_);
  and (_26856_, _26506_, p3in_reg[2]);
  and (_26857_, _26505_, p3_in[2]);
  or (_26858_, _26857_, _26856_);
  or (_26859_, _26858_, _26504_);
  or (_26860_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_26861_, _26860_, _26859_);
  and (_26862_, _26861_, _24467_);
  or (_26863_, _26862_, _26855_);
  and (_26864_, _26863_, _26443_);
  or (_26865_, _26864_, _26848_);
  and (_26866_, _26506_, p3in_reg[3]);
  and (_26867_, _26505_, p3_in[3]);
  or (_26868_, _26867_, _26866_);
  or (_26869_, _26868_, _26504_);
  or (_26870_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_26871_, _26870_, _26869_);
  and (_26872_, _26871_, _26437_);
  and (_26873_, _26506_, p3in_reg[1]);
  and (_26874_, _26505_, p3_in[1]);
  or (_26875_, _26874_, _26873_);
  or (_26876_, _26875_, _26504_);
  or (_26877_, _26511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_26878_, _26877_, _26876_);
  and (_26879_, _26878_, _26440_);
  or (_26880_, _26879_, _26872_);
  and (_26881_, _26880_, _24467_);
  or (_26882_, _26881_, _26865_);
  or (_26883_, _26882_, _26832_);
  and (_26884_, _26883_, _26387_);
  nor (_26885_, _26884_, _26816_);
  nand (_26886_, _26885_, _26434_);
  or (_26887_, _26886_, _26797_);
  or (_26888_, _26887_, _26645_);
  nand (_26889_, _26888_, _26435_);
  nor (_26890_, _26889_, _26368_);
  not (_26891_, _26400_);
  nor (_26892_, _26504_, _26390_);
  not (_26893_, _26892_);
  and (_26894_, _26420_, _23247_);
  and (_26895_, _26894_, _26893_);
  and (_26896_, _26895_, _26891_);
  nand (_26897_, _26436_, _23404_);
  nand (_26898_, _24467_, _23359_);
  and (_26899_, _26898_, _26440_);
  and (_26900_, _26899_, _26897_);
  nor (_26901_, _24467_, _23415_);
  nor (_26902_, _26436_, _23369_);
  or (_26903_, _26902_, _26901_);
  and (_26904_, _26903_, _26443_);
  nor (_26905_, _24467_, _23394_);
  nor (_26906_, _26436_, _23348_);
  or (_26907_, _26906_, _26905_);
  and (_26908_, _26907_, _26445_);
  nand (_26909_, _26436_, _23334_);
  nand (_26910_, _24467_, _23379_);
  and (_26911_, _26910_, _26437_);
  and (_26912_, _26911_, _26909_);
  or (_26913_, _26912_, _26908_);
  or (_26914_, _26913_, _26904_);
  or (_26915_, _26914_, _26900_);
  and (_26916_, _26915_, _26368_);
  or (_26917_, _26916_, _26896_);
  or (_26918_, _26917_, _26890_);
  and (_26919_, _26445_, ABINPUT[3]);
  and (_26920_, _26443_, ABINPUT[5]);
  or (_26921_, _26920_, _26919_);
  and (_26922_, _26921_, _24467_);
  nor (_26923_, _24467_, _23293_);
  and (_26924_, _24467_, ABINPUT[4]);
  or (_26925_, _26924_, _26923_);
  and (_26926_, _26925_, _26440_);
  nand (_26927_, _24467_, _23519_);
  or (_26928_, _24467_, ABINPUT[10]);
  and (_26929_, _26928_, _26927_);
  and (_26930_, _26929_, _26437_);
  or (_26931_, _26930_, _26926_);
  and (_26932_, _26445_, ABINPUT[7]);
  and (_26933_, _26443_, ABINPUT[9]);
  or (_26934_, _26933_, _26932_);
  and (_26935_, _26934_, _26436_);
  or (_26936_, _26935_, _26931_);
  nor (_26937_, _26936_, _26922_);
  nand (_26938_, _26937_, _26896_);
  and (_26939_, _26938_, _25964_);
  and (_01520_, _26939_, _26918_);
  and (_26940_, _26445_, _24467_);
  and (_26941_, _26940_, _26367_);
  and (_26942_, _26941_, _23310_);
  not (_26943_, _23241_);
  and (_26944_, _24511_, _24467_);
  and (_26945_, _26944_, _26445_);
  and (_26946_, _26945_, _26371_);
  and (_26947_, _26946_, _26943_);
  nor (_26948_, _26947_, _26942_);
  and (_26949_, _26944_, _26437_);
  and (_26950_, _26949_, _26383_);
  and (_26951_, _26950_, _23141_);
  not (_26953_, _26951_);
  and (_26955_, _26953_, _26948_);
  nor (_26957_, _26955_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_26959_, _26957_);
  nor (_26961_, _22615_, _16205_);
  and (_26963_, _26961_, _26432_);
  not (_26965_, _26963_);
  and (_26967_, _26437_, _26436_);
  not (_26969_, _26967_);
  and (_26971_, _26969_, _23385_);
  and (_26973_, _26971_, _26420_);
  and (_26975_, _26940_, _26368_);
  nor (_26977_, _26975_, _26973_);
  and (_26979_, _26977_, _26965_);
  and (_26981_, _26979_, _26959_);
  and (_26983_, _26944_, _26443_);
  and (_26985_, _26983_, _26383_);
  and (_26987_, _26985_, _23141_);
  or (_26989_, _26987_, rst);
  nor (_01522_, _26989_, _26981_);
  not (_26992_, _26987_);
  and (_26994_, _26940_, _26391_);
  and (_26996_, _26994_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_26998_, _26985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or (_27000_, _26998_, _26996_);
  and (_27002_, _26940_, _24512_);
  and (_27004_, _27002_, _26383_);
  and (_27006_, _27004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_27008_, _27002_, _26381_);
  and (_27010_, _27008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_27012_, _27010_, _27006_);
  or (_27013_, _27012_, _27000_);
  and (_27014_, _26940_, _26396_);
  and (_27015_, _27014_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_27016_, _26950_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_27017_, _27016_, _27015_);
  and (_27018_, _26945_, _26386_);
  and (_27019_, _27018_, _26822_);
  not (_27020_, _23072_);
  and (_27021_, _26944_, _26440_);
  and (_27022_, _27021_, _26383_);
  and (_27023_, _27022_, _27020_);
  or (_27024_, _27023_, _27019_);
  or (_27025_, _27024_, _27017_);
  or (_27026_, _27025_, _27013_);
  and (_27027_, _26941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_27028_, _26945_, _26381_);
  and (_27029_, _27028_, _26636_);
  and (_27030_, _26945_, _26375_);
  and (_27031_, _27030_, _26757_);
  or (_27032_, _27031_, _27029_);
  and (_27033_, _26946_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_27034_, _26945_, _26383_);
  and (_27035_, _27034_, _26545_);
  or (_27036_, _27035_, _27033_);
  or (_27037_, _27036_, _27032_);
  or (_27038_, _27037_, _27027_);
  nor (_27039_, _27038_, _27026_);
  and (_27040_, _26969_, _26420_);
  and (_27041_, _27040_, _23385_);
  not (_27042_, _27041_);
  and (_27043_, _26941_, _23313_);
  and (_27044_, _26432_, _17151_);
  and (_27045_, _27044_, _16216_);
  nor (_27046_, _27045_, _27043_);
  and (_27047_, _27046_, _27042_);
  and (_27048_, _27047_, _26959_);
  and (_27049_, _27048_, _27039_);
  nor (_27050_, _27048_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_27051_, _27050_, _27049_);
  nand (_27052_, _27051_, _26992_);
  nand (_27053_, _26987_, _17086_);
  and (_27054_, _27053_, _25964_);
  and (_01524_, _27054_, _27052_);
  nor (_01527_, _24391_, rst);
  and (_27055_, _26994_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_27056_, _26985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or (_27057_, _27056_, _27055_);
  and (_27058_, _27004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_27059_, _27008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_27060_, _27059_, _27058_);
  or (_27061_, _27060_, _27057_);
  and (_27062_, _27014_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_27063_, _26950_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_27064_, _27063_, _27062_);
  and (_27065_, _27018_, _26845_);
  and (_27066_, _27022_, _24543_);
  or (_27067_, _27066_, _27065_);
  or (_27068_, _27067_, _27064_);
  or (_27069_, _27068_, _27061_);
  and (_27070_, _26941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_27071_, _27028_, _26620_);
  and (_27072_, _27030_, _26789_);
  or (_27073_, _27072_, _27071_);
  and (_27074_, _27034_, _26561_);
  and (_27075_, _26946_, _26688_);
  or (_27076_, _27075_, _27074_);
  or (_27077_, _27076_, _27073_);
  or (_27078_, _27077_, _27070_);
  nor (_27079_, _27078_, _27069_);
  nand (_27080_, _27079_, _26981_);
  or (_27081_, _26981_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_27082_, _27081_, _27080_);
  or (_27083_, _27082_, _26987_);
  nand (_27084_, _26987_, _23162_);
  and (_27085_, _27084_, _25964_);
  and (_02203_, _27085_, _27083_);
  and (_27086_, _26994_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_27087_, _26985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or (_27088_, _27087_, _27086_);
  and (_27089_, _27004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_27090_, _27008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_27091_, _27090_, _27089_);
  or (_27092_, _27091_, _27088_);
  and (_27094_, _27014_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_27095_, _26950_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_27096_, _27095_, _27094_);
  and (_27097_, _27018_, _26878_);
  and (_27098_, _27022_, _24646_);
  or (_27099_, _27098_, _27097_);
  or (_27100_, _27099_, _27096_);
  or (_27101_, _27100_, _27092_);
  and (_27102_, _26941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_27103_, _27028_, _26604_);
  and (_27104_, _27030_, _26767_);
  or (_27106_, _27104_, _27103_);
  and (_27107_, _26946_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_27108_, _27034_, _26529_);
  or (_27109_, _27108_, _27107_);
  or (_27110_, _27109_, _27106_);
  or (_27111_, _27110_, _27102_);
  nor (_27112_, _27111_, _27101_);
  and (_27113_, _27112_, _27048_);
  nor (_27114_, _27048_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or (_27115_, _27114_, _27113_);
  nand (_27116_, _27115_, _26992_);
  nand (_27117_, _26987_, _17475_);
  and (_27118_, _27117_, _25964_);
  and (_02205_, _27118_, _27116_);
  and (_27119_, _26985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_27120_, _26994_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_27121_, _27120_, _27119_);
  and (_27122_, _27004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_27123_, _27008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_27124_, _27123_, _27122_);
  or (_27125_, _27124_, _27121_);
  and (_27126_, _27014_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_27127_, _26950_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_27128_, _27127_, _27126_);
  and (_27129_, _27018_, _26861_);
  and (_27130_, _27022_, _24462_);
  or (_27131_, _27130_, _27129_);
  or (_27132_, _27131_, _27128_);
  or (_27133_, _27132_, _27125_);
  and (_27134_, _26941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_27136_, _27028_, _26581_);
  and (_27137_, _27030_, _26782_);
  or (_27138_, _27137_, _27136_);
  and (_27139_, _27034_, _26520_);
  and (_27140_, _26946_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_27141_, _27140_, _27139_);
  or (_27142_, _27141_, _27138_);
  or (_27143_, _27142_, _27134_);
  nor (_27144_, _27143_, _27133_);
  nand (_27145_, _27144_, _26981_);
  or (_27146_, _26981_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_27147_, _27146_, _27145_);
  or (_27148_, _27147_, _26987_);
  nand (_27149_, _26987_, _17670_);
  and (_27150_, _27149_, _25964_);
  and (_02207_, _27150_, _27148_);
  and (_27151_, _26994_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_27152_, _26985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_27153_, _27152_, _27151_);
  and (_27154_, _27004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_27156_, _27008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_27157_, _27156_, _27154_);
  or (_27158_, _27157_, _27153_);
  and (_27159_, _27014_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_27160_, _26950_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_27161_, _27160_, _27159_);
  and (_27162_, _27018_, _26871_);
  and (_27163_, _27022_, _24495_);
  or (_27164_, _27163_, _27162_);
  or (_27165_, _27164_, _27161_);
  or (_27166_, _27165_, _27158_);
  and (_27167_, _26941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_27168_, _27028_, _26629_);
  and (_27169_, _27030_, _26774_);
  or (_27170_, _27169_, _27168_);
  and (_27171_, _26946_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_27172_, _27034_, _26552_);
  or (_27173_, _27172_, _27171_);
  or (_27174_, _27173_, _27170_);
  or (_27175_, _27174_, _27167_);
  nor (_27176_, _27175_, _27166_);
  and (_27177_, _27176_, _27048_);
  nor (_27178_, _27048_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or (_27179_, _27178_, _27177_);
  nand (_27180_, _27179_, _26992_);
  nand (_27181_, _26987_, _17845_);
  and (_27182_, _27181_, _25964_);
  and (_02209_, _27182_, _27180_);
  and (_27183_, _26994_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_27184_, _26985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  or (_27185_, _27184_, _27183_);
  and (_27186_, _27004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_27187_, _27008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_27188_, _27187_, _27186_);
  or (_27189_, _27188_, _27185_);
  and (_27190_, _27014_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_27191_, _26950_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_27192_, _27191_, _27190_);
  and (_27193_, _27018_, _26838_);
  and (_27194_, _27022_, _24617_);
  or (_27195_, _27194_, _27193_);
  or (_27196_, _27195_, _27192_);
  or (_27197_, _27196_, _27189_);
  and (_27198_, _26941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_27199_, _27028_, _26613_);
  and (_27200_, _27030_, _26735_);
  or (_27201_, _27200_, _27199_);
  and (_27202_, _26946_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_27203_, _27034_, _26568_);
  or (_27204_, _27203_, _27202_);
  or (_27205_, _27204_, _27201_);
  or (_27206_, _27205_, _27198_);
  nor (_27207_, _27206_, _27197_);
  and (_27208_, _27207_, _27048_);
  nor (_27209_, _27048_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or (_27210_, _27209_, _27208_);
  nand (_27211_, _27210_, _26992_);
  nand (_27212_, _26987_, _18019_);
  and (_27213_, _27212_, _25964_);
  and (_02211_, _27213_, _27211_);
  and (_27214_, _26994_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_27215_, _26985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_27216_, _27215_, _27214_);
  and (_27217_, _27004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_27218_, _27008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_27219_, _27218_, _27217_);
  or (_27220_, _27219_, _27216_);
  and (_27221_, _27014_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_27222_, _26950_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_27223_, _27222_, _27221_);
  and (_27224_, _27018_, _26829_);
  not (_27225_, _23133_);
  and (_27226_, _27022_, _27225_);
  or (_27227_, _27226_, _27224_);
  or (_27228_, _27227_, _27223_);
  or (_27229_, _27228_, _27220_);
  and (_27230_, _26941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_27231_, _27028_, _26597_);
  and (_27232_, _27030_, _26750_);
  or (_27233_, _27232_, _27231_);
  and (_27234_, _26946_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_27235_, _27034_, _26536_);
  or (_27236_, _27235_, _27234_);
  or (_27237_, _27236_, _27233_);
  or (_27238_, _27237_, _27230_);
  nor (_27239_, _27238_, _27229_);
  and (_27240_, _27239_, _27048_);
  nor (_27241_, _27048_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or (_27242_, _27241_, _27240_);
  nand (_27243_, _27242_, _26992_);
  nand (_27244_, _26987_, _18194_);
  and (_27245_, _27244_, _25964_);
  and (_02213_, _27245_, _27243_);
  and (_27246_, _26994_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_27247_, _26985_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_27248_, _27247_, _27246_);
  and (_27249_, _27004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_27250_, _27008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_27251_, _27250_, _27249_);
  or (_27252_, _27251_, _27248_);
  and (_27253_, _27014_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_27254_, _26950_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_27255_, _27254_, _27253_);
  and (_27256_, _27018_, _26854_);
  and (_27257_, _27022_, _24570_);
  or (_27258_, _27257_, _27256_);
  or (_27259_, _27258_, _27255_);
  or (_27260_, _27259_, _27252_);
  and (_27261_, _26941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_27262_, _27028_, _26588_);
  and (_27263_, _27030_, _26742_);
  or (_27264_, _27263_, _27262_);
  and (_27265_, _26946_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_27266_, _27034_, _26513_);
  or (_27267_, _27266_, _27265_);
  or (_27268_, _27267_, _27264_);
  or (_27269_, _27268_, _27261_);
  nor (_27270_, _27269_, _27260_);
  and (_27271_, _27270_, _27048_);
  nor (_27272_, _27048_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or (_27273_, _27272_, _27271_);
  nand (_27274_, _27273_, _26992_);
  nand (_27275_, _26987_, _18368_);
  and (_27276_, _27275_, _25964_);
  and (_02215_, _27276_, _27274_);
  or (_27277_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_27278_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_27279_, _26505_, _27278_);
  and (_27280_, _27279_, _25964_);
  and (_02771_, _27280_, _27277_);
  and (_27281_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_27282_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  or (_27283_, _27282_, _27281_);
  and (_02775_, _27283_, _25964_);
  nor (_03153_, _24377_, rst);
  nor (_03160_, _24637_, rst);
  nor (_03164_, _24368_, rst);
  and (_27284_, \oc8051_top_1.oc8051_decoder1.state [0], _15520_);
  nor (_27285_, _21476_, _27284_);
  nor (_27286_, _22615_, _16988_);
  and (_27287_, _27286_, _27285_);
  and (_27288_, _27287_, _26420_);
  nor (_27289_, _27285_, _20774_);
  nor (_27290_, _27289_, _20982_);
  nand (_27291_, _27290_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_27292_, ABINPUT[28], ABINPUT[27]);
  nor (_27293_, ABINPUT[30], ABINPUT[29]);
  and (_27294_, _27293_, _27292_);
  nor (_27295_, ABINPUT[32], ABINPUT[31]);
  nor (_27296_, ABINPUT[33], ABINPUT[34]);
  and (_27297_, _27296_, _27295_);
  and (_27298_, _27297_, _27294_);
  nor (_27299_, _27285_, _20971_);
  and (_27300_, _27299_, _27298_);
  nor (_27301_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_27302_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_27303_, _27302_, _27301_);
  nor (_27304_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_27305_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_27306_, _27305_, _27304_);
  and (_27307_, _27306_, _27303_);
  and (_27308_, _27307_, _22528_);
  nor (_27309_, _27308_, _27300_);
  and (_27310_, _27309_, _27291_);
  not (_27311_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_27312_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _27311_);
  and (_27313_, _24793_, _24789_);
  and (_27314_, _24804_, _24801_);
  nor (_27315_, _27314_, _27313_);
  and (_27316_, _24819_, _24817_);
  and (_27317_, _24835_, _24834_);
  nor (_27318_, _27317_, _27316_);
  and (_27319_, _27318_, _27315_);
  and (_27320_, _24876_, _24875_);
  and (_27321_, _24848_, _24847_);
  nor (_27322_, _27321_, _27320_);
  and (_27323_, _24767_, _24766_);
  and (_27324_, _24862_, _24861_);
  nor (_27325_, _27324_, _27323_);
  and (_27326_, _27325_, _27322_);
  and (_27327_, _27326_, _27319_);
  nor (_27328_, _27327_, _27312_);
  and (_27329_, _27312_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_27330_, _27329_, _27328_);
  not (_27331_, _27330_);
  and (_27332_, _27331_, _27285_);
  not (_27333_, _27332_);
  and (_27334_, _27333_, _27310_);
  and (_27335_, _20960_, _19475_);
  nor (_27336_, _27335_, _22101_);
  or (_27337_, _27336_, _27334_);
  and (_27338_, _20949_, _20993_);
  nor (_27339_, _27338_, _20850_);
  not (_27340_, _27339_);
  and (_27341_, _26480_, _21311_);
  not (_27342_, _27341_);
  and (_27343_, _26492_, _21783_);
  nor (_27344_, _27343_, _21837_);
  and (_27345_, _27344_, _27342_);
  and (_27346_, _22221_, _21508_);
  and (_27347_, _26480_, _21508_);
  nor (_27348_, _27347_, _27346_);
  and (_27349_, _27348_, _27345_);
  or (_27350_, _20840_, _21421_);
  or (_27351_, _27350_, _21190_);
  and (_27352_, _27351_, _20949_);
  not (_27353_, _27352_);
  and (_27354_, _27353_, _27349_);
  not (_27355_, _27354_);
  and (_27356_, _27355_, _27334_);
  nor (_27357_, _27356_, _27340_);
  and (_27358_, _27357_, _27337_);
  nor (_27359_, _27358_, _24389_);
  and (_27360_, _21245_, _20719_);
  and (_27361_, _21432_, _21147_);
  nor (_27362_, _27361_, _27360_);
  nor (_27363_, _27362_, _18477_);
  nor (_27364_, _27363_, _22123_);
  not (_27365_, _27364_);
  nor (_27366_, _27365_, _27359_);
  not (_27367_, _22528_);
  nor (_27368_, _23337_, _23326_);
  nor (_27369_, _27368_, _27367_);
  not (_27370_, _23235_);
  nor (_27371_, _23248_, _26943_);
  and (_27372_, _27371_, _27370_);
  not (_27373_, _27372_);
  and (_27374_, _27373_, _27290_);
  nor (_27375_, _27374_, _27369_);
  not (_27376_, _27375_);
  nor (_27377_, _27376_, _27366_);
  not (_27378_, _27377_);
  nor (_27379_, _27378_, _27288_);
  and (_27380_, _27379_, _26965_);
  nor (_27381_, _22134_, rst);
  and (_03173_, _27381_, _27380_);
  and (_03177_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _25964_);
  and (_03180_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _25964_);
  and (_27383_, _20850_, _20916_);
  nor (_27384_, _27383_, _27363_);
  nor (_27385_, _24389_, _21476_);
  and (_27386_, _21388_, _24378_);
  nor (_27387_, _27386_, _27385_);
  and (_27389_, _27348_, _27344_);
  nor (_27390_, _27389_, _24389_);
  and (_27391_, _20905_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_27392_, _27391_, _21574_);
  and (_27393_, _27361_, _24378_);
  nor (_27395_, _27393_, _27392_);
  not (_27396_, _27395_);
  nor (_27397_, _27396_, _27390_);
  and (_27398_, _27397_, _27387_);
  and (_27399_, _27349_, _27339_);
  nor (_27401_, _27399_, _24389_);
  not (_27402_, _27401_);
  and (_27403_, _27387_, _20982_);
  and (_27404_, _27403_, _27402_);
  and (_27405_, _27404_, _27398_);
  and (_27407_, _27405_, _27384_);
  and (_27408_, _27407_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_27409_, _27393_, _24336_);
  and (_27410_, _27392_, ABINPUT[26]);
  or (_27411_, _27410_, _27409_);
  or (_27413_, _27411_, _27408_);
  and (_27414_, _27398_, _24336_);
  nor (_27415_, _27398_, _26244_);
  nor (_27416_, _27415_, _27414_);
  not (_27417_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_27419_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_27420_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_27422_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_27423_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_27424_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not (_27425_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_27426_, _27416_, _27425_);
  and (_27427_, _27416_, _27425_);
  not (_27428_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_27430_, _27398_, _24587_);
  nor (_27431_, _27398_, _26363_);
  nor (_27432_, _27431_, _27430_);
  nor (_27434_, _27432_, _27428_);
  and (_27435_, _27432_, _27428_);
  nor (_27436_, _27435_, _27434_);
  not (_27438_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_27439_, _27398_, _24421_);
  nor (_27440_, _27398_, _26346_);
  nor (_27442_, _27440_, _27439_);
  nor (_27443_, _27442_, _27438_);
  and (_27444_, _27442_, _27438_);
  not (_27446_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_27447_, _27398_, _24634_);
  nor (_27448_, _27398_, _26329_);
  nor (_27450_, _27448_, _27447_);
  or (_27451_, _27450_, _27446_);
  not (_27452_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_27454_, _27398_, _24492_);
  nor (_27455_, _27398_, _26312_);
  nor (_27457_, _27455_, _27454_);
  nor (_27458_, _27457_, _27452_);
  and (_27459_, _27457_, _27452_);
  not (_27460_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_27461_, _27398_, _24447_);
  nor (_27462_, _27398_, _26295_);
  nor (_27463_, _27462_, _27461_);
  nor (_27465_, _27463_, _27460_);
  not (_27466_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_27467_, _27398_, _24676_);
  nor (_27469_, _27398_, _26278_);
  nor (_27470_, _27469_, _27467_);
  nor (_27471_, _27470_, _27466_);
  not (_27473_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_27474_, _27398_, _24528_);
  nor (_27475_, _27398_, _26261_);
  nor (_27477_, _27475_, _27474_);
  nor (_27478_, _27477_, _27473_);
  and (_27479_, _27470_, _27466_);
  nor (_27481_, _27479_, _27471_);
  and (_27482_, _27481_, _27478_);
  nor (_27483_, _27482_, _27471_);
  not (_27485_, _27483_);
  and (_27486_, _27463_, _27460_);
  nor (_27487_, _27486_, _27465_);
  and (_27489_, _27487_, _27485_);
  nor (_27490_, _27489_, _27465_);
  nor (_27492_, _27490_, _27459_);
  or (_27493_, _27492_, _27458_);
  nand (_27494_, _27450_, _27446_);
  and (_27495_, _27494_, _27451_);
  nand (_27496_, _27495_, _27493_);
  and (_27498_, _27496_, _27451_);
  nor (_27499_, _27498_, _27444_);
  or (_27500_, _27499_, _27443_);
  and (_27502_, _27500_, _27436_);
  nor (_27503_, _27502_, _27434_);
  nor (_27504_, _27503_, _27427_);
  or (_27506_, _27504_, _27426_);
  nor (_27507_, _27506_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_27508_, _27507_, _27424_);
  and (_27510_, _27508_, _27423_);
  and (_27511_, _27510_, _27422_);
  and (_27512_, _27511_, _27420_);
  and (_27514_, _27512_, _27419_);
  and (_27515_, _27514_, _27417_);
  nor (_27516_, _27515_, _27416_);
  not (_27518_, _27416_);
  and (_27519_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_27520_, _27519_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_27522_, _27520_, _27506_);
  and (_27523_, _27522_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_27525_, _27523_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_27526_, _27525_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_27527_, _27526_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_27528_, _27527_, _27518_);
  nor (_27529_, _27528_, _27516_);
  or (_27530_, _27529_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_27531_, _27529_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_27533_, _27531_, _27530_);
  not (_27534_, _27384_);
  and (_27535_, _27534_, _27398_);
  not (_27537_, _27348_);
  nor (_27538_, _27537_, _20960_);
  and (_27539_, _27538_, _27339_);
  and (_27541_, _27539_, _27345_);
  nor (_27542_, _27541_, _24389_);
  and (_27543_, _21366_, _19732_);
  and (_27545_, _27543_, _20949_);
  not (_27546_, _27545_);
  and (_27547_, _24388_, _27546_);
  nor (_27549_, _24389_, _27547_);
  and (_27550_, _20949_, _24378_);
  and (_27551_, _27550_, _21377_);
  nor (_27553_, _27551_, _27549_);
  not (_27554_, _27553_);
  nor (_27555_, _27554_, _27542_);
  nor (_27557_, _27555_, _27535_);
  and (_27558_, _27557_, _27533_);
  or (_27560_, _27558_, _27413_);
  and (_27561_, _27383_, ABINPUT[18]);
  and (_27562_, _27555_, _27535_);
  and (_27563_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_27565_, _27563_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_27566_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_27567_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_27569_, _27567_, _27566_);
  and (_27570_, _27569_, _27565_);
  and (_27571_, _27570_, _27520_);
  and (_27573_, _27571_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_27574_, _27573_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_27575_, _27574_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_27577_, _27575_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_27578_, _27577_, _27278_);
  and (_27579_, _27577_, _27278_);
  or (_27581_, _27579_, _27578_);
  and (_27582_, _27581_, _27562_);
  nor (_27583_, _27582_, _27561_);
  nand (_27585_, _27583_, _27380_);
  or (_27586_, _27585_, _27560_);
  and (_27587_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_27589_, _18685_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_27590_, _27589_, _24319_);
  nor (_27592_, _27590_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_27593_, _27592_);
  and (_27594_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_27595_, _27594_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_27597_, _27595_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_27598_, _27597_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_27599_, _27598_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_27601_, _27599_, _27593_);
  and (_27602_, _27601_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_27603_, _27602_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_27605_, _27603_, _27587_);
  and (_27606_, _27605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_27607_, _27606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_27609_, _27607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_27610_, _27609_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_27611_, _27609_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_27613_, _27611_, _27610_);
  or (_27614_, _27613_, _27380_);
  and (_27615_, _27614_, _25964_);
  and (_03183_, _27615_, _27586_);
  and (_27617_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _25964_);
  and (_27618_, _27617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_27620_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_27621_, _18521_, _27620_);
  not (_27623_, _27621_);
  not (_27624_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_27625_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_27626_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_27628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_27629_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_27630_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_27632_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_27633_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_27634_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_27636_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_27637_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_27638_, _27637_, _27636_);
  and (_27640_, _27638_, _27634_);
  and (_27641_, _27640_, _27633_);
  and (_27642_, _27641_, _27632_);
  and (_27644_, _27642_, _27630_);
  and (_27645_, _27644_, _27629_);
  and (_27646_, _27645_, _27628_);
  and (_27648_, _27646_, _27626_);
  and (_27649_, _27648_, _27625_);
  nor (_27650_, _27649_, _27624_);
  and (_27652_, _27649_, _27624_);
  nor (_27653_, _27652_, _27650_);
  not (_27655_, _27653_);
  and (_27656_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_27657_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_27658_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_27659_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_27660_, _27659_, _27657_);
  and (_27661_, _27660_, _27658_);
  nor (_27663_, _27661_, _27657_);
  nor (_27664_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_27665_, _27664_, _27656_);
  not (_27667_, _27665_);
  nor (_27668_, _27667_, _27663_);
  nor (_27669_, _27668_, _27656_);
  and (_27671_, _27669_, _27648_);
  nor (_27672_, _27671_, _27625_);
  and (_27673_, _27669_, _27649_);
  nor (_27675_, _27673_, _27672_);
  not (_27676_, _27675_);
  and (_27677_, _27669_, _27646_);
  nor (_27679_, _27677_, _27626_);
  nor (_27680_, _27679_, _27671_);
  not (_27681_, _27680_);
  and (_27683_, _27669_, _27645_);
  and (_27684_, _27669_, _27642_);
  and (_27685_, _27684_, _27630_);
  nor (_27687_, _27685_, _27629_);
  nor (_27688_, _27687_, _27683_);
  not (_27690_, _27688_);
  nor (_27691_, _27684_, _27630_);
  or (_27692_, _27691_, _27685_);
  not (_27693_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_27695_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_27696_, _27669_, _27641_);
  and (_27697_, _27696_, _27695_);
  nor (_27699_, _27697_, _27693_);
  nor (_27700_, _27699_, _27684_);
  not (_27701_, _27700_);
  and (_27703_, _27669_, _27638_);
  and (_27704_, _27703_, _27634_);
  nor (_27705_, _27704_, _27633_);
  nor (_27707_, _27705_, _27696_);
  not (_27708_, _27707_);
  nor (_27709_, _27703_, _27634_);
  or (_27711_, _27709_, _27704_);
  nand (_27712_, _27669_, _27637_);
  and (_27713_, _27712_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_27715_, _27713_, _27703_);
  not (_27716_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_27717_, _27669_, _27716_);
  nor (_27721_, _27669_, _27716_);
  nor (_27722_, _27721_, _27717_);
  not (_27730_, _27722_);
  not (_27731_, _18905_);
  and (_27738_, _19135_, _27731_);
  nor (_27746_, _19699_, _19442_);
  and (_27748_, _27746_, _27738_);
  not (_27749_, _27748_);
  and (_27762_, _20686_, _20445_);
  and (_27767_, _27762_, _20214_);
  not (_27768_, _20445_);
  not (_27775_, _20214_);
  and (_27784_, _20686_, _27775_);
  and (_27785_, _27784_, _27768_);
  nor (_27793_, _27785_, _27767_);
  nor (_27795_, _27793_, _27749_);
  not (_27796_, _19962_);
  and (_27804_, _27785_, _27796_);
  not (_27813_, _19699_);
  and (_27814_, _19135_, _18905_);
  and (_27821_, _27814_, _27813_);
  and (_27826_, _27821_, _27804_);
  nor (_27827_, _27826_, _27795_);
  not (_27840_, _19135_);
  and (_27846_, _27840_, _18905_);
  and (_27847_, _27846_, _27746_);
  and (_27859_, _27813_, _19442_);
  and (_27860_, _27859_, _27738_);
  nor (_27867_, _27860_, _27847_);
  nor (_27876_, _27867_, _20686_);
  and (_27885_, _27785_, _19962_);
  not (_27886_, _27885_);
  and (_27894_, _19699_, _19442_);
  and (_27903_, _27894_, _27846_);
  nor (_27904_, _27903_, _27860_);
  nor (_27912_, _27904_, _27886_);
  nor (_27918_, _27912_, _27876_);
  and (_27919_, _27918_, _27827_);
  and (_27933_, _27767_, _19962_);
  not (_27940_, _19442_);
  and (_27941_, _19699_, _27940_);
  and (_27953_, _27941_, _27846_);
  and (_27958_, _27953_, _27933_);
  and (_27959_, _27814_, _19699_);
  and (_27967_, _27959_, _27804_);
  nor (_27969_, _27967_, _27958_);
  not (_27970_, _27933_);
  nor (_27971_, _19135_, _18905_);
  and (_27973_, _27971_, _27894_);
  nor (_27974_, _27973_, _27860_);
  nor (_27976_, _27974_, _27970_);
  and (_27977_, _27821_, _27885_);
  nor (_27978_, _27977_, _27976_);
  and (_27979_, _27978_, _27969_);
  and (_27980_, _27979_, _27919_);
  and (_27982_, _27767_, _27796_);
  and (_27983_, _27941_, _27738_);
  and (_27984_, _27983_, _27982_);
  and (_27986_, _27775_, _19962_);
  and (_27987_, _27986_, _27762_);
  and (_27988_, _27987_, _27903_);
  nor (_27990_, _27988_, _27984_);
  not (_27991_, _27990_);
  and (_27992_, _27859_, _27846_);
  and (_27994_, _27992_, _27804_);
  and (_27995_, _27894_, _27738_);
  and (_27996_, _27995_, _27982_);
  or (_27998_, _27996_, _27994_);
  nor (_27999_, _27998_, _27991_);
  or (_28000_, _27903_, _27847_);
  and (_28002_, _28000_, _27933_);
  not (_28003_, _27987_);
  and (_28004_, _27971_, _19699_);
  nor (_28006_, _28004_, _27847_);
  nor (_28007_, _28006_, _28003_);
  nor (_28009_, _28007_, _28002_);
  not (_28010_, _27804_);
  and (_28011_, _27971_, _27941_);
  nor (_28012_, _28011_, _27903_);
  nor (_28014_, _28012_, _28010_);
  nor (_28015_, _28011_, _27992_);
  nor (_28016_, _28015_, _27970_);
  nor (_28018_, _28016_, _28014_);
  and (_28019_, _28018_, _28009_);
  and (_28020_, _28019_, _27999_);
  and (_28022_, _28020_, _27980_);
  nor (_28023_, _27933_, _27785_);
  not (_28024_, _28023_);
  and (_28026_, _28024_, _27983_);
  and (_28027_, _27971_, _27813_);
  and (_28028_, _28027_, _27804_);
  nor (_28030_, _28028_, _28026_);
  not (_28031_, _27814_);
  or (_28032_, _27859_, _28031_);
  nor (_28034_, _28032_, _27941_);
  and (_28035_, _28034_, _27987_);
  and (_28036_, _27973_, _27804_);
  nor (_28038_, _28036_, _28035_);
  and (_28039_, _27959_, _27933_);
  not (_28041_, _28039_);
  or (_28042_, _27953_, _27860_);
  and (_28043_, _28042_, _27804_);
  and (_28044_, _27992_, _27885_);
  nor (_28046_, _28044_, _28043_);
  and (_28047_, _28046_, _28041_);
  and (_28048_, _28047_, _28038_);
  and (_28050_, _27738_, _27813_);
  and (_28051_, _27987_, _28050_);
  not (_28052_, _28051_);
  and (_28054_, _27846_, _27940_);
  nor (_28055_, _20445_, _27775_);
  and (_28056_, _28055_, _20686_);
  and (_28058_, _28056_, _28054_);
  nor (_28059_, _20214_, _19962_);
  and (_28060_, _28059_, _27762_);
  nor (_28062_, _28060_, _28058_);
  and (_28063_, _28062_, _28052_);
  and (_28064_, _27992_, _27987_);
  or (_28066_, _27846_, _27738_);
  and (_28067_, _28066_, _27859_);
  and (_28068_, _28067_, _28056_);
  nor (_28070_, _28068_, _28064_);
  and (_28071_, _28070_, _28063_);
  nor (_28073_, _27992_, _27953_);
  nor (_28074_, _28073_, _20686_);
  and (_28075_, _27995_, _27987_);
  and (_28076_, _27859_, _27814_);
  and (_28078_, _28076_, _27987_);
  nor (_28079_, _28078_, _28075_);
  not (_28080_, _28079_);
  nor (_28082_, _28080_, _28074_);
  and (_28083_, _28082_, _28071_);
  and (_28084_, _28024_, _27995_);
  not (_28086_, _28084_);
  and (_28087_, _27987_, _27953_);
  not (_28088_, _28087_);
  and (_28090_, _27987_, _27983_);
  not (_28091_, _20686_);
  and (_28092_, _27973_, _28091_);
  nor (_28094_, _28092_, _28090_);
  and (_28095_, _28094_, _28088_);
  and (_28096_, _28095_, _28086_);
  and (_28098_, _28096_, _28083_);
  and (_28099_, _28098_, _28048_);
  and (_28100_, _28099_, _28030_);
  and (_28102_, _28100_, _28022_);
  not (_28103_, _28102_);
  nor (_28104_, _27660_, _27658_);
  nor (_28105_, _28104_, _27661_);
  nand (_28106_, _28105_, _28103_);
  and (_28107_, _27982_, _27748_);
  or (_28108_, _28055_, _28091_);
  and (_28109_, _28108_, _27992_);
  or (_28110_, _28109_, _28078_);
  nor (_28111_, _28110_, _28107_);
  and (_28112_, _28111_, _27999_);
  nand (_28113_, _28112_, _28048_);
  nor (_28114_, _28113_, _28102_);
  not (_28115_, _28114_);
  nor (_28116_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_28117_, _28116_, _27658_);
  and (_28118_, _28117_, _28115_);
  or (_28119_, _28105_, _28103_);
  and (_28120_, _28119_, _28106_);
  nand (_28121_, _28120_, _28118_);
  and (_28122_, _28121_, _28106_);
  not (_28123_, _28122_);
  and (_28124_, _27667_, _27663_);
  nor (_28125_, _28124_, _27668_);
  and (_28126_, _28125_, _28123_);
  and (_28127_, _28126_, _27730_);
  not (_28128_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_28129_, _27717_, _28128_);
  nand (_28130_, _28129_, _27712_);
  and (_28131_, _28130_, _28127_);
  and (_28132_, _28131_, _27715_);
  and (_28133_, _28132_, _27711_);
  and (_28134_, _28133_, _27708_);
  nor (_28135_, _27696_, _27695_);
  or (_28136_, _28135_, _27697_);
  and (_28137_, _28136_, _28134_);
  and (_28138_, _28137_, _27701_);
  and (_28139_, _28138_, _27692_);
  and (_28140_, _28139_, _27690_);
  nor (_28141_, _27683_, _27628_);
  or (_28142_, _28141_, _27677_);
  and (_28143_, _28142_, _28140_);
  and (_28144_, _28143_, _27681_);
  and (_28145_, _28144_, _27676_);
  not (_28146_, _27669_);
  and (_28147_, _28146_, _27649_);
  nor (_28148_, _28147_, _28145_);
  nor (_28149_, _28148_, _27655_);
  and (_28150_, _28148_, _27655_);
  or (_28151_, _28150_, _28149_);
  or (_28152_, _28151_, _27623_);
  or (_28153_, _27621_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_28154_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_28155_, _28154_, _28153_);
  and (_28156_, _28155_, _28152_);
  or (_03186_, _28156_, _27618_);
  nor (_28157_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_03191_, _28157_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_03194_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _25964_);
  nor (_28158_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_28159_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_28160_, _28159_, _28158_);
  nor (_28161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_28162_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_28163_, _28162_, _28161_);
  and (_28164_, _28163_, _28160_);
  nor (_28165_, _28164_, rst);
  and (_28166_, \oc8051_top_1.oc8051_rom1.ea_int , _18488_);
  nand (_28167_, _28166_, _18521_);
  and (_28168_, _28167_, _03194_);
  or (_03197_, _28168_, _28165_);
  and (_28169_, _28164_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_28170_, _28169_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_03200_, _28170_, _25964_);
  nor (_28171_, _27592_, _24319_);
  or (_28172_, _28102_, _18631_);
  nor (_28173_, _28114_, _18718_);
  nand (_28174_, _28102_, _18631_);
  and (_28175_, _28174_, _28172_);
  nand (_28176_, _28175_, _28173_);
  and (_28177_, _28176_, _28172_);
  nor (_28178_, _28177_, _24319_);
  and (_28179_, _28178_, _18620_);
  nor (_28180_, _28178_, _18620_);
  nor (_28181_, _28180_, _28179_);
  nor (_28182_, _28181_, _28171_);
  and (_28183_, _18642_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_28184_, _28183_, _28171_);
  and (_28185_, _28184_, _28113_);
  or (_28186_, _28185_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_28187_, _28186_, _28182_);
  and (_03202_, _28187_, _25964_);
  not (_28188_, _20148_);
  and (_28189_, _28188_, _18839_);
  not (_28190_, _19366_);
  and (_28191_, _19091_, _28190_);
  and (_28192_, _28191_, _28189_);
  and (_28193_, _18521_, _25964_);
  and (_28194_, _28193_, _18510_);
  nand (_28195_, _28194_, _20401_);
  nor (_28196_, _28195_, _20642_);
  not (_28197_, _19918_);
  and (_28198_, _28197_, _19655_);
  and (_28199_, _28198_, _28196_);
  and (_03210_, _28199_, _28192_);
  not (_28200_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_28201_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_28202_, _28201_, _28200_);
  or (_28203_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_28204_, _28203_, _25964_);
  and (_03212_, _28204_, _28202_);
  and (_03215_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _25964_);
  not (_28205_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_28206_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_28207_, _28206_, _28205_);
  and (_28208_, _28206_, _28205_);
  nor (_28209_, _28208_, _28207_);
  not (_28210_, _28209_);
  and (_28211_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_28212_, _28211_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_28213_, _28211_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_28214_, _28213_, _28212_);
  or (_28215_, _28214_, _28206_);
  and (_28216_, _28215_, _28210_);
  nor (_28217_, _28207_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_28218_, _28207_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_28219_, _28218_, _28217_);
  or (_28220_, _28212_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_03221_, _28220_, _25964_);
  and (_28221_, _03221_, _28219_);
  and (_03218_, _28221_, _28216_);
  not (_28222_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_28223_, _27592_, _28222_);
  and (_28224_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_28225_, _28223_);
  and (_28226_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_28227_, _28226_, _28224_);
  and (_03224_, _28227_, _25964_);
  and (_28228_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_28229_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_28230_, _28229_, _28228_);
  and (_03226_, _28230_, _25964_);
  and (_28231_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_28232_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_28233_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _28232_);
  and (_28234_, _28233_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_28235_, _28234_, _28231_);
  and (_03228_, _28235_, _25964_);
  and (_28236_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_28237_, _28236_, _28233_);
  and (_03230_, _28237_, _25964_);
  or (_28238_, _28232_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_03232_, _28238_, _25964_);
  not (_28239_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_28240_, _28239_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_28241_, _28240_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_28242_, _28232_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_28243_, _28242_, _25964_);
  and (_03234_, _28243_, _28241_);
  or (_28244_, _28232_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_03236_, _28244_, _25964_);
  nor (_28245_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_28246_, _28245_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_28247_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_28248_, _28247_, _28246_);
  and (_03238_, _28248_, _25964_);
  and (_28249_, _28222_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_28250_, _28249_, _28246_);
  and (_03240_, _28250_, _25964_);
  or (_28251_, _28246_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  nand (_28252_, _28246_, _23149_);
  and (_28253_, _28252_, _25964_);
  and (_03242_, _28253_, _28251_);
  nand (_28254_, _21114_, _25964_);
  nor (_03244_, _28254_, _22572_);
  or (_28255_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nand (_28256_, _26505_, _27473_);
  and (_28257_, _28256_, _25964_);
  and (_03626_, _28257_, _28255_);
  or (_28258_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_28259_, _26505_, _27466_);
  and (_28260_, _28259_, _25964_);
  and (_03628_, _28260_, _28258_);
  or (_28261_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_28262_, _26505_, _27460_);
  and (_28263_, _28262_, _25964_);
  and (_03630_, _28263_, _28261_);
  or (_28264_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_28265_, _26505_, _27452_);
  and (_28266_, _28265_, _25964_);
  and (_03632_, _28266_, _28264_);
  or (_28267_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_28268_, _26505_, _27446_);
  and (_28269_, _28268_, _25964_);
  and (_03634_, _28269_, _28267_);
  or (_28270_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_28271_, _26505_, _27438_);
  and (_28272_, _28271_, _25964_);
  and (_03636_, _28272_, _28270_);
  or (_28273_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_28274_, _26505_, _27428_);
  and (_28275_, _28274_, _25964_);
  and (_03638_, _28275_, _28273_);
  or (_28276_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand (_28277_, _26505_, _27425_);
  and (_28278_, _28277_, _25964_);
  and (_03640_, _28278_, _28276_);
  or (_28279_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  not (_28280_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nand (_28281_, _26505_, _28280_);
  and (_28282_, _28281_, _25964_);
  and (_03642_, _28282_, _28279_);
  or (_28283_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_28284_, _26505_, _27424_);
  and (_28285_, _28284_, _25964_);
  and (_03644_, _28285_, _28283_);
  or (_28286_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_28287_, _26505_, _27423_);
  and (_28288_, _28287_, _25964_);
  and (_03646_, _28288_, _28286_);
  or (_28289_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_28290_, _26505_, _27422_);
  and (_28291_, _28290_, _25964_);
  and (_03648_, _28291_, _28289_);
  or (_28292_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_28293_, _26505_, _27420_);
  and (_28294_, _28293_, _25964_);
  and (_03650_, _28294_, _28292_);
  or (_28295_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_28296_, _26505_, _27419_);
  and (_28297_, _28296_, _25964_);
  and (_03652_, _28297_, _28295_);
  or (_28298_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_28299_, _26505_, _27417_);
  and (_28300_, _28299_, _25964_);
  and (_03654_, _28300_, _28298_);
  and (_28301_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_28302_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_28303_, _28302_, _28301_);
  and (_03686_, _28303_, _25964_);
  and (_28304_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_28305_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_28306_, _28305_, _28304_);
  and (_03688_, _28306_, _25964_);
  and (_28307_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_28308_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_28309_, _28308_, _28307_);
  and (_03690_, _28309_, _25964_);
  and (_28310_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_28311_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_28312_, _28311_, _28310_);
  and (_03692_, _28312_, _25964_);
  and (_28313_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_28314_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_28315_, _28314_, _28313_);
  and (_03694_, _28315_, _25964_);
  and (_28316_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_28317_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or (_28318_, _28317_, _28316_);
  and (_03696_, _28318_, _25964_);
  and (_28319_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_28320_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or (_28321_, _28320_, _28319_);
  and (_03698_, _28321_, _25964_);
  and (_28322_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_28323_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_28324_, _28323_, _28322_);
  and (_03700_, _28324_, _25964_);
  and (_28325_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_28326_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  or (_28327_, _28326_, _28325_);
  and (_03702_, _28327_, _25964_);
  and (_28328_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and (_28329_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  or (_28330_, _28329_, _28328_);
  and (_03704_, _28330_, _25964_);
  and (_28331_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_28333_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or (_28334_, _28333_, _28331_);
  and (_03706_, _28334_, _25964_);
  and (_28335_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_28336_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  or (_28337_, _28336_, _28335_);
  and (_03708_, _28337_, _25964_);
  and (_28338_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_28339_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or (_28340_, _28339_, _28338_);
  and (_03710_, _28340_, _25964_);
  and (_28342_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_28343_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_28344_, _28343_, _28342_);
  and (_03712_, _28344_, _25964_);
  and (_28345_, _26506_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and (_28346_, _26505_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_28347_, _28346_, _28345_);
  and (_03714_, _28347_, _25964_);
  and (_28348_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_28350_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_28351_, _28350_, _28223_);
  or (_28352_, _28351_, _28348_);
  and (_05586_, _28352_, _25964_);
  and (_28353_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_28354_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_28355_, _28354_, _28353_);
  and (_05588_, _28355_, _25964_);
  and (_28356_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_28357_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_28359_, _28357_, _28223_);
  or (_28360_, _28359_, _28356_);
  and (_05590_, _28360_, _25964_);
  and (_28361_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_28362_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or (_28363_, _28362_, _28361_);
  and (_05592_, _28363_, _25964_);
  and (_28364_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_28365_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_28366_, _28365_, _28223_);
  or (_28368_, _28366_, _28364_);
  and (_05594_, _28368_, _25964_);
  and (_28369_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_28370_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_28371_, _28370_, _28223_);
  or (_28372_, _28371_, _28369_);
  and (_05596_, _28372_, _25964_);
  and (_28373_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_28374_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_28375_, _28374_, _28223_);
  or (_28377_, _28375_, _28373_);
  and (_05598_, _28377_, _25964_);
  and (_28378_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_28379_, _28223_, _28201_);
  or (_28380_, _28379_, _28378_);
  and (_05600_, _28380_, _25964_);
  and (_28381_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_28382_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_28383_, _28382_, _28381_);
  and (_05602_, _28383_, _25964_);
  and (_28385_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_28386_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_28387_, _28386_, _28385_);
  and (_05604_, _28387_, _25964_);
  and (_28388_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_28389_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_28390_, _28389_, _28388_);
  and (_05606_, _28390_, _25964_);
  and (_28391_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_28392_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_28394_, _28392_, _28391_);
  and (_05608_, _28394_, _25964_);
  and (_28395_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_28396_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_28397_, _28396_, _28395_);
  and (_05610_, _28397_, _25964_);
  and (_28398_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_28399_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_28400_, _28399_, _28398_);
  and (_05612_, _28400_, _25964_);
  and (_28402_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_28403_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_28404_, _28403_, _28402_);
  and (_05614_, _28404_, _25964_);
  and (_28405_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_28406_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_28407_, _28406_, _28405_);
  and (_05616_, _28407_, _25964_);
  and (_28408_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_28409_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_28411_, _28409_, _28408_);
  and (_05618_, _28411_, _25964_);
  and (_28412_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_28413_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_28414_, _28413_, _28412_);
  and (_05620_, _28414_, _25964_);
  and (_28415_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_28416_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_28417_, _28416_, _28415_);
  and (_05622_, _28417_, _25964_);
  and (_28419_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_28420_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_28421_, _28420_, _28419_);
  and (_05624_, _28421_, _25964_);
  and (_28422_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_28423_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_28424_, _28423_, _28422_);
  and (_05626_, _28424_, _25964_);
  and (_28425_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_28426_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_28428_, _28426_, _28425_);
  and (_05628_, _28428_, _25964_);
  and (_28429_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_28430_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_28431_, _28430_, _28429_);
  and (_05630_, _28431_, _25964_);
  and (_28432_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_28433_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_28434_, _28433_, _28432_);
  and (_05632_, _28434_, _25964_);
  and (_28436_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_28437_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_28438_, _28437_, _28436_);
  and (_05634_, _28438_, _25964_);
  and (_28439_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_28440_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_28441_, _28440_, _28439_);
  and (_05636_, _28441_, _25964_);
  and (_28442_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_28443_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_28445_, _28443_, _28442_);
  and (_05638_, _28445_, _25964_);
  and (_28446_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_28447_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_28448_, _28447_, _28446_);
  and (_05640_, _28448_, _25964_);
  and (_28449_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_28450_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_28451_, _28450_, _28449_);
  and (_05642_, _28451_, _25964_);
  and (_28452_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_28453_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_28454_, _28453_, _28452_);
  and (_05644_, _28454_, _25964_);
  and (_28455_, _28223_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_28456_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_28457_, _28456_, _28455_);
  and (_05646_, _28457_, _25964_);
  and (_05649_, _19984_, _25964_);
  and (_05652_, _20236_, _25964_);
  and (_05655_, _20467_, _25964_);
  nor (_05657_, _24350_, rst);
  nor (_05660_, _24539_, rst);
  nor (_05663_, _24659_, rst);
  nor (_05666_, _24458_, rst);
  nor (_05669_, _24507_, rst);
  nor (_05672_, _24612_, rst);
  nor (_05675_, _24403_, rst);
  nor (_05678_, _24567_, rst);
  and (_05708_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _25964_);
  and (_05710_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _25964_);
  and (_05712_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _25964_);
  and (_05714_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _25964_);
  and (_05716_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _25964_);
  and (_05718_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _25964_);
  and (_05720_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _25964_);
  or (_28458_, _27407_, _27383_);
  and (_28459_, _28458_, ABINPUT[19]);
  not (_28460_, _27393_);
  nor (_28461_, _28460_, _26261_);
  and (_28462_, _27562_, _24528_);
  or (_28463_, _28462_, _28461_);
  and (_28464_, _27392_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_28465_, _28464_, _28463_);
  nand (_28466_, _27477_, _27473_);
  not (_28467_, _27557_);
  nor (_28468_, _28467_, _27478_);
  and (_28469_, _28468_, _28466_);
  or (_28470_, _28469_, _28465_);
  nor (_28471_, _28470_, _28459_);
  nand (_28472_, _28471_, _27380_);
  or (_28473_, _27380_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_28474_, _28473_, _25964_);
  and (_05722_, _28474_, _28472_);
  and (_28475_, _28458_, ABINPUT[20]);
  nor (_28476_, _28460_, _26278_);
  and (_28477_, _27467_, _27363_);
  and (_28478_, _22134_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_28479_, _28478_, _28477_);
  or (_28480_, _28479_, _28476_);
  or (_28481_, _28480_, _28475_);
  nor (_28482_, _27481_, _27478_);
  nor (_28483_, _28482_, _27482_);
  and (_28484_, _28483_, _27557_);
  nor (_28485_, _28484_, _28481_);
  nand (_28486_, _28485_, _27380_);
  or (_28487_, _27380_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_28488_, _28487_, _25964_);
  and (_05724_, _28488_, _28486_);
  and (_28489_, _28458_, ABINPUT[21]);
  nor (_28490_, _28460_, _26295_);
  and (_28491_, _27461_, _27363_);
  and (_28492_, _22134_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_28493_, _28492_, _28491_);
  or (_28494_, _28493_, _28490_);
  or (_28495_, _28494_, _28489_);
  nor (_28496_, _27487_, _27485_);
  nor (_28497_, _28496_, _27489_);
  and (_28498_, _28497_, _27557_);
  or (_28499_, _28498_, _28495_);
  and (_28500_, _28499_, _27380_);
  not (_28501_, _27380_);
  not (_28502_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_28503_, _27592_, _28502_);
  and (_28504_, _27592_, _28502_);
  nor (_28505_, _28504_, _28503_);
  and (_28506_, _28505_, _28501_);
  or (_28507_, _28506_, _28500_);
  and (_05726_, _28507_, _25964_);
  and (_28508_, _28458_, ABINPUT[22]);
  nor (_28509_, _28460_, _26312_);
  and (_28510_, _27454_, _27363_);
  and (_28511_, _22134_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_28512_, _28511_, _28510_);
  or (_28513_, _28512_, _28509_);
  or (_28514_, _28513_, _28508_);
  or (_28515_, _27459_, _27458_);
  or (_28516_, _28515_, _27490_);
  nand (_28517_, _28515_, _27490_);
  and (_28518_, _28517_, _28516_);
  and (_28519_, _28518_, _27557_);
  or (_28520_, _28519_, _28514_);
  and (_28521_, _28520_, _27380_);
  and (_28522_, _28503_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_28523_, _28503_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_28524_, _28523_, _28522_);
  and (_28525_, _28524_, _28501_);
  or (_28526_, _28525_, _28521_);
  and (_05728_, _28526_, _25964_);
  and (_28527_, _28458_, ABINPUT[23]);
  nor (_28528_, _28460_, _26329_);
  and (_28529_, _27447_, _27363_);
  and (_28530_, _22134_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_28531_, _28530_, _28529_);
  or (_28532_, _28531_, _28528_);
  or (_28533_, _28532_, _28527_);
  or (_28534_, _27495_, _27493_);
  and (_28535_, _28534_, _27496_);
  and (_28536_, _28535_, _27557_);
  or (_28537_, _28536_, _28533_);
  and (_28538_, _28537_, _27380_);
  and (_28539_, _28503_, _27594_);
  nor (_28540_, _28522_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_28541_, _28540_, _28539_);
  nor (_28542_, _28541_, _27380_);
  or (_28543_, _28542_, _28538_);
  and (_05730_, _28543_, _25964_);
  and (_28544_, _28458_, ABINPUT[24]);
  nor (_28545_, _28460_, _26346_);
  and (_28546_, _27439_, _27363_);
  and (_28547_, _22134_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_28548_, _28547_, _28546_);
  or (_28549_, _28548_, _28545_);
  or (_28550_, _28549_, _28544_);
  or (_28551_, _27444_, _27443_);
  nand (_28552_, _28551_, _27498_);
  or (_28553_, _28551_, _27498_);
  and (_28554_, _28553_, _28552_);
  and (_28555_, _28554_, _27557_);
  or (_28556_, _28555_, _28550_);
  and (_28557_, _28556_, _27380_);
  and (_28558_, _28539_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_28559_, _28539_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_28560_, _28559_, _28558_);
  nor (_28561_, _28560_, _27380_);
  or (_28562_, _28561_, _28557_);
  and (_05732_, _28562_, _25964_);
  and (_28563_, _28458_, ABINPUT[25]);
  nor (_28564_, _28460_, _26363_);
  and (_28565_, _27430_, _27363_);
  and (_28566_, _22134_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_28567_, _28566_, _28565_);
  or (_28568_, _28567_, _28564_);
  or (_28569_, _28568_, _28563_);
  nor (_28570_, _27500_, _27436_);
  nor (_28571_, _28570_, _27502_);
  and (_28572_, _28571_, _27557_);
  or (_28573_, _28572_, _28569_);
  and (_28574_, _28573_, _27380_);
  and (_28575_, _28558_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_28576_, _28558_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_28577_, _28576_, _28575_);
  nor (_28578_, _28577_, _27380_);
  or (_28579_, _28578_, _28574_);
  and (_05734_, _28579_, _25964_);
  and (_28580_, _28458_, ABINPUT[26]);
  nor (_28581_, _28460_, _26244_);
  and (_28582_, _27414_, _27363_);
  and (_28583_, _22134_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_28584_, _28583_, _28582_);
  or (_28585_, _28584_, _28581_);
  or (_28586_, _28585_, _28580_);
  or (_28587_, _27426_, _27427_);
  nand (_28588_, _28587_, _27503_);
  or (_28589_, _28587_, _27503_);
  and (_28590_, _28589_, _28588_);
  and (_28591_, _28590_, _27557_);
  or (_28592_, _28591_, _28586_);
  and (_28593_, _28592_, _27380_);
  nor (_28594_, _28575_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_28595_, _28594_, _27601_);
  nor (_28596_, _28595_, _27380_);
  or (_28597_, _28596_, _28593_);
  and (_05736_, _28597_, _25964_);
  and (_28598_, _27506_, _28280_);
  nor (_28599_, _27506_, _28280_);
  nor (_28600_, _28599_, _28598_);
  or (_28601_, _28600_, _27416_);
  nor (_28602_, _27404_, _27535_);
  nand (_28603_, _28600_, _27416_);
  and (_28604_, _28603_, _28602_);
  and (_28605_, _28604_, _28601_);
  and (_28606_, _27407_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_28607_, _27383_, ABINPUT[11]);
  and (_28608_, _22134_, ABINPUT[19]);
  or (_28609_, _28608_, _28607_);
  nor (_28610_, _28609_, _28606_);
  and (_28611_, _27393_, _24528_);
  and (_28612_, _27562_, _27813_);
  nor (_28613_, _28612_, _28611_);
  and (_28614_, _28613_, _28610_);
  nand (_28615_, _28614_, _27380_);
  or (_28616_, _28615_, _28605_);
  nor (_28617_, _27601_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_28618_, _28617_, _27602_);
  or (_28619_, _28618_, _27380_);
  and (_28620_, _28619_, _25964_);
  and (_05738_, _28620_, _28616_);
  and (_28621_, _27506_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_28622_, _28621_, _27416_);
  and (_28623_, _27507_, _27518_);
  nor (_28624_, _28623_, _28622_);
  nand (_28625_, _28624_, _27424_);
  or (_28626_, _28624_, _27424_);
  and (_28627_, _28626_, _28602_);
  and (_28628_, _28627_, _28625_);
  and (_28629_, _27407_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_28630_, _27383_, ABINPUT[12]);
  and (_28631_, _22134_, ABINPUT[20]);
  or (_28632_, _28631_, _28630_);
  nor (_28633_, _28632_, _28629_);
  and (_28634_, _27393_, _24676_);
  and (_28635_, _27562_, _27731_);
  nor (_28636_, _28635_, _28634_);
  and (_28637_, _28636_, _28633_);
  nand (_28638_, _28637_, _27380_);
  or (_28639_, _28638_, _28628_);
  and (_28640_, _27599_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_28641_, _28640_, _27593_);
  nor (_28642_, _28641_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_28643_, _28641_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_28644_, _28643_, _28642_);
  or (_28645_, _28644_, _27380_);
  and (_28646_, _28645_, _25964_);
  and (_05740_, _28646_, _28639_);
  and (_28647_, _27508_, _27518_);
  and (_28648_, _28622_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_28649_, _28648_, _28647_);
  nand (_28650_, _28649_, _27423_);
  or (_28651_, _28649_, _27423_);
  and (_28652_, _28651_, _28602_);
  and (_28653_, _28652_, _28650_);
  and (_28654_, _27407_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_28655_, _27383_, ABINPUT[13]);
  and (_28656_, _22134_, ABINPUT[21]);
  or (_28657_, _28656_, _28655_);
  nor (_28658_, _28657_, _28654_);
  and (_28659_, _27393_, _24447_);
  and (_28660_, _27562_, _27840_);
  nor (_28661_, _28660_, _28659_);
  and (_28662_, _28661_, _28658_);
  nand (_28663_, _28662_, _27380_);
  or (_28664_, _28663_, _28653_);
  nor (_28665_, _28643_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_28666_, _28643_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_28667_, _28666_, _28665_);
  or (_28668_, _28667_, _27380_);
  and (_28669_, _28668_, _25964_);
  and (_05742_, _28669_, _28664_);
  and (_28670_, _27522_, _27416_);
  and (_28671_, _27510_, _27518_);
  nor (_28672_, _28671_, _28670_);
  nand (_28673_, _28672_, _27422_);
  or (_28674_, _28672_, _27422_);
  and (_28675_, _28674_, _28602_);
  and (_28676_, _28675_, _28673_);
  nor (_28677_, _27571_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_28678_, _28677_, _27573_);
  and (_28679_, _28678_, _27562_);
  and (_28680_, _27383_, ABINPUT[14]);
  and (_28681_, _22134_, ABINPUT[22]);
  or (_28682_, _28681_, _28680_);
  nor (_28683_, _28682_, _28679_);
  and (_28684_, _27393_, _24492_);
  and (_28685_, _27407_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_28686_, _28685_, _28684_);
  and (_28687_, _28686_, _28683_);
  nand (_28688_, _28687_, _27380_);
  or (_28689_, _28688_, _28676_);
  nor (_28690_, _28666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_28691_, _28690_, _27605_);
  or (_28692_, _28691_, _27380_);
  and (_28693_, _28692_, _25964_);
  and (_05744_, _28693_, _28689_);
  nand (_28694_, _27383_, ABINPUT[15]);
  nand (_28695_, _27393_, _24634_);
  nand (_28696_, _27392_, ABINPUT[23]);
  and (_28697_, _28696_, _28695_);
  and (_28698_, _28697_, _28694_);
  nor (_28699_, _27573_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_28700_, _28699_, _27574_);
  and (_28701_, _28700_, _27562_);
  and (_28702_, _27407_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_28703_, _28702_, _28701_);
  and (_28704_, _27523_, _27416_);
  and (_28705_, _27511_, _27518_);
  nor (_28706_, _28705_, _28704_);
  and (_28707_, _28706_, _27420_);
  nor (_28708_, _28706_, _27420_);
  or (_28709_, _28708_, _28707_);
  or (_28710_, _28709_, _28467_);
  and (_28711_, _28710_, _28703_);
  and (_28712_, _28711_, _28698_);
  nand (_28713_, _28712_, _27380_);
  nor (_28714_, _27605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_28715_, _28714_, _27606_);
  or (_28716_, _28715_, _27380_);
  and (_28717_, _28716_, _25964_);
  and (_05746_, _28717_, _28713_);
  and (_28718_, _27407_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_28719_, _27393_, _24421_);
  and (_28720_, _27392_, ABINPUT[24]);
  or (_28721_, _28720_, _28719_);
  or (_28722_, _28721_, _28718_);
  and (_28723_, _27525_, _27416_);
  and (_28724_, _27512_, _27518_);
  nor (_28725_, _28724_, _28723_);
  nor (_28726_, _28725_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_28727_, _28725_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_28728_, _28727_, _28726_);
  and (_28729_, _28728_, _27557_);
  or (_28730_, _28729_, _28722_);
  and (_28731_, _27383_, ABINPUT[16]);
  nor (_28732_, _27574_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_28733_, _28732_, _27575_);
  and (_28734_, _28733_, _27562_);
  nor (_28735_, _28734_, _28731_);
  nand (_28736_, _28735_, _27380_);
  or (_28737_, _28736_, _28730_);
  nor (_28738_, _27606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_28739_, _28738_, _27607_);
  or (_28740_, _28739_, _27380_);
  and (_28741_, _28740_, _25964_);
  and (_05748_, _28741_, _28737_);
  nor (_28742_, _27416_, _27419_);
  and (_28743_, _27416_, _27419_);
  nor (_28744_, _28743_, _28742_);
  not (_28745_, _28744_);
  nor (_28746_, _28745_, _28725_);
  nor (_28747_, _28746_, _27417_);
  and (_28748_, _28746_, _27417_);
  or (_28749_, _28748_, _28747_);
  and (_28750_, _28749_, _28602_);
  nor (_28751_, _27575_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_28752_, _28751_, _27577_);
  and (_28753_, _28752_, _27562_);
  and (_28754_, _27383_, ABINPUT[17]);
  and (_28755_, _22134_, ABINPUT[25]);
  or (_28756_, _28755_, _28754_);
  or (_28757_, _28756_, _28753_);
  and (_28758_, _27393_, _24587_);
  and (_28759_, _27407_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_28760_, _28759_, _28758_);
  or (_28761_, _28760_, _28757_);
  or (_28762_, _28761_, _28750_);
  or (_28763_, _28762_, _28501_);
  nor (_28764_, _27607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_28765_, _28764_, _27609_);
  or (_28766_, _28765_, _27380_);
  and (_28767_, _28766_, _25964_);
  and (_05750_, _28767_, _28763_);
  or (_28768_, _28117_, _28115_);
  nor (_28769_, _27623_, _28118_);
  and (_28770_, _28769_, _28768_);
  nor (_28771_, _27621_, _27473_);
  or (_28772_, _28771_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_28773_, _28772_, _28770_);
  or (_28774_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _18488_);
  and (_28775_, _28774_, _25964_);
  and (_05752_, _28775_, _28773_);
  or (_28776_, _28120_, _28118_);
  and (_28777_, _28776_, _28121_);
  or (_28778_, _28777_, _27623_);
  or (_28779_, _27621_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_28780_, _28779_, _28154_);
  and (_28781_, _28780_, _28778_);
  and (_28782_, _27617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_05754_, _28782_, _28781_);
  or (_28783_, _28125_, _28123_);
  nor (_28784_, _27623_, _28126_);
  and (_28785_, _28784_, _28783_);
  nor (_28786_, _27621_, _27460_);
  or (_28787_, _28786_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_28788_, _28787_, _28785_);
  or (_28789_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _18488_);
  and (_28790_, _28789_, _25964_);
  and (_05756_, _28790_, _28788_);
  and (_28791_, _27617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_28792_, _28126_, _27730_);
  nor (_28793_, _28792_, _28127_);
  or (_28794_, _28793_, _27623_);
  or (_28795_, _27621_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_28796_, _28795_, _28154_);
  and (_28797_, _28796_, _28794_);
  or (_05758_, _28797_, _28791_);
  and (_28798_, _27617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_28799_, _28130_, _28127_);
  nor (_28800_, _28799_, _28131_);
  or (_28801_, _28800_, _27623_);
  or (_28802_, _27621_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_28803_, _28802_, _28154_);
  and (_28804_, _28803_, _28801_);
  or (_05760_, _28804_, _28798_);
  or (_28805_, _28131_, _27715_);
  nor (_28806_, _27623_, _28132_);
  and (_28807_, _28806_, _28805_);
  nor (_28808_, _27621_, _27438_);
  or (_28809_, _28808_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_28810_, _28809_, _28807_);
  or (_28811_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _18488_);
  and (_28812_, _28811_, _25964_);
  and (_05762_, _28812_, _28810_);
  and (_28813_, _27617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_28814_, _28132_, _27711_);
  nor (_28815_, _28814_, _28133_);
  or (_28816_, _28815_, _27623_);
  or (_28817_, _27621_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_28818_, _28817_, _28154_);
  and (_28819_, _28818_, _28816_);
  or (_05764_, _28819_, _28813_);
  and (_28820_, _27617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_28821_, _28133_, _27708_);
  nor (_28822_, _28821_, _28134_);
  or (_28823_, _28822_, _27623_);
  or (_28824_, _27621_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_28825_, _28824_, _28154_);
  and (_28826_, _28825_, _28823_);
  or (_05766_, _28826_, _28820_);
  nor (_28827_, _28136_, _28134_);
  nor (_28828_, _28827_, _28137_);
  or (_28829_, _28828_, _27623_);
  or (_28830_, _27621_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_28831_, _28830_, _28154_);
  and (_28832_, _28831_, _28829_);
  and (_28833_, _27617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_05768_, _28833_, _28832_);
  and (_28834_, _27617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_28835_, _28137_, _27701_);
  nor (_28836_, _28835_, _28138_);
  or (_28837_, _28836_, _27623_);
  or (_28838_, _27621_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_28839_, _28838_, _28154_);
  and (_28840_, _28839_, _28837_);
  or (_05770_, _28840_, _28834_);
  or (_28841_, _28138_, _27692_);
  nor (_28842_, _27623_, _28139_);
  and (_28843_, _28842_, _28841_);
  nor (_28844_, _27621_, _27423_);
  or (_28845_, _28844_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_28846_, _28845_, _28843_);
  or (_28847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _18488_);
  and (_28848_, _28847_, _25964_);
  and (_05772_, _28848_, _28846_);
  nor (_28849_, _28139_, _27690_);
  nor (_28850_, _28849_, _28140_);
  or (_28851_, _28850_, _27623_);
  or (_28852_, _27621_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_28853_, _28852_, _28154_);
  and (_28854_, _28853_, _28851_);
  and (_28855_, _27617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_05774_, _28855_, _28854_);
  and (_28856_, _27617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_28857_, _28142_, _28140_);
  nor (_28858_, _28857_, _28143_);
  or (_28859_, _28858_, _27623_);
  or (_28860_, _27621_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_28861_, _28860_, _28154_);
  and (_28862_, _28861_, _28859_);
  or (_05775_, _28862_, _28856_);
  nor (_28863_, _28143_, _27681_);
  nor (_28864_, _28863_, _28144_);
  or (_28865_, _28864_, _27623_);
  or (_28866_, _27621_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_28867_, _28866_, _28154_);
  and (_28868_, _28867_, _28865_);
  and (_28869_, _27617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_05777_, _28869_, _28868_);
  and (_28870_, _27617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_28871_, _28144_, _27676_);
  nor (_28872_, _28871_, _28145_);
  or (_28873_, _28872_, _27623_);
  or (_28874_, _27621_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_28875_, _28874_, _28154_);
  and (_28876_, _28875_, _28873_);
  or (_05779_, _28876_, _28870_);
  and (_28877_, _28164_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_28878_, _28877_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_05781_, _28878_, _25964_);
  and (_28879_, _28164_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_28880_, _28879_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_05783_, _28880_, _25964_);
  and (_28881_, _28164_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_28882_, _28881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_05785_, _28882_, _25964_);
  and (_28883_, _28164_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_28884_, _28883_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_05787_, _28884_, _25964_);
  and (_28885_, _28164_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_28886_, _28885_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_05789_, _28886_, _25964_);
  and (_28887_, _28164_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_28888_, _28887_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_05791_, _28888_, _25964_);
  and (_28889_, _28164_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_28890_, _28889_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_05793_, _28890_, _25964_);
  nor (_28891_, _28114_, _24319_);
  nand (_28892_, _28891_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_28893_, _28891_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_28894_, _28893_, _28154_);
  and (_05795_, _28894_, _28892_);
  or (_28895_, _28175_, _28173_);
  and (_28896_, _28895_, _28176_);
  or (_28897_, _28896_, _24319_);
  or (_28898_, _18521_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_28899_, _28898_, _28154_);
  and (_05797_, _28899_, _28897_);
  or (_28900_, _28350_, _28200_);
  or (_28901_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_28902_, _28901_, _25964_);
  and (_05827_, _28902_, _28900_);
  and (_28903_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  or (_28904_, _28903_, _28200_);
  or (_28905_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_28906_, _28905_, _25964_);
  and (_05829_, _28906_, _28904_);
  or (_28907_, _28357_, _28200_);
  or (_28908_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_28909_, _28908_, _25964_);
  and (_05831_, _28909_, _28907_);
  and (_28910_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_28911_, _28910_, _28200_);
  or (_28912_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_28913_, _28912_, _25964_);
  and (_05833_, _28913_, _28911_);
  or (_28914_, _28365_, _28200_);
  or (_28915_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_28916_, _28915_, _25964_);
  and (_05835_, _28916_, _28914_);
  or (_28917_, _28370_, _28200_);
  or (_28918_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_28919_, _28918_, _25964_);
  and (_05837_, _28919_, _28917_);
  or (_28920_, _28374_, _28200_);
  or (_28921_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_28922_, _28921_, _25964_);
  and (_05839_, _28922_, _28920_);
  and (_05841_, _28209_, _25964_);
  nor (_05843_, _28219_, rst);
  and (_05845_, _28215_, _25964_);
  and (_28923_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_28924_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_28925_, _28924_, _28923_);
  and (_05847_, _28925_, _25964_);
  and (_28926_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_28927_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_28928_, _28927_, _28926_);
  and (_05849_, _28928_, _25964_);
  and (_28929_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_28930_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_28931_, _28930_, _28929_);
  and (_05851_, _28931_, _25964_);
  and (_28932_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_28933_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_28934_, _28933_, _28932_);
  and (_05853_, _28934_, _25964_);
  and (_28935_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_28936_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_28937_, _28936_, _28935_);
  and (_05855_, _28937_, _25964_);
  and (_28938_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_28939_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_28940_, _28939_, _28938_);
  and (_05857_, _28940_, _25964_);
  and (_28941_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_28942_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_28943_, _28942_, _28941_);
  and (_05859_, _28943_, _25964_);
  and (_28944_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_28945_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_28946_, _28945_, _28944_);
  and (_05861_, _28946_, _25964_);
  and (_28947_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_28948_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_28949_, _28948_, _28947_);
  and (_05863_, _28949_, _25964_);
  and (_28950_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_28951_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_28952_, _28951_, _28950_);
  and (_05865_, _28952_, _25964_);
  and (_28953_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_28954_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_28955_, _28954_, _28953_);
  and (_05867_, _28955_, _25964_);
  and (_28956_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_28957_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_28958_, _28957_, _28956_);
  and (_05869_, _28958_, _25964_);
  and (_28959_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_28960_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_28961_, _28960_, _28959_);
  and (_05871_, _28961_, _25964_);
  and (_28962_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_28963_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_28964_, _28963_, _28962_);
  and (_05873_, _28964_, _25964_);
  and (_28965_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_28966_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_28967_, _28966_, _28965_);
  and (_05875_, _28967_, _25964_);
  and (_28968_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_28969_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_28970_, _28969_, _28968_);
  and (_05877_, _28970_, _25964_);
  and (_28971_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_28972_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_28973_, _28972_, _28971_);
  and (_05879_, _28973_, _25964_);
  and (_28974_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_28975_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_28976_, _28975_, _28974_);
  and (_05881_, _28976_, _25964_);
  and (_28977_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_28978_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_28979_, _28978_, _28977_);
  and (_05883_, _28979_, _25964_);
  and (_28980_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_28981_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_28982_, _28981_, _28980_);
  and (_05885_, _28982_, _25964_);
  and (_28983_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_28984_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_28985_, _28984_, _28983_);
  and (_05887_, _28985_, _25964_);
  and (_28986_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_28987_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_28988_, _28987_, _28986_);
  and (_05889_, _28988_, _25964_);
  and (_28989_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_28990_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_28991_, _28990_, _28989_);
  and (_05891_, _28991_, _25964_);
  and (_28992_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_28993_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_28994_, _28993_, _28992_);
  and (_05893_, _28994_, _25964_);
  and (_28995_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_28996_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_28997_, _28996_, _28995_);
  and (_05895_, _28997_, _25964_);
  and (_28998_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_28999_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_29000_, _28999_, _28998_);
  and (_05897_, _29000_, _25964_);
  and (_29001_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_29002_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_29003_, _29002_, _29001_);
  and (_05899_, _29003_, _25964_);
  and (_29004_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_29005_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_29006_, _29005_, _29004_);
  and (_05901_, _29006_, _25964_);
  and (_29007_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_29008_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_29009_, _29008_, _29007_);
  and (_05903_, _29009_, _25964_);
  and (_29010_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_29011_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_29012_, _29011_, _29010_);
  and (_05905_, _29012_, _25964_);
  and (_29013_, _28223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_29014_, _28225_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_29015_, _29014_, _29013_);
  and (_05907_, _29015_, _25964_);
  and (_29016_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_29017_, _28233_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_29018_, _29017_, _29016_);
  and (_05909_, _29018_, _25964_);
  and (_29019_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_29020_, _28233_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_29021_, _29020_, _29019_);
  and (_05911_, _29021_, _25964_);
  and (_29022_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_29023_, _28233_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_29024_, _29023_, _29022_);
  and (_05913_, _29024_, _25964_);
  and (_29025_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_29026_, _28233_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_29027_, _29026_, _29025_);
  and (_05915_, _29027_, _25964_);
  and (_29028_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_29029_, _28233_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_29030_, _29029_, _29028_);
  and (_05917_, _29030_, _25964_);
  and (_29031_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_29032_, _28233_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_29033_, _29032_, _29031_);
  and (_05919_, _29033_, _25964_);
  and (_29034_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_29035_, _28233_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_29036_, _29035_, _29034_);
  and (_05921_, _29036_, _25964_);
  and (_29037_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_29038_, _24539_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_29039_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_29040_, _29039_, _28232_);
  and (_29041_, _29040_, _29038_);
  or (_29042_, _29041_, _29037_);
  and (_05923_, _29042_, _25964_);
  and (_29043_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_29044_, _24659_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_29045_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_29046_, _29045_, _28232_);
  and (_29047_, _29046_, _29044_);
  or (_29048_, _29047_, _29043_);
  and (_05925_, _29048_, _25964_);
  and (_29049_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_29050_, _24458_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_29051_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_29052_, _29051_, _28232_);
  and (_29053_, _29052_, _29050_);
  or (_29054_, _29053_, _29049_);
  and (_05927_, _29054_, _25964_);
  and (_29055_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_29056_, _24507_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_29057_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_29058_, _29057_, _28232_);
  and (_29059_, _29058_, _29056_);
  or (_29060_, _29059_, _29055_);
  and (_05929_, _29060_, _25964_);
  and (_29061_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_29062_, _24612_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_29063_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_29064_, _29063_, _28232_);
  and (_29065_, _29064_, _29062_);
  or (_29066_, _29065_, _29061_);
  and (_05931_, _29066_, _25964_);
  and (_29067_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_29068_, _24403_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_29069_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_29070_, _29069_, _28232_);
  and (_29071_, _29070_, _29068_);
  or (_29072_, _29071_, _29067_);
  and (_05933_, _29072_, _25964_);
  and (_29073_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_29074_, _24567_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_29075_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_29076_, _29075_, _28232_);
  and (_29077_, _29076_, _29074_);
  or (_29078_, _29077_, _29073_);
  and (_05935_, _29078_, _25964_);
  and (_29079_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_29080_, _24368_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_29081_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_29082_, _29081_, _28232_);
  and (_29083_, _29082_, _29080_);
  or (_29084_, _29083_, _29079_);
  and (_05937_, _29084_, _25964_);
  and (_29085_, _28239_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_29086_, _29085_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_29087_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _28232_);
  and (_29088_, _29087_, _25964_);
  and (_05938_, _29088_, _29086_);
  and (_29089_, _28239_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_29090_, _29089_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_29091_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _28232_);
  and (_29092_, _29091_, _25964_);
  and (_05940_, _29092_, _29090_);
  and (_29093_, _28239_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_29094_, _29093_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_29095_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _28232_);
  and (_29096_, _29095_, _25964_);
  and (_05942_, _29096_, _29094_);
  and (_29097_, _28239_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_29098_, _29097_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_29099_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _28232_);
  and (_29100_, _29099_, _25964_);
  and (_05944_, _29100_, _29098_);
  and (_29101_, _28239_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_29102_, _29101_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_29103_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _28232_);
  and (_29104_, _29103_, _25964_);
  and (_05946_, _29104_, _29102_);
  and (_29105_, _28239_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_29106_, _29105_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_29107_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _28232_);
  and (_29108_, _29107_, _25964_);
  and (_05948_, _29108_, _29106_);
  and (_29109_, _28239_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_29110_, _29109_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_29111_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _28232_);
  and (_29112_, _29111_, _25964_);
  and (_05950_, _29112_, _29110_);
  not (_29113_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor (_29114_, _28246_, _29113_);
  and (_29115_, _28246_, ABINPUT[19]);
  or (_29116_, _29115_, _29114_);
  and (_05952_, _29116_, _25964_);
  not (_29117_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nor (_29118_, _28246_, _29117_);
  and (_29119_, _28246_, ABINPUT[20]);
  or (_29120_, _29119_, _29118_);
  and (_05954_, _29120_, _25964_);
  not (_29121_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor (_29122_, _28246_, _29121_);
  and (_29123_, _28246_, ABINPUT[21]);
  or (_29124_, _29123_, _29122_);
  and (_05956_, _29124_, _25964_);
  not (_29125_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nor (_29126_, _28246_, _29125_);
  and (_29127_, _28246_, ABINPUT[22]);
  or (_29128_, _29127_, _29126_);
  and (_05958_, _29128_, _25964_);
  or (_29129_, _28246_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  nand (_29130_, _28246_, _18019_);
  and (_29131_, _29130_, _25964_);
  and (_05960_, _29131_, _29129_);
  or (_29132_, _28246_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  nand (_29133_, _28246_, _18194_);
  and (_29134_, _29133_, _25964_);
  and (_05962_, _29134_, _29132_);
  or (_29135_, _28246_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  nand (_29136_, _28246_, _18368_);
  and (_29137_, _29136_, _25964_);
  and (_05964_, _29137_, _29135_);
  or (_29138_, _28246_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  nand (_29139_, _28246_, _17086_);
  and (_29140_, _29139_, _25964_);
  and (_05966_, _29140_, _29138_);
  or (_29141_, _28246_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  nand (_29142_, _28246_, _23166_);
  and (_29143_, _29142_, _25964_);
  and (_05968_, _29143_, _29141_);
  or (_29144_, _28246_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  nand (_29145_, _28246_, _23173_);
  and (_29146_, _29145_, _25964_);
  and (_05970_, _29146_, _29144_);
  or (_29147_, _28246_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  nand (_29148_, _28246_, _23180_);
  and (_29149_, _29148_, _25964_);
  and (_05972_, _29149_, _29147_);
  or (_29150_, _28246_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  nand (_29151_, _28246_, _23187_);
  and (_29152_, _29151_, _25964_);
  and (_05974_, _29152_, _29150_);
  or (_29153_, _28246_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  nand (_29154_, _28246_, _23194_);
  and (_29155_, _29154_, _25964_);
  and (_05976_, _29155_, _29153_);
  or (_29156_, _28246_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  nand (_29157_, _28246_, _23201_);
  and (_29158_, _29157_, _25964_);
  and (_05978_, _29158_, _29156_);
  or (_29159_, _28246_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  nand (_29160_, _28246_, _23208_);
  and (_29161_, _29160_, _25964_);
  and (_05980_, _29161_, _29159_);
  and (_08290_, _24695_, _25964_);
  and (_08293_, _24773_, _25964_);
  nor (_08298_, _24467_, rst);
  and (_08451_, _24795_, _25964_);
  and (_08453_, _24811_, _25964_);
  and (_08455_, _24826_, _25964_);
  and (_08457_, _24841_, _25964_);
  and (_08459_, _24855_, _25964_);
  and (_08461_, _24869_, _25964_);
  and (_08463_, _24883_, _25964_);
  nor (_08465_, _24547_, rst);
  nor (_08467_, _24680_, rst);
  nor (_12124_, _21092_, rst);
  nand (_29162_, _28193_, _22430_);
  nor (_29163_, _20949_, _20730_);
  or (_12127_, _29163_, _29162_);
  and (_29164_, _27814_, _27746_);
  and (_29165_, _29164_, _27933_);
  and (_29166_, _27846_, _19699_);
  and (_29167_, _29166_, _27982_);
  or (_29168_, _29167_, _29165_);
  and (_29169_, _28027_, _27987_);
  and (_29170_, _28027_, _27767_);
  or (_29171_, _29170_, _28109_);
  nor (_29172_, _29171_, _29169_);
  nand (_29173_, _29172_, _28038_);
  or (_29174_, _29173_, _29168_);
  and (_29175_, _27860_, _27982_);
  or (_29176_, _29175_, _28039_);
  and (_29177_, _28054_, _27885_);
  and (_29178_, _28076_, _27933_);
  or (_29179_, _29178_, _29177_);
  or (_29180_, _29179_, _29176_);
  and (_29181_, _27992_, _27785_);
  nor (_29182_, _28087_, _29181_);
  nand (_29183_, _29182_, _28094_);
  nor (_29184_, _28060_, _28051_);
  nand (_29185_, _29184_, _28079_);
  or (_29186_, _29185_, _29183_);
  or (_29187_, _29186_, _29180_);
  or (_29188_, _29187_, _29174_);
  and (_29189_, _29188_, _18532_);
  not (_29190_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_29191_, _18510_, _15520_);
  and (_29192_, _29191_, _20894_);
  nor (_29193_, _29192_, _29190_);
  or (_29194_, _29193_, rst);
  or (_12130_, _29194_, _29189_);
  nand (_29195_, _19135_, _18466_);
  or (_29196_, _18466_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_29197_, _29196_, _25964_);
  and (_12133_, _29197_, _29195_);
  and (_29198_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _25964_);
  and (_29199_, _29198_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_29200_, _20741_, _21322_);
  or (_29201_, _29200_, _21333_);
  nor (_29202_, _29201_, _21914_);
  nand (_29203_, _29202_, _27547_);
  and (_29204_, _21026_, _21969_);
  and (_29205_, _20741_, _20993_);
  or (_29206_, _29205_, _29204_);
  and (_29207_, _20741_, _21629_);
  or (_29208_, _29207_, _27338_);
  or (_29209_, _29208_, _20960_);
  or (_29210_, _29209_, _29206_);
  or (_29211_, _29210_, _29203_);
  and (_29212_, _29211_, _28193_);
  or (_12136_, _29212_, _29199_);
  and (_29213_, _20949_, _20796_);
  or (_29214_, _29213_, _20752_);
  and (_29215_, _21585_, _21311_);
  or (_29216_, _29215_, _22397_);
  and (_29217_, _26492_, _21629_);
  or (_29218_, _29217_, _29216_);
  or (_29219_, _29218_, _29214_);
  and (_29220_, _29219_, _18521_);
  and (_29221_, _27284_, _29190_);
  not (_29222_, _21059_);
  and (_29223_, _29222_, _29221_);
  and (_29224_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_29225_, _29224_, _29223_);
  or (_29226_, _29225_, _29220_);
  and (_12139_, _29226_, _25964_);
  and (_29227_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], _25964_);
  and (_29228_, _29227_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_29229_, _21026_, _21980_);
  or (_29230_, _26484_, _21837_);
  or (_29231_, _29230_, _29229_);
  and (_29232_, _26492_, _21443_);
  or (_29233_, _29232_, _29231_);
  or (_29234_, _27347_, _26498_);
  and (_29235_, _21026_, _19464_);
  nand (_29236_, _29235_, _19179_);
  nand (_29237_, _29236_, _22331_);
  or (_29238_, _29237_, _29214_);
  or (_29239_, _29238_, _29234_);
  or (_29240_, _29239_, _29233_);
  and (_29241_, _29240_, _28193_);
  or (_12142_, _29241_, _29228_);
  and (_29242_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_29243_, _21267_, _18521_);
  or (_29244_, _29243_, _29242_);
  or (_29245_, _29244_, _29223_);
  and (_12145_, _29245_, _25964_);
  not (_29246_, _27284_);
  and (_29247_, _21443_, _21147_);
  and (_29248_, _27360_, _19464_);
  or (_29249_, _29248_, _29247_);
  and (_29250_, _29249_, _29246_);
  and (_29251_, _20741_, _20785_);
  not (_29252_, _21969_);
  nor (_29253_, _29163_, _29252_);
  nor (_29254_, _29253_, _29251_);
  not (_29255_, _29254_);
  and (_29256_, _29255_, _29221_);
  and (_29257_, _29251_, _19475_);
  and (_29258_, _29257_, _24378_);
  or (_29259_, _29258_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_29260_, _29259_, _29256_);
  or (_29261_, _29260_, _29250_);
  or (_29262_, _15520_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_29263_, _29262_, _25964_);
  and (_12148_, _29263_, _29261_);
  and (_29264_, \oc8051_top_1.oc8051_sfr1.wait_data , _25964_);
  and (_29265_, _29264_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_29266_, _21432_, _21311_);
  and (_29267_, _29266_, _26480_);
  or (_29268_, _21629_, _21443_);
  and (_29269_, _29268_, _21530_);
  or (_29270_, _29269_, _29267_);
  and (_29271_, _21508_, _21147_);
  and (_29272_, _21322_, _20730_);
  or (_29273_, _29232_, _29272_);
  or (_29274_, _29273_, _29271_);
  or (_29275_, _20752_, _21837_);
  or (_29276_, _29215_, _21640_);
  or (_29277_, _29276_, _29275_);
  or (_29278_, _29277_, _29274_);
  or (_29279_, _29278_, _29270_);
  and (_29280_, _29279_, _28193_);
  or (_12151_, _29280_, _29265_);
  and (_29281_, _29264_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_29282_, _21541_, _21169_);
  or (_29283_, _29282_, _22353_);
  and (_29284_, _21530_, _21322_);
  or (_29285_, _29284_, _29283_);
  not (_29286_, _26500_);
  and (_29287_, _26492_, _21750_);
  and (_29288_, _29287_, _21136_);
  or (_29289_, _21827_, _21761_);
  or (_29290_, _29289_, _29288_);
  or (_29291_, _29290_, _29286_);
  or (_29292_, _29291_, _29285_);
  and (_29293_, _21585_, _21169_);
  and (_29294_, _26485_, _19721_);
  or (_29295_, _29294_, _29293_);
  and (_29296_, _20741_, _21366_);
  and (_29297_, _26492_, _21651_);
  or (_29298_, _29297_, _29296_);
  or (_29299_, _29298_, _29295_);
  nor (_29300_, _29217_, _21794_);
  nand (_29301_, _29300_, _21892_);
  or (_29302_, _29301_, _29299_);
  or (_29303_, _29302_, _29233_);
  or (_29304_, _29303_, _29292_);
  and (_29305_, _29304_, _28193_);
  or (_12154_, _29305_, _29281_);
  and (_29306_, _22221_, _20785_);
  and (_29307_, _26492_, _21377_);
  or (_29308_, _29307_, _29306_);
  and (_29309_, _26480_, _20785_);
  or (_29310_, _29309_, _22243_);
  and (_29311_, _21377_, _20708_);
  or (_29312_, _29311_, _29310_);
  or (_29313_, _29312_, _29308_);
  and (_29314_, _26492_, _20796_);
  or (_29315_, _29314_, _29222_);
  or (_29316_, _29315_, _29313_);
  and (_29317_, _29316_, _28193_);
  nor (_29318_, _21059_, _24378_);
  and (_29319_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_29320_, _29319_, _29318_);
  and (_29321_, _29320_, _25964_);
  or (_12157_, _29321_, _29317_);
  not (_29322_, _21278_);
  or (_29323_, _29230_, _29322_);
  or (_29324_, _21640_, _21333_);
  or (_29325_, _29324_, _29247_);
  or (_29326_, _29325_, _29323_);
  and (_29327_, _20818_, _19464_);
  and (_29328_, _29327_, _21256_);
  or (_29329_, _22287_, _21772_);
  or (_29330_, _29329_, _29328_);
  or (_29331_, _21761_, _21201_);
  or (_29332_, _29331_, _29330_);
  nand (_29333_, _21925_, _21706_);
  or (_29334_, _29333_, _29332_);
  or (_29335_, _29334_, _29326_);
  and (_29336_, _21585_, _20785_);
  or (_29337_, _29336_, _29248_);
  and (_29338_, _26480_, _20818_);
  or (_29339_, _29338_, _21596_);
  or (_29340_, _29339_, _29216_);
  or (_29341_, _29340_, _29337_);
  and (_29342_, _29327_, _21530_);
  or (_29343_, _29342_, _22309_);
  or (_29344_, _29343_, _21552_);
  or (_29345_, _29344_, _26498_);
  or (_29346_, _29345_, _29341_);
  or (_29347_, _29346_, _29335_);
  and (_29348_, _29347_, _18521_);
  and (_29349_, _29249_, _20916_);
  or (_29350_, _29349_, _29223_);
  and (_29351_, _20916_, _22090_);
  or (_29352_, _29351_, _29350_);
  and (_29353_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_29354_, _29353_, _29352_);
  or (_29355_, _29354_, _29348_);
  and (_12160_, _29355_, _25964_);
  nor (_12208_, _22550_, rst);
  nor (_12210_, _22166_, rst);
  nand (_12213_, _29255_, _28193_);
  nand (_29356_, _29251_, _28193_);
  not (_29357_, _20949_);
  or (_29358_, _29162_, _29357_);
  and (_12216_, _29358_, _29356_);
  or (_29359_, _29177_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_29360_, _29359_, _29178_);
  or (_29361_, _29360_, _29168_);
  and (_29362_, _29361_, _29192_);
  nor (_29363_, _29191_, _20894_);
  or (_29364_, _29363_, rst);
  or (_12219_, _29364_, _29362_);
  nand (_29365_, _19962_, _18466_);
  or (_29366_, _18466_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_29367_, _29366_, _25964_);
  and (_12222_, _29367_, _29365_);
  not (_29368_, _18466_);
  or (_29369_, _20214_, _29368_);
  or (_29370_, _18466_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_29371_, _29370_, _25964_);
  and (_12225_, _29371_, _29369_);
  nand (_29372_, _20445_, _18466_);
  or (_29373_, _18466_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_29374_, _29373_, _25964_);
  and (_12228_, _29374_, _29372_);
  nand (_29375_, _20686_, _18466_);
  or (_29376_, _18466_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_29377_, _29376_, _25964_);
  and (_12231_, _29377_, _29375_);
  or (_29378_, _19442_, _29368_);
  or (_29379_, _18466_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_29380_, _29379_, _25964_);
  and (_12234_, _29380_, _29378_);
  nand (_29381_, _19699_, _18466_);
  or (_29382_, _18466_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_29383_, _29382_, _25964_);
  and (_12237_, _29383_, _29381_);
  nand (_29384_, _18905_, _18466_);
  or (_29385_, _18466_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_29386_, _29385_, _25964_);
  and (_12240_, _29386_, _29384_);
  or (_29387_, _29287_, _29213_);
  or (_29388_, _29311_, _26481_);
  or (_29389_, _29388_, _29387_);
  not (_29390_, _26497_);
  and (_29391_, _29390_, _21026_);
  or (_29392_, _29294_, _22408_);
  or (_29393_, _29314_, _29307_);
  or (_29394_, _29393_, _29392_);
  or (_29395_, _29394_, _29391_);
  or (_29396_, _29395_, _29389_);
  and (_29397_, _21969_, _21256_);
  or (_29398_, _29310_, _29397_);
  and (_29399_, _29235_, _20818_);
  and (_29400_, _22441_, _21585_);
  or (_29401_, _29400_, _29399_);
  or (_29402_, _29401_, _29398_);
  or (_29403_, _29204_, _26493_);
  or (_29404_, _29403_, _29298_);
  or (_29405_, _20752_, _22353_);
  and (_29406_, _21530_, _21190_);
  or (_29407_, _29406_, _22451_);
  or (_29408_, _29407_, _29405_);
  or (_29409_, _29408_, _29404_);
  or (_29410_, _29409_, _29402_);
  or (_29411_, _29410_, _29396_);
  and (_29412_, _29411_, _18521_);
  and (_29413_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_29414_, _29413_, _29256_);
  or (_29415_, _29414_, _29412_);
  and (_24286_, _29415_, _25964_);
  and (_29416_, _29264_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_29417_, _29257_, _29204_);
  and (_29418_, _21783_, _20708_);
  or (_29419_, _29418_, _22320_);
  and (_29420_, _21026_, _20796_);
  or (_29421_, _29420_, _29419_);
  or (_29422_, _21508_, _21180_);
  and (_29423_, _29422_, _29235_);
  or (_29424_, _29423_, _29295_);
  or (_29425_, _29424_, _29421_);
  or (_29426_, _29425_, _29417_);
  or (_29427_, _29426_, _29285_);
  or (_29428_, _29307_, _21761_);
  or (_29429_, _29428_, _21695_);
  and (_29430_, _29429_, _21136_);
  and (_29431_, _29297_, _21136_);
  not (_29432_, _21673_);
  or (_29433_, _29387_, _29432_);
  or (_29434_, _29433_, _29431_);
  or (_29435_, _29434_, _29430_);
  or (_29436_, _29435_, _29427_);
  and (_29437_, _29436_, _28193_);
  or (_24287_, _29437_, _29416_);
  or (_29438_, _29337_, _29335_);
  and (_29439_, _29438_, _18521_);
  and (_29440_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_29441_, _29440_, _29352_);
  or (_29442_, _29441_, _29439_);
  and (_24288_, _29442_, _25964_);
  and (_29443_, _21684_, _19475_);
  or (_29444_, _29443_, _22397_);
  or (_29445_, _29444_, _29344_);
  or (_29446_, _29445_, _29249_);
  and (_29447_, _29446_, _18521_);
  or (_29448_, _29447_, _29350_);
  and (_29449_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_29450_, _29449_, _29448_);
  and (_24289_, _29450_, _25964_);
  and (_29451_, _29399_, _19157_);
  or (_29452_, _29204_, _27343_);
  or (_29453_, _29452_, _29391_);
  or (_29454_, _29453_, _29451_);
  and (_29455_, _21026_, _21629_);
  or (_29456_, _29314_, _29455_);
  or (_29457_, _29309_, _21037_);
  or (_29458_, _29457_, _22254_);
  or (_29459_, _29458_, _29456_);
  or (_29460_, _29459_, _29454_);
  or (_29461_, _29338_, _22408_);
  or (_29462_, _29461_, _29342_);
  and (_29463_, _29328_, _19157_);
  or (_29464_, _29463_, _20850_);
  or (_29465_, _29464_, _29462_);
  or (_29466_, _29431_, _29288_);
  or (_29467_, _29466_, _29465_);
  and (_29468_, _21026_, _20840_);
  and (_29469_, _21190_, _21147_);
  and (_29470_, _29307_, _19475_);
  or (_29471_, _29470_, _29469_);
  or (_29472_, _29471_, _29468_);
  or (_29473_, _29472_, _29249_);
  or (_29474_, _29388_, _29296_);
  or (_29475_, _26493_, _21048_);
  and (_29476_, _29307_, _19464_);
  or (_29477_, _29476_, _29251_);
  or (_29478_, _29477_, _29475_);
  or (_29479_, _29478_, _29474_);
  or (_29480_, _29479_, _29473_);
  or (_29481_, _29480_, _29467_);
  or (_29482_, _29481_, _29460_);
  and (_29483_, _29482_, _28193_);
  or (_29484_, _29256_, _29318_);
  and (_29485_, _29484_, _25964_);
  and (_29486_, _29264_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_29487_, _29486_, _29485_);
  or (_24290_, _29487_, _29483_);
  or (_29488_, _21048_, _22408_);
  or (_29489_, _29328_, _29213_);
  nor (_29490_, _29489_, _29488_);
  nand (_29491_, _29490_, _20861_);
  not (_29492_, _21256_);
  nor (_29493_, _21958_, _29492_);
  or (_29494_, _21750_, _21651_);
  and (_29495_, _29494_, _20741_);
  or (_29496_, _29495_, _29493_);
  or (_29497_, _29496_, _29491_);
  and (_29498_, _29338_, _19157_);
  and (_29499_, _29342_, _19157_);
  or (_29500_, _29499_, _21201_);
  or (_29501_, _29500_, _29498_);
  or (_29502_, _29501_, _29474_);
  or (_29503_, _29502_, _29497_);
  or (_29504_, _29503_, _29460_);
  and (_29505_, _29504_, _28193_);
  and (_29506_, _29264_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or (_29507_, _29506_, _29485_);
  or (_24291_, _29507_, _29505_);
  and (_29508_, _29264_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_29509_, _20741_, _21443_);
  or (_29510_, _29509_, _29200_);
  or (_29511_, _29270_, _24381_);
  or (_29512_, _29511_, _29510_);
  and (_29513_, _29235_, _29266_);
  or (_29514_, _29513_, _21772_);
  or (_29515_, _29324_, _29275_);
  or (_29516_, _29515_, _29514_);
  and (_29517_, _20741_, _21783_);
  or (_29518_, _29309_, _29215_);
  or (_29519_, _29518_, _29517_);
  and (_29520_, _22221_, _21377_);
  and (_29521_, _20741_, _21421_);
  or (_29522_, _29521_, _29520_);
  or (_29523_, _29522_, _29519_);
  and (_29524_, _21421_, _20708_);
  or (_29525_, _29314_, _22408_);
  or (_29526_, _29525_, _29524_);
  or (_29527_, _29476_, _21223_);
  or (_29528_, _29527_, _29526_);
  or (_29529_, _29528_, _29523_);
  or (_29530_, _29529_, _29516_);
  or (_29531_, _29530_, _29512_);
  and (_29532_, _29531_, _28193_);
  or (_24292_, _29532_, _29508_);
  or (_29533_, _29282_, _29217_);
  or (_29534_, _29470_, _29284_);
  or (_29535_, _29534_, _29533_);
  or (_29536_, _29535_, _29290_);
  or (_29537_, _29536_, _29478_);
  and (_29538_, _29235_, _21311_);
  or (_29539_, _29538_, _29521_);
  or (_29540_, _29388_, _29509_);
  or (_29541_, _29540_, _29539_);
  or (_29542_, _20850_, _21881_);
  or (_29543_, _29293_, _20752_);
  or (_29544_, _29543_, _29542_);
  nand (_29545_, _22265_, _21212_);
  or (_29546_, _29545_, _29544_);
  or (_29547_, _29546_, _29541_);
  or (_29548_, _29547_, _29537_);
  and (_29549_, _29548_, _28193_);
  and (_29550_, _18477_, _25964_);
  and (_29551_, _29550_, _21048_);
  and (_29552_, _29264_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_29553_, _29552_, _29551_);
  or (_24293_, _29553_, _29549_);
  and (_29554_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_29555_, _21048_, _15520_);
  or (_29556_, _29555_, _29554_);
  and (_29557_, _29556_, _25964_);
  and (_29558_, _20741_, _21377_);
  or (_29559_, _22408_, _22397_);
  or (_29560_, _29518_, _29559_);
  nor (_29561_, _29560_, _29558_);
  and (_29562_, _29561_, _26495_);
  or (_29563_, _29517_, _21903_);
  or (_29564_, _29563_, _29451_);
  nor (_29565_, _29564_, _29234_);
  and (_29566_, _29565_, _29562_);
  not (_29567_, _26482_);
  or (_29568_, _22342_, _21870_);
  or (_29569_, _29568_, _29567_);
  or (_29570_, _29314_, _29217_);
  or (_29571_, _29570_, _29452_);
  or (_29572_, _29571_, _29569_);
  nor (_29573_, _29572_, _29233_);
  nand (_29574_, _29573_, _29566_);
  and (_29575_, _29574_, _28193_);
  or (_24294_, _29575_, _29557_);
  or (_29576_, _29276_, _29567_);
  or (_29577_, _29576_, _29514_);
  or (_29578_, _22397_, _22309_);
  or (_29579_, _29578_, _21794_);
  and (_29580_, _20741_, _21432_);
  or (_29581_, _29580_, _26493_);
  or (_29582_, _29581_, _29579_);
  nand (_29583_, _26499_, _21212_);
  or (_29584_, _29583_, _29582_);
  or (_29585_, _29564_, _29231_);
  or (_29586_, _29585_, _29584_);
  or (_29587_, _29586_, _29577_);
  and (_29588_, _29587_, _28193_);
  or (_29589_, _21037_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_29590_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _15520_);
  and (_29591_, _29590_, _25964_);
  and (_29592_, _29591_, _29589_);
  or (_24295_, _29592_, _29588_);
  and (_29593_, _29264_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_29594_, _29314_, _27343_);
  or (_29595_, _29594_, _21344_);
  or (_29596_, _29595_, _24379_);
  or (_29597_, _29539_, _24380_);
  or (_29598_, _29597_, _29596_);
  or (_29599_, _29207_, _29419_);
  or (_29600_, _29599_, _29517_);
  or (_29601_, _29600_, _29313_);
  or (_29602_, _29601_, _29510_);
  or (_29603_, _29602_, _29598_);
  and (_29604_, _29603_, _28193_);
  or (_24297_, _29604_, _29593_);
  not (_29605_, _25847_);
  nor (_29606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_29607_, _29113_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_29608_, _29607_, _29606_);
  nor (_29609_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_29610_, _29117_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_29611_, _29610_, _29609_);
  nor (_29612_, _29611_, _29608_);
  nor (_29613_, _28505_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_29614_, _29121_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_29615_, _29614_, _29613_);
  and (_29616_, _29615_, _29612_);
  nor (_29617_, _28524_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_29618_, _29125_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_29619_, _29618_, _29617_);
  not (_29620_, _29619_);
  and (_29621_, _29620_, _29616_);
  and (_29622_, _29621_, _29605_);
  not (_29623_, _25974_);
  and (_29624_, _29611_, _29608_);
  not (_29625_, _29612_);
  and (_29626_, _29615_, _29625_);
  nor (_29627_, _29615_, _29625_);
  nor (_29628_, _29627_, _29626_);
  not (_29629_, _29628_);
  nor (_29630_, _29619_, _29626_);
  and (_29631_, _29619_, _29626_);
  nor (_29632_, _29631_, _29630_);
  and (_29633_, _29632_, _29629_);
  and (_29634_, _29633_, _29624_);
  and (_29635_, _29634_, _29623_);
  not (_00007_, _25929_);
  not (_00008_, _29611_);
  nor (_00009_, _00008_, _29608_);
  and (_00010_, _29633_, _00009_);
  and (_00011_, _00010_, _00007_);
  or (_00012_, _00011_, _29635_);
  or (_00013_, _00012_, _29622_);
  not (_00014_, _26067_);
  and (_00015_, _00008_, _29608_);
  and (_00016_, _29619_, _29628_);
  and (_00017_, _00016_, _00015_);
  and (_00018_, _00017_, _00014_);
  not (_00019_, _26149_);
  and (_00020_, _00016_, _29624_);
  and (_00021_, _00020_, _00019_);
  not (_00022_, _26108_);
  and (_00023_, _00016_, _00009_);
  and (_00024_, _00023_, _00022_);
  or (_00025_, _00024_, _00021_);
  or (_00026_, _00025_, _00018_);
  not (_00027_, _26023_);
  and (_00028_, _29619_, _29627_);
  and (_00029_, _00028_, _00027_);
  not (_00030_, _25888_);
  and (_00031_, _00015_, _29633_);
  and (_00032_, _00031_, _00030_);
  or (_00033_, _00032_, _00029_);
  or (_00034_, _00033_, _00026_);
  or (_00035_, _00034_, _00013_);
  not (_00036_, _25601_);
  nor (_00037_, _29632_, _29628_);
  and (_00038_, _00037_, _00009_);
  and (_00039_, _00038_, _00036_);
  not (_00040_, _25765_);
  and (_00041_, _29630_, _00009_);
  and (_00042_, _00041_, _00040_);
  not (_00043_, _25806_);
  and (_00044_, _29630_, _29624_);
  and (_00045_, _00044_, _00043_);
  or (_00047_, _00045_, _00042_);
  not (_00049_, _25683_);
  and (_00051_, _29620_, _29627_);
  and (_00053_, _00051_, _00049_);
  not (_00055_, _25724_);
  and (_00057_, _00015_, _29630_);
  and (_00059_, _00057_, _00055_);
  or (_00060_, _00059_, _00053_);
  or (_00061_, _00060_, _00047_);
  or (_00062_, _00061_, _00039_);
  not (_00063_, _26190_);
  and (_00064_, _29619_, _29616_);
  and (_00065_, _00064_, _00063_);
  not (_00067_, _25558_);
  and (_00068_, _00015_, _00037_);
  and (_00070_, _00068_, _00067_);
  not (_00071_, _25642_);
  and (_00072_, _00037_, _29624_);
  and (_00073_, _00072_, _00071_);
  or (_00074_, _00073_, _00070_);
  or (_00075_, _00074_, _00065_);
  or (_00076_, _00075_, _00062_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _00076_, _00035_);
  and (_00077_, _00068_, _00019_);
  and (_00078_, _00023_, _00027_);
  and (_00079_, _00020_, _00014_);
  or (_00080_, _00079_, _00078_);
  or (_00081_, _00080_, _00077_);
  and (_00082_, _29634_, _00030_);
  and (_00083_, _00038_, _00063_);
  or (_00084_, _00083_, _00082_);
  or (_00085_, _00084_, _00081_);
  and (_00086_, _29621_, _00040_);
  and (_00087_, _00044_, _00055_);
  and (_00088_, _00041_, _00049_);
  or (_00089_, _00088_, _00087_);
  or (_00090_, _00089_, _00086_);
  and (_00091_, _00031_, _00043_);
  and (_00092_, _00051_, _00036_);
  or (_00093_, _00092_, _00091_);
  or (_00094_, _00093_, _00090_);
  or (_00095_, _00094_, _00085_);
  and (_00096_, _00064_, _00022_);
  and (_00097_, _00072_, _00067_);
  and (_00099_, _00057_, _00071_);
  or (_00101_, _00099_, _00097_);
  and (_00103_, _00010_, _29605_);
  and (_00105_, _00028_, _00007_);
  and (_00107_, _00017_, _29623_);
  or (_00109_, _00107_, _00105_);
  or (_00111_, _00109_, _00103_);
  or (_00112_, _00111_, _00101_);
  or (_00113_, _00112_, _00096_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _00113_, _00095_);
  and (_00114_, _00010_, _00030_);
  and (_00115_, _00031_, _29605_);
  and (_00116_, _00038_, _00067_);
  or (_00118_, _00116_, _00115_);
  or (_00119_, _00118_, _00114_);
  and (_00121_, _00023_, _00014_);
  and (_00122_, _00017_, _00027_);
  or (_00123_, _00122_, _00121_);
  and (_00124_, _00020_, _00022_);
  and (_00125_, _00028_, _29623_);
  and (_00126_, _00051_, _00071_);
  or (_00127_, _00126_, _00125_);
  and (_00128_, _00064_, _00019_);
  and (_00129_, _29621_, _00043_);
  or (_00130_, _00129_, _00128_);
  or (_00131_, _00130_, _00127_);
  or (_00132_, _00131_, _00124_);
  or (_00133_, _00132_, _00123_);
  and (_00134_, _29634_, _00007_);
  and (_00135_, _00057_, _00049_);
  and (_00136_, _00044_, _00040_);
  and (_00137_, _00041_, _00055_);
  or (_00138_, _00137_, _00136_);
  or (_00139_, _00138_, _00135_);
  or (_00140_, _00139_, _00134_);
  and (_00141_, _00068_, _00063_);
  and (_00142_, _00072_, _00036_);
  or (_00143_, _00142_, _00141_);
  or (_00144_, _00143_, _00140_);
  or (_00145_, _00144_, _00133_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _00145_, _00119_);
  and (_00146_, _29634_, _29605_);
  and (_00147_, _00010_, _00043_);
  and (_00148_, _00068_, _00022_);
  or (_00150_, _00148_, _00147_);
  or (_00152_, _00150_, _00146_);
  and (_00154_, _00017_, _00007_);
  and (_00156_, _00051_, _00067_);
  and (_00158_, _29621_, _00055_);
  or (_00160_, _00158_, _00156_);
  and (_00162_, _00028_, _00030_);
  and (_00163_, _00064_, _00014_);
  or (_00164_, _00163_, _00162_);
  or (_00165_, _00164_, _00160_);
  or (_00166_, _00165_, _00154_);
  and (_00167_, _00023_, _29623_);
  and (_00168_, _00020_, _00027_);
  or (_00170_, _00168_, _00167_);
  or (_00171_, _00170_, _00166_);
  and (_00173_, _00072_, _00063_);
  and (_00174_, _00038_, _00019_);
  or (_00175_, _00174_, _00173_);
  and (_00176_, _00031_, _00040_);
  and (_00177_, _00041_, _00071_);
  and (_00178_, _00057_, _00036_);
  or (_00179_, _00178_, _00177_);
  and (_00180_, _00044_, _00049_);
  or (_00181_, _00180_, _00179_);
  or (_00182_, _00181_, _00176_);
  or (_00183_, _00182_, _00175_);
  or (_00184_, _00183_, _00171_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _00184_, _00152_);
  not (_00185_, _25893_);
  and (_00186_, _00010_, _00185_);
  not (_00187_, _25852_);
  and (_00188_, _00031_, _00187_);
  not (_00189_, _25563_);
  and (_00190_, _00038_, _00189_);
  or (_00191_, _00190_, _00188_);
  or (_00192_, _00191_, _00186_);
  not (_00193_, _26072_);
  and (_00194_, _00023_, _00193_);
  not (_00195_, _26031_);
  and (_00196_, _00017_, _00195_);
  or (_00197_, _00196_, _00194_);
  not (_00198_, _26113_);
  and (_00199_, _00020_, _00198_);
  not (_00200_, _25983_);
  and (_00202_, _00028_, _00200_);
  not (_00204_, _25647_);
  and (_00206_, _00051_, _00204_);
  or (_00208_, _00206_, _00202_);
  not (_00210_, _26154_);
  and (_00212_, _00064_, _00210_);
  not (_00214_, _25811_);
  and (_00215_, _29621_, _00214_);
  or (_00216_, _00215_, _00212_);
  or (_00217_, _00216_, _00208_);
  or (_00218_, _00217_, _00199_);
  or (_00219_, _00218_, _00197_);
  not (_00220_, _25934_);
  and (_00222_, _29634_, _00220_);
  not (_00223_, _25729_);
  and (_00225_, _00041_, _00223_);
  not (_00226_, _25688_);
  and (_00227_, _00057_, _00226_);
  or (_00228_, _00227_, _00225_);
  not (_00229_, _25770_);
  and (_00230_, _00044_, _00229_);
  or (_00231_, _00230_, _00228_);
  or (_00232_, _00231_, _00222_);
  not (_00233_, _26195_);
  and (_00234_, _00068_, _00233_);
  not (_00235_, _25606_);
  and (_00236_, _00072_, _00235_);
  or (_00237_, _00236_, _00234_);
  or (_00238_, _00237_, _00232_);
  or (_00239_, _00238_, _00219_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _00239_, _00192_);
  not (_00240_, _26200_);
  and (_00241_, _00068_, _00240_);
  not (_00242_, _25898_);
  and (_00243_, _00010_, _00242_);
  or (_00244_, _00243_, _00241_);
  not (_00245_, _26118_);
  and (_00246_, _00020_, _00245_);
  not (_00247_, _26036_);
  and (_00248_, _00017_, _00247_);
  not (_00249_, _26077_);
  and (_00250_, _00023_, _00249_);
  or (_00251_, _00250_, _00248_);
  or (_00252_, _00251_, _00246_);
  or (_00254_, _00252_, _00244_);
  not (_00256_, _25734_);
  and (_00258_, _00041_, _00256_);
  not (_00260_, _25816_);
  and (_00262_, _29621_, _00260_);
  not (_00264_, _25775_);
  and (_00266_, _00044_, _00264_);
  or (_00267_, _00266_, _00262_);
  or (_00268_, _00267_, _00258_);
  not (_00269_, _25611_);
  and (_00270_, _00072_, _00269_);
  not (_00271_, _25693_);
  and (_00272_, _00057_, _00271_);
  or (_00274_, _00272_, _00270_);
  or (_00275_, _00274_, _00268_);
  or (_00277_, _00275_, _00254_);
  not (_00278_, _25857_);
  and (_00279_, _00031_, _00278_);
  not (_00280_, _25939_);
  and (_00281_, _29634_, _00280_);
  not (_00282_, _25988_);
  and (_00283_, _00028_, _00282_);
  or (_00284_, _00283_, _00281_);
  or (_00285_, _00284_, _00279_);
  not (_00286_, _26159_);
  and (_00287_, _00064_, _00286_);
  not (_00288_, _25568_);
  and (_00289_, _00038_, _00288_);
  not (_00290_, _25652_);
  and (_00291_, _00051_, _00290_);
  or (_00292_, _00291_, _00289_);
  or (_00293_, _00292_, _00287_);
  or (_00294_, _00293_, _00285_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _00294_, _00277_);
  not (_00295_, _25944_);
  and (_00296_, _29634_, _00295_);
  not (_00297_, _25862_);
  and (_00298_, _00031_, _00297_);
  not (_00299_, _25616_);
  and (_00300_, _00072_, _00299_);
  or (_00301_, _00300_, _00298_);
  or (_00302_, _00301_, _00296_);
  not (_00303_, _26041_);
  and (_00304_, _00017_, _00303_);
  not (_00306_, _26164_);
  and (_00308_, _00064_, _00306_);
  not (_00310_, _25821_);
  and (_00312_, _29621_, _00310_);
  or (_00314_, _00312_, _00308_);
  not (_00316_, _25993_);
  and (_00318_, _00028_, _00316_);
  not (_00319_, _25657_);
  and (_00320_, _00051_, _00319_);
  or (_00321_, _00320_, _00318_);
  or (_00322_, _00321_, _00314_);
  or (_00323_, _00322_, _00304_);
  not (_00324_, _26082_);
  and (_00326_, _00023_, _00324_);
  not (_00327_, _26123_);
  and (_00329_, _00020_, _00327_);
  or (_00330_, _00329_, _00326_);
  or (_00331_, _00330_, _00323_);
  not (_00332_, _25903_);
  and (_00333_, _00010_, _00332_);
  not (_00334_, _25739_);
  and (_00335_, _00041_, _00334_);
  not (_00336_, _25780_);
  and (_00337_, _00044_, _00336_);
  not (_00338_, _25698_);
  and (_00339_, _00057_, _00338_);
  or (_00340_, _00339_, _00337_);
  or (_00341_, _00340_, _00335_);
  or (_00342_, _00341_, _00333_);
  not (_00343_, _26205_);
  and (_00344_, _00068_, _00343_);
  not (_00345_, _25575_);
  and (_00346_, _00038_, _00345_);
  or (_00347_, _00346_, _00344_);
  or (_00348_, _00347_, _00342_);
  or (_00349_, _00348_, _00331_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _00349_, _00302_);
  not (_00350_, _26210_);
  and (_00351_, _00068_, _00350_);
  not (_00352_, _25867_);
  and (_00353_, _00031_, _00352_);
  not (_00354_, _25580_);
  and (_00355_, _00038_, _00354_);
  or (_00356_, _00355_, _00353_);
  or (_00358_, _00356_, _00351_);
  not (_00360_, _26087_);
  and (_00362_, _00023_, _00360_);
  not (_00364_, _26046_);
  and (_00366_, _00017_, _00364_);
  or (_00368_, _00366_, _00362_);
  not (_00370_, _26128_);
  and (_00371_, _00020_, _00370_);
  not (_00372_, _25826_);
  and (_00373_, _29621_, _00372_);
  not (_00374_, _25662_);
  and (_00375_, _00051_, _00374_);
  or (_00376_, _00375_, _00373_);
  not (_00378_, _26169_);
  and (_00379_, _00064_, _00378_);
  not (_00381_, _25998_);
  and (_00382_, _00028_, _00381_);
  or (_00383_, _00382_, _00379_);
  or (_00384_, _00383_, _00376_);
  or (_00385_, _00384_, _00371_);
  or (_00386_, _00385_, _00368_);
  not (_00387_, _25621_);
  and (_00388_, _00072_, _00387_);
  not (_00389_, _25703_);
  and (_00390_, _00057_, _00389_);
  not (_00391_, _25785_);
  and (_00392_, _00044_, _00391_);
  not (_00393_, _25744_);
  and (_00394_, _00041_, _00393_);
  or (_00395_, _00394_, _00392_);
  or (_00396_, _00395_, _00390_);
  or (_00397_, _00396_, _00388_);
  not (_00398_, _25949_);
  and (_00399_, _29634_, _00398_);
  not (_00400_, _25908_);
  and (_00401_, _00010_, _00400_);
  or (_00402_, _00401_, _00399_);
  or (_00403_, _00402_, _00397_);
  or (_00404_, _00403_, _00386_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _00404_, _00358_);
  not (_00405_, _25872_);
  and (_00406_, _00031_, _00405_);
  not (_00407_, _25585_);
  and (_00408_, _00038_, _00407_);
  not (_00410_, _25954_);
  and (_00412_, _29634_, _00410_);
  or (_00414_, _00412_, _00408_);
  or (_00416_, _00414_, _00406_);
  not (_00418_, _26051_);
  and (_00420_, _00017_, _00418_);
  not (_00422_, _25667_);
  and (_00423_, _00051_, _00422_);
  not (_00424_, _26003_);
  and (_00425_, _00028_, _00424_);
  or (_00426_, _00425_, _00423_);
  not (_00427_, _25831_);
  and (_00428_, _29621_, _00427_);
  not (_00430_, _26174_);
  and (_00431_, _00064_, _00430_);
  or (_00433_, _00431_, _00428_);
  or (_00434_, _00433_, _00426_);
  or (_00435_, _00434_, _00420_);
  not (_00436_, _26092_);
  and (_00437_, _00023_, _00436_);
  not (_00438_, _26133_);
  and (_00439_, _00020_, _00438_);
  or (_00440_, _00439_, _00437_);
  or (_00441_, _00440_, _00435_);
  not (_00442_, _26215_);
  and (_00443_, _00068_, _00442_);
  not (_00444_, _25708_);
  and (_00445_, _00057_, _00444_);
  not (_00446_, _25749_);
  and (_00447_, _00041_, _00446_);
  or (_00448_, _00447_, _00445_);
  not (_00449_, _25790_);
  and (_00450_, _00044_, _00449_);
  or (_00451_, _00450_, _00448_);
  or (_00452_, _00451_, _00443_);
  not (_00453_, _25626_);
  and (_00454_, _00072_, _00453_);
  not (_00455_, _25913_);
  and (_00456_, _00010_, _00455_);
  or (_00457_, _00456_, _00454_);
  or (_00458_, _00457_, _00452_);
  or (_00459_, _00458_, _00441_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _00459_, _00416_);
  not (_00460_, _26220_);
  and (_00462_, _00068_, _00460_);
  not (_00464_, _25918_);
  and (_00466_, _00010_, _00464_);
  or (_00468_, _00466_, _00462_);
  not (_00470_, _26138_);
  and (_00472_, _00020_, _00470_);
  not (_00474_, _26056_);
  and (_00475_, _00017_, _00474_);
  not (_00476_, _26097_);
  and (_00477_, _00023_, _00476_);
  or (_00478_, _00477_, _00475_);
  or (_00479_, _00478_, _00472_);
  or (_00480_, _00479_, _00468_);
  not (_00482_, _25754_);
  and (_00483_, _00041_, _00482_);
  not (_00485_, _25836_);
  and (_00486_, _29621_, _00485_);
  not (_00487_, _25795_);
  and (_00488_, _00044_, _00487_);
  or (_00489_, _00488_, _00486_);
  or (_00490_, _00489_, _00483_);
  not (_00491_, _25631_);
  and (_00492_, _00072_, _00491_);
  not (_00493_, _25713_);
  and (_00494_, _00057_, _00493_);
  or (_00495_, _00494_, _00492_);
  or (_00496_, _00495_, _00490_);
  or (_00497_, _00496_, _00480_);
  not (_00498_, _25877_);
  and (_00499_, _00031_, _00498_);
  not (_00500_, _25959_);
  and (_00501_, _29634_, _00500_);
  not (_00502_, _26008_);
  and (_00503_, _00028_, _00502_);
  or (_00504_, _00503_, _00501_);
  or (_00505_, _00504_, _00499_);
  not (_00506_, _26179_);
  and (_00507_, _00064_, _00506_);
  not (_00508_, _25590_);
  and (_00509_, _00038_, _00508_);
  not (_00510_, _25672_);
  and (_00511_, _00051_, _00510_);
  or (_00512_, _00511_, _00509_);
  or (_00513_, _00512_, _00507_);
  or (_00515_, _00513_, _00505_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _00515_, _00497_);
  not (_00518_, _25965_);
  and (_00520_, _29634_, _00518_);
  not (_00522_, _26225_);
  and (_00524_, _00068_, _00522_);
  not (_00526_, _25923_);
  and (_00527_, _00010_, _00526_);
  or (_00528_, _00527_, _00524_);
  or (_00529_, _00528_, _00520_);
  not (_00530_, _26061_);
  and (_00531_, _00017_, _00530_);
  not (_00532_, _26102_);
  and (_00534_, _00023_, _00532_);
  or (_00535_, _00534_, _00531_);
  not (_00537_, _26143_);
  and (_00538_, _00020_, _00537_);
  not (_00539_, _25677_);
  and (_00540_, _00051_, _00539_);
  not (_00541_, _26184_);
  and (_00542_, _00064_, _00541_);
  or (_00543_, _00542_, _00540_);
  not (_00544_, _25841_);
  and (_00545_, _29621_, _00544_);
  not (_00546_, _26013_);
  and (_00547_, _00028_, _00546_);
  or (_00548_, _00547_, _00545_);
  or (_00549_, _00548_, _00543_);
  or (_00550_, _00549_, _00538_);
  or (_00551_, _00550_, _00535_);
  not (_00552_, _25636_);
  and (_00553_, _00072_, _00552_);
  not (_00554_, _25718_);
  and (_00555_, _00057_, _00554_);
  not (_00556_, _25800_);
  and (_00557_, _00044_, _00556_);
  not (_00558_, _25759_);
  and (_00559_, _00041_, _00558_);
  or (_00560_, _00559_, _00557_);
  or (_00561_, _00560_, _00555_);
  or (_00562_, _00561_, _00553_);
  not (_00563_, _25595_);
  and (_00564_, _00038_, _00563_);
  not (_00565_, _25882_);
  and (_00567_, _00031_, _00565_);
  or (_00569_, _00567_, _00564_);
  or (_00571_, _00569_, _00562_);
  or (_00573_, _00571_, _00551_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _00573_, _00529_);
  and (_00576_, _00068_, _00210_);
  and (_00578_, _00023_, _00195_);
  and (_00579_, _00020_, _00193_);
  or (_00580_, _00579_, _00578_);
  or (_00581_, _00580_, _00576_);
  and (_00582_, _29634_, _00185_);
  and (_00583_, _00038_, _00233_);
  or (_00584_, _00583_, _00582_);
  or (_00586_, _00584_, _00581_);
  and (_00587_, _29621_, _00229_);
  and (_00589_, _00044_, _00223_);
  and (_00590_, _00041_, _00226_);
  or (_00591_, _00590_, _00589_);
  or (_00592_, _00591_, _00587_);
  and (_00593_, _00031_, _00214_);
  and (_00594_, _00051_, _00235_);
  or (_00595_, _00594_, _00593_);
  or (_00596_, _00595_, _00592_);
  or (_00597_, _00596_, _00586_);
  and (_00598_, _00064_, _00198_);
  and (_00599_, _00072_, _00189_);
  and (_00600_, _00057_, _00204_);
  or (_00601_, _00600_, _00599_);
  and (_00602_, _00010_, _00187_);
  and (_00603_, _00028_, _00220_);
  and (_00604_, _00017_, _00200_);
  or (_00605_, _00604_, _00603_);
  or (_00606_, _00605_, _00602_);
  or (_00607_, _00606_, _00601_);
  or (_00608_, _00607_, _00598_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _00608_, _00597_);
  and (_00609_, _00068_, _00286_);
  and (_00610_, _00023_, _00247_);
  and (_00611_, _00020_, _00249_);
  or (_00612_, _00611_, _00610_);
  or (_00613_, _00612_, _00609_);
  and (_00614_, _29634_, _00242_);
  and (_00615_, _00038_, _00240_);
  or (_00616_, _00615_, _00614_);
  or (_00618_, _00616_, _00613_);
  and (_00620_, _29621_, _00264_);
  and (_00622_, _00041_, _00271_);
  and (_00624_, _00044_, _00256_);
  or (_00626_, _00624_, _00622_);
  or (_00628_, _00626_, _00620_);
  and (_00630_, _00051_, _00269_);
  and (_00631_, _00031_, _00260_);
  or (_00632_, _00631_, _00630_);
  or (_00633_, _00632_, _00628_);
  or (_00634_, _00633_, _00618_);
  and (_00635_, _00064_, _00245_);
  and (_00636_, _00072_, _00288_);
  and (_00638_, _00057_, _00290_);
  or (_00639_, _00638_, _00636_);
  and (_00641_, _00010_, _00278_);
  and (_00642_, _00028_, _00280_);
  and (_00643_, _00017_, _00282_);
  or (_00644_, _00643_, _00642_);
  or (_00645_, _00644_, _00641_);
  or (_00646_, _00645_, _00639_);
  or (_00647_, _00646_, _00635_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _00647_, _00634_);
  and (_00648_, _00028_, _00295_);
  and (_00649_, _00017_, _00316_);
  or (_00650_, _00649_, _00648_);
  and (_00651_, _00010_, _00297_);
  and (_00652_, _29634_, _00332_);
  or (_00653_, _00652_, _00651_);
  or (_00654_, _00653_, _00650_);
  and (_00655_, _29621_, _00336_);
  and (_00656_, _00041_, _00338_);
  and (_00657_, _00044_, _00334_);
  or (_00658_, _00657_, _00656_);
  or (_00659_, _00658_, _00655_);
  and (_00660_, _00031_, _00310_);
  and (_00661_, _00051_, _00299_);
  or (_00662_, _00661_, _00660_);
  or (_00663_, _00662_, _00659_);
  or (_00664_, _00663_, _00654_);
  and (_00665_, _00038_, _00343_);
  and (_00666_, _00068_, _00306_);
  and (_00667_, _00023_, _00303_);
  and (_00668_, _00020_, _00324_);
  or (_00670_, _00668_, _00667_);
  or (_00672_, _00670_, _00666_);
  or (_00674_, _00672_, _00665_);
  and (_00676_, _00064_, _00327_);
  and (_00678_, _00057_, _00319_);
  and (_00680_, _00072_, _00345_);
  or (_00682_, _00680_, _00678_);
  or (_00683_, _00682_, _00676_);
  or (_00684_, _00683_, _00674_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _00684_, _00664_);
  and (_00685_, _00068_, _00378_);
  and (_00686_, _00023_, _00364_);
  and (_00687_, _00020_, _00360_);
  or (_00689_, _00687_, _00686_);
  or (_00690_, _00689_, _00685_);
  and (_00692_, _00010_, _00352_);
  and (_00693_, _00038_, _00350_);
  or (_00694_, _00693_, _00692_);
  or (_00695_, _00694_, _00690_);
  and (_00696_, _29621_, _00391_);
  and (_00697_, _00044_, _00393_);
  and (_00698_, _00041_, _00389_);
  or (_00699_, _00698_, _00697_);
  or (_00700_, _00699_, _00696_);
  and (_00701_, _00031_, _00372_);
  and (_00702_, _00051_, _00387_);
  or (_00703_, _00702_, _00701_);
  or (_00704_, _00703_, _00700_);
  or (_00705_, _00704_, _00695_);
  and (_00706_, _00064_, _00370_);
  and (_00707_, _00072_, _00354_);
  and (_00708_, _00057_, _00374_);
  or (_00709_, _00708_, _00707_);
  and (_00710_, _29634_, _00400_);
  and (_00711_, _00028_, _00398_);
  and (_00712_, _00017_, _00381_);
  or (_00713_, _00712_, _00711_);
  or (_00714_, _00713_, _00710_);
  or (_00715_, _00714_, _00709_);
  or (_00716_, _00715_, _00706_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _00716_, _00705_);
  and (_00717_, _00017_, _00424_);
  and (_00718_, _00028_, _00410_);
  or (_00719_, _00718_, _00717_);
  and (_00721_, _29634_, _00455_);
  and (_00723_, _00010_, _00405_);
  or (_00725_, _00723_, _00721_);
  or (_00727_, _00725_, _00719_);
  and (_00729_, _29621_, _00449_);
  and (_00731_, _00044_, _00446_);
  and (_00733_, _00041_, _00444_);
  or (_00734_, _00733_, _00731_);
  or (_00735_, _00734_, _00729_);
  and (_00736_, _00051_, _00453_);
  and (_00737_, _00031_, _00427_);
  or (_00738_, _00737_, _00736_);
  or (_00739_, _00738_, _00735_);
  or (_00741_, _00739_, _00727_);
  and (_00742_, _00038_, _00442_);
  and (_00744_, _00023_, _00418_);
  and (_00745_, _00020_, _00436_);
  or (_00746_, _00745_, _00744_);
  and (_00747_, _00068_, _00430_);
  or (_00748_, _00747_, _00746_);
  or (_00749_, _00748_, _00742_);
  and (_00750_, _00064_, _00438_);
  and (_00751_, _00072_, _00407_);
  and (_00752_, _00057_, _00422_);
  or (_00753_, _00752_, _00751_);
  or (_00754_, _00753_, _00750_);
  or (_00755_, _00754_, _00749_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _00755_, _00741_);
  and (_00756_, _00041_, _00493_);
  and (_00757_, _00044_, _00482_);
  or (_00758_, _00757_, _00756_);
  and (_00759_, _00031_, _00485_);
  and (_00760_, _29621_, _00487_);
  or (_00761_, _00760_, _00759_);
  or (_00762_, _00761_, _00758_);
  and (_00763_, _00068_, _00506_);
  and (_00764_, _00023_, _00474_);
  and (_00765_, _00020_, _00476_);
  or (_00766_, _00765_, _00764_);
  or (_00767_, _00766_, _00763_);
  and (_00768_, _29634_, _00464_);
  and (_00769_, _00038_, _00460_);
  or (_00770_, _00769_, _00768_);
  or (_00771_, _00770_, _00767_);
  or (_00773_, _00771_, _00762_);
  and (_00775_, _00072_, _00508_);
  and (_00777_, _00051_, _00491_);
  and (_00779_, _00057_, _00510_);
  or (_00781_, _00779_, _00777_);
  or (_00783_, _00781_, _00775_);
  and (_00785_, _00064_, _00470_);
  and (_00786_, _00010_, _00498_);
  and (_00787_, _00028_, _00500_);
  and (_00788_, _00017_, _00502_);
  or (_00789_, _00788_, _00787_);
  or (_00790_, _00789_, _00786_);
  or (_00791_, _00790_, _00785_);
  or (_00793_, _00791_, _00783_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _00793_, _00773_);
  and (_00795_, _00038_, _00522_);
  and (_00796_, _00010_, _00565_);
  or (_00797_, _00796_, _00795_);
  and (_00798_, _00068_, _00541_);
  and (_00799_, _00020_, _00532_);
  and (_00800_, _00023_, _00530_);
  or (_00801_, _00800_, _00799_);
  or (_00802_, _00801_, _00798_);
  or (_00803_, _00802_, _00797_);
  and (_00804_, _29621_, _00556_);
  and (_00805_, _00044_, _00558_);
  and (_00806_, _00041_, _00554_);
  or (_00807_, _00806_, _00805_);
  or (_00808_, _00807_, _00804_);
  and (_00809_, _00031_, _00544_);
  and (_00810_, _00051_, _00552_);
  or (_00811_, _00810_, _00809_);
  or (_00812_, _00811_, _00808_);
  or (_00813_, _00812_, _00803_);
  and (_00814_, _00064_, _00537_);
  and (_00815_, _00072_, _00563_);
  and (_00816_, _00057_, _00539_);
  or (_00817_, _00816_, _00815_);
  and (_00818_, _29634_, _00526_);
  and (_00819_, _00017_, _00546_);
  and (_00820_, _00028_, _00518_);
  or (_00821_, _00820_, _00819_);
  or (_00822_, _00821_, _00818_);
  or (_00823_, _00822_, _00817_);
  or (_00825_, _00823_, _00814_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _00825_, _00813_);
  and (_00828_, _00010_, _00220_);
  and (_00830_, _29634_, _00200_);
  or (_00832_, _00830_, _00828_);
  and (_00834_, _00031_, _00185_);
  and (_00836_, _29621_, _00187_);
  or (_00837_, _00836_, _00834_);
  or (_00838_, _00837_, _00832_);
  and (_00839_, _00051_, _00226_);
  and (_00840_, _00041_, _00229_);
  and (_00841_, _00044_, _00214_);
  or (_00842_, _00841_, _00840_);
  or (_00844_, _00842_, _00839_);
  and (_00845_, _00038_, _00235_);
  and (_00847_, _00057_, _00223_);
  or (_00848_, _00847_, _00845_);
  or (_00849_, _00848_, _00844_);
  or (_00850_, _00849_, _00838_);
  and (_00851_, _00023_, _00198_);
  and (_00852_, _00020_, _00210_);
  or (_00853_, _00852_, _00851_);
  and (_00854_, _00017_, _00193_);
  and (_00855_, _00028_, _00195_);
  or (_00856_, _00855_, _00854_);
  or (_00857_, _00856_, _00853_);
  and (_00858_, _00064_, _00233_);
  and (_00859_, _00072_, _00204_);
  and (_00860_, _00068_, _00189_);
  or (_00861_, _00860_, _00859_);
  or (_00862_, _00861_, _00858_);
  or (_00863_, _00862_, _00857_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _00863_, _00850_);
  and (_00864_, _00031_, _00242_);
  and (_00865_, _00010_, _00280_);
  and (_00866_, _00038_, _00269_);
  or (_00867_, _00866_, _00865_);
  or (_00868_, _00867_, _00864_);
  and (_00869_, _00023_, _00245_);
  and (_00870_, _00020_, _00286_);
  or (_00871_, _00870_, _00869_);
  and (_00872_, _00017_, _00249_);
  and (_00873_, _00028_, _00247_);
  and (_00874_, _29621_, _00278_);
  or (_00876_, _00874_, _00873_);
  and (_00878_, _00064_, _00240_);
  and (_00880_, _00051_, _00271_);
  or (_00882_, _00880_, _00878_);
  or (_00884_, _00882_, _00876_);
  or (_00886_, _00884_, _00872_);
  or (_00888_, _00886_, _00871_);
  and (_00889_, _00068_, _00288_);
  and (_00890_, _00072_, _00290_);
  or (_00891_, _00890_, _00889_);
  and (_00892_, _29634_, _00282_);
  and (_00893_, _00041_, _00264_);
  and (_00894_, _00044_, _00260_);
  or (_00895_, _00894_, _00893_);
  and (_00896_, _00057_, _00256_);
  or (_00897_, _00896_, _00895_);
  or (_00898_, _00897_, _00892_);
  or (_00899_, _00898_, _00891_);
  or (_00900_, _00899_, _00888_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _00900_, _00868_);
  and (_00901_, _00023_, _00327_);
  and (_00902_, _00020_, _00306_);
  or (_00903_, _00902_, _00901_);
  and (_00904_, _00028_, _00303_);
  or (_00905_, _00904_, _00903_);
  and (_00906_, _00017_, _00324_);
  and (_00907_, _29621_, _00297_);
  or (_00908_, _00907_, _00906_);
  or (_00909_, _00908_, _00905_);
  and (_00910_, _00051_, _00338_);
  and (_00911_, _00044_, _00310_);
  and (_00912_, _00041_, _00336_);
  or (_00913_, _00912_, _00911_);
  or (_00914_, _00913_, _00910_);
  and (_00915_, _00057_, _00334_);
  and (_00916_, _00038_, _00299_);
  or (_00917_, _00916_, _00915_);
  or (_00919_, _00917_, _00914_);
  or (_00920_, _00919_, _00909_);
  and (_00921_, _00031_, _00332_);
  and (_00923_, _29634_, _00316_);
  and (_00924_, _00010_, _00295_);
  or (_00925_, _00924_, _00923_);
  or (_00927_, _00925_, _00921_);
  and (_00928_, _00068_, _00345_);
  and (_00929_, _00072_, _00319_);
  or (_00930_, _00929_, _00928_);
  and (_00931_, _00064_, _00343_);
  or (_00932_, _00931_, _00930_);
  or (_00933_, _00932_, _00927_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _00933_, _00920_);
  and (_00934_, _00028_, _00364_);
  and (_00935_, _00020_, _00378_);
  and (_00936_, _00023_, _00370_);
  or (_00937_, _00936_, _00935_);
  or (_00938_, _00937_, _00934_);
  and (_00939_, _29621_, _00352_);
  and (_00940_, _00017_, _00360_);
  or (_00941_, _00940_, _00939_);
  or (_00942_, _00941_, _00938_);
  and (_00943_, _00051_, _00389_);
  and (_00944_, _00041_, _00391_);
  and (_00945_, _00044_, _00372_);
  or (_00946_, _00945_, _00944_);
  or (_00947_, _00946_, _00943_);
  and (_00948_, _00038_, _00387_);
  and (_00949_, _00057_, _00393_);
  or (_00950_, _00949_, _00948_);
  or (_00951_, _00950_, _00947_);
  or (_00952_, _00951_, _00942_);
  and (_00953_, _00031_, _00400_);
  and (_00954_, _00010_, _00398_);
  and (_00955_, _29634_, _00381_);
  or (_00956_, _00955_, _00954_);
  or (_00957_, _00956_, _00953_);
  and (_00958_, _00064_, _00350_);
  and (_00959_, _00072_, _00374_);
  and (_00960_, _00068_, _00354_);
  or (_00961_, _00960_, _00959_);
  or (_00962_, _00961_, _00958_);
  or (_00963_, _00962_, _00957_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _00963_, _00952_);
  and (_00964_, _00010_, _00410_);
  and (_00965_, _00072_, _00422_);
  and (_00966_, _00038_, _00453_);
  or (_00967_, _00966_, _00965_);
  or (_00968_, _00967_, _00964_);
  and (_00969_, _00020_, _00430_);
  and (_00970_, _00023_, _00438_);
  or (_00971_, _00970_, _00969_);
  and (_00972_, _00017_, _00436_);
  and (_00973_, _29621_, _00405_);
  and (_00974_, _00051_, _00444_);
  or (_00975_, _00974_, _00973_);
  and (_00976_, _00064_, _00442_);
  and (_00977_, _00028_, _00418_);
  or (_00978_, _00977_, _00976_);
  or (_00979_, _00978_, _00975_);
  or (_00980_, _00979_, _00972_);
  or (_00981_, _00980_, _00971_);
  and (_00982_, _00031_, _00455_);
  and (_00983_, _00057_, _00446_);
  and (_00984_, _00044_, _00427_);
  and (_00985_, _00041_, _00449_);
  or (_00986_, _00985_, _00984_);
  or (_00987_, _00986_, _00983_);
  or (_00988_, _00987_, _00982_);
  and (_00989_, _29634_, _00424_);
  and (_00990_, _00068_, _00407_);
  or (_00991_, _00990_, _00989_);
  or (_00992_, _00991_, _00988_);
  or (_00993_, _00992_, _00981_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _00993_, _00968_);
  and (_00994_, _00031_, _00464_);
  and (_00995_, _00010_, _00500_);
  and (_00996_, _00038_, _00491_);
  or (_00997_, _00996_, _00995_);
  or (_00998_, _00997_, _00994_);
  and (_00999_, _00023_, _00470_);
  and (_01000_, _00028_, _00474_);
  and (_01001_, _29621_, _00498_);
  or (_01002_, _01001_, _01000_);
  and (_01003_, _00064_, _00460_);
  and (_01004_, _00051_, _00493_);
  or (_01005_, _01004_, _01003_);
  or (_01006_, _01005_, _01002_);
  or (_01007_, _01006_, _00999_);
  and (_01008_, _00020_, _00506_);
  and (_01009_, _00017_, _00476_);
  or (_01010_, _01009_, _01008_);
  or (_01011_, _01010_, _01007_);
  and (_01012_, _00068_, _00508_);
  and (_01013_, _00072_, _00510_);
  or (_01014_, _01013_, _01012_);
  and (_01015_, _29634_, _00502_);
  and (_01016_, _00044_, _00485_);
  and (_01017_, _00041_, _00487_);
  or (_01018_, _01017_, _01016_);
  and (_01019_, _00057_, _00482_);
  or (_01020_, _01019_, _01018_);
  or (_01021_, _01020_, _01015_);
  or (_01022_, _01021_, _01014_);
  or (_01023_, _01022_, _01011_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _01023_, _00998_);
  and (_01024_, _29634_, _00546_);
  and (_01025_, _00031_, _00526_);
  and (_01026_, _00038_, _00552_);
  or (_01027_, _01026_, _01025_);
  or (_01028_, _01027_, _01024_);
  and (_01029_, _00023_, _00537_);
  and (_01030_, _00064_, _00522_);
  and (_01031_, _29621_, _00565_);
  or (_01032_, _01031_, _01030_);
  and (_01033_, _00028_, _00530_);
  and (_01034_, _00051_, _00554_);
  or (_01035_, _01034_, _01033_);
  or (_01036_, _01035_, _01032_);
  or (_01037_, _01036_, _01029_);
  and (_01038_, _00020_, _00541_);
  and (_01039_, _00017_, _00532_);
  or (_01040_, _01039_, _01038_);
  or (_01041_, _01040_, _01037_);
  and (_01042_, _00068_, _00563_);
  and (_01043_, _00072_, _00539_);
  or (_01044_, _01043_, _01042_);
  and (_01045_, _00010_, _00518_);
  and (_01046_, _00041_, _00556_);
  and (_01048_, _00044_, _00544_);
  or (_01049_, _01048_, _01046_);
  and (_01051_, _00057_, _00558_);
  or (_01052_, _01051_, _01049_);
  or (_01054_, _01052_, _01045_);
  or (_01055_, _01054_, _01044_);
  or (_01057_, _01055_, _01041_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _01057_, _01028_);
  and (_01059_, _00038_, _00210_);
  and (_01060_, _00068_, _00198_);
  and (_01062_, _00031_, _00229_);
  or (_01063_, _01062_, _01060_);
  or (_01065_, _01063_, _01059_);
  and (_01066_, _00023_, _00200_);
  and (_01068_, _00064_, _00193_);
  and (_01069_, _00051_, _00189_);
  or (_01071_, _01069_, _01068_);
  and (_01072_, _00028_, _00185_);
  and (_01074_, _29621_, _00223_);
  or (_01075_, _01074_, _01072_);
  or (_01077_, _01075_, _01071_);
  or (_01078_, _01077_, _01066_);
  and (_01080_, _00020_, _00195_);
  and (_01081_, _00017_, _00220_);
  or (_01083_, _01081_, _01080_);
  or (_01084_, _01083_, _01078_);
  and (_01086_, _29634_, _00187_);
  and (_01087_, _00057_, _00235_);
  and (_01089_, _00041_, _00204_);
  or (_01090_, _01089_, _01087_);
  and (_01092_, _00044_, _00226_);
  or (_01093_, _01092_, _01090_);
  or (_01095_, _01093_, _01086_);
  and (_01096_, _00072_, _00233_);
  and (_01098_, _00010_, _00214_);
  or (_01099_, _01098_, _01096_);
  or (_01101_, _01099_, _01095_);
  or (_01102_, _01101_, _01084_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _01102_, _01065_);
  and (_01104_, _29634_, _00278_);
  and (_01106_, _00023_, _00282_);
  and (_01107_, _00017_, _00280_);
  or (_01108_, _01107_, _01106_);
  or (_01109_, _01108_, _01104_);
  and (_01110_, _00028_, _00242_);
  and (_01111_, _00068_, _00245_);
  or (_01112_, _01111_, _01110_);
  or (_01113_, _01112_, _01109_);
  and (_01114_, _00010_, _00260_);
  and (_01115_, _00057_, _00269_);
  and (_01116_, _00051_, _00288_);
  and (_01117_, _00041_, _00290_);
  or (_01118_, _01117_, _01116_);
  or (_01119_, _01118_, _01115_);
  or (_01120_, _01119_, _01114_);
  or (_01121_, _01120_, _01113_);
  and (_01122_, _00020_, _00247_);
  and (_01123_, _00072_, _00240_);
  and (_01124_, _00038_, _00286_);
  or (_01125_, _01124_, _01123_);
  or (_01126_, _01125_, _01122_);
  and (_01127_, _00064_, _00249_);
  and (_01128_, _00031_, _00264_);
  and (_01129_, _29621_, _00256_);
  and (_01130_, _00044_, _00271_);
  or (_01131_, _01130_, _01129_);
  or (_01132_, _01131_, _01128_);
  or (_01133_, _01132_, _01127_);
  or (_01134_, _01133_, _01126_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _01134_, _01121_);
  and (_01135_, _29634_, _00297_);
  and (_01136_, _00010_, _00310_);
  and (_01137_, _00068_, _00327_);
  or (_01138_, _01137_, _01136_);
  or (_01139_, _01138_, _01135_);
  and (_01140_, _00017_, _00295_);
  and (_01141_, _00051_, _00345_);
  and (_01142_, _29621_, _00334_);
  or (_01143_, _01142_, _01141_);
  and (_01144_, _00028_, _00332_);
  and (_01145_, _00064_, _00324_);
  or (_01146_, _01145_, _01144_);
  or (_01147_, _01146_, _01143_);
  or (_01148_, _01147_, _01140_);
  and (_01149_, _00023_, _00316_);
  and (_01150_, _00020_, _00303_);
  or (_01151_, _01150_, _01149_);
  or (_01152_, _01151_, _01148_);
  and (_01153_, _00072_, _00343_);
  and (_01154_, _00038_, _00306_);
  or (_01155_, _01154_, _01153_);
  and (_01156_, _00031_, _00336_);
  and (_01157_, _00041_, _00319_);
  and (_01158_, _00057_, _00299_);
  or (_01159_, _01158_, _01157_);
  and (_01160_, _00044_, _00338_);
  or (_01161_, _01160_, _01159_);
  or (_01162_, _01161_, _01156_);
  or (_01163_, _01162_, _01155_);
  or (_01164_, _01163_, _01152_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _01164_, _01139_);
  and (_01165_, _00010_, _00372_);
  and (_01166_, _00031_, _00391_);
  and (_01167_, _00068_, _00370_);
  or (_01168_, _01167_, _01166_);
  or (_01169_, _01168_, _01165_);
  and (_01170_, _00017_, _00398_);
  and (_01171_, _00023_, _00381_);
  or (_01172_, _01171_, _01170_);
  and (_01173_, _00020_, _00364_);
  and (_01174_, _00051_, _00354_);
  and (_01175_, _00064_, _00360_);
  or (_01176_, _01175_, _01174_);
  and (_01177_, _29621_, _00393_);
  and (_01178_, _00028_, _00400_);
  or (_01179_, _01178_, _01177_);
  or (_01180_, _01179_, _01176_);
  or (_01181_, _01180_, _01173_);
  or (_01182_, _01181_, _01172_);
  and (_01183_, _00038_, _00378_);
  and (_01184_, _00057_, _00387_);
  and (_01185_, _00041_, _00374_);
  or (_01186_, _01185_, _01184_);
  and (_01187_, _00044_, _00389_);
  or (_01188_, _01187_, _01186_);
  or (_01189_, _01188_, _01183_);
  and (_01190_, _00072_, _00350_);
  and (_01191_, _29634_, _00352_);
  or (_01192_, _01191_, _01190_);
  or (_01193_, _01192_, _01189_);
  or (_01194_, _01193_, _01182_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _01194_, _01169_);
  and (_01195_, _00010_, _00427_);
  and (_01196_, _00038_, _00430_);
  and (_01197_, _00031_, _00449_);
  or (_01198_, _01197_, _01196_);
  or (_01199_, _01198_, _01195_);
  and (_01200_, _00017_, _00410_);
  and (_01201_, _00064_, _00436_);
  and (_01202_, _00028_, _00455_);
  or (_01203_, _01202_, _01201_);
  and (_01204_, _00051_, _00407_);
  and (_01205_, _29621_, _00446_);
  or (_01206_, _01205_, _01204_);
  or (_01207_, _01206_, _01203_);
  or (_01208_, _01207_, _01200_);
  and (_01209_, _00020_, _00418_);
  and (_01210_, _00023_, _00424_);
  or (_01211_, _01210_, _01209_);
  or (_01212_, _01211_, _01208_);
  and (_01213_, _00068_, _00438_);
  and (_01214_, _00041_, _00422_);
  and (_01215_, _00057_, _00453_);
  and (_01216_, _00044_, _00444_);
  or (_01217_, _01216_, _01215_);
  or (_01218_, _01217_, _01214_);
  or (_01219_, _01218_, _01213_);
  and (_01220_, _00072_, _00442_);
  and (_01221_, _29634_, _00405_);
  or (_01222_, _01221_, _01220_);
  or (_01223_, _01222_, _01219_);
  or (_01224_, _01223_, _01212_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _01224_, _01199_);
  and (_01225_, _29634_, _00498_);
  and (_01226_, _00023_, _00502_);
  and (_01227_, _00017_, _00500_);
  or (_01228_, _01227_, _01226_);
  or (_01229_, _01228_, _01225_);
  and (_01230_, _00028_, _00464_);
  and (_01231_, _00020_, _00474_);
  or (_01232_, _01231_, _01230_);
  or (_01233_, _01232_, _01229_);
  and (_01234_, _00010_, _00485_);
  and (_01235_, _00057_, _00491_);
  and (_01236_, _00051_, _00508_);
  and (_01237_, _00041_, _00510_);
  or (_01238_, _01237_, _01236_);
  or (_01239_, _01238_, _01235_);
  or (_01240_, _01239_, _01234_);
  or (_01241_, _01240_, _01233_);
  and (_01242_, _00068_, _00470_);
  and (_01243_, _00072_, _00460_);
  and (_01244_, _00038_, _00506_);
  or (_01245_, _01244_, _01243_);
  or (_01246_, _01245_, _01242_);
  and (_01247_, _00064_, _00476_);
  and (_01248_, _00031_, _00487_);
  and (_01249_, _29621_, _00482_);
  and (_01250_, _00044_, _00493_);
  or (_01251_, _01250_, _01249_);
  or (_01252_, _01251_, _01248_);
  or (_01253_, _01252_, _01247_);
  or (_01254_, _01253_, _01246_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _01254_, _01241_);
  and (_01255_, _29634_, _00565_);
  and (_01256_, _00010_, _00544_);
  and (_01257_, _00068_, _00537_);
  or (_01258_, _01257_, _01256_);
  or (_01259_, _01258_, _01255_);
  and (_01260_, _00017_, _00518_);
  and (_01261_, _00051_, _00563_);
  and (_01262_, _29621_, _00558_);
  or (_01263_, _01262_, _01261_);
  and (_01264_, _00028_, _00526_);
  and (_01265_, _00064_, _00532_);
  or (_01266_, _01265_, _01264_);
  or (_01267_, _01266_, _01263_);
  or (_01268_, _01267_, _01260_);
  and (_01269_, _00023_, _00546_);
  and (_01270_, _00020_, _00530_);
  or (_01271_, _01270_, _01269_);
  or (_01272_, _01271_, _01268_);
  and (_01273_, _00072_, _00522_);
  and (_01274_, _00038_, _00541_);
  or (_01275_, _01274_, _01273_);
  and (_01276_, _00031_, _00556_);
  and (_01277_, _00041_, _00539_);
  and (_01278_, _00057_, _00552_);
  or (_01279_, _01278_, _01277_);
  and (_01280_, _00044_, _00554_);
  or (_01281_, _01280_, _01279_);
  or (_01282_, _01281_, _01276_);
  or (_01283_, _01282_, _01275_);
  or (_01284_, _01283_, _01272_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _01284_, _01259_);
  and (_01285_, _26506_, \oc8051_golden_model_1.P3INREG [7]);
  or (_01286_, _01285_, _26818_);
  and (_25303_, _01286_, _25964_);
  and (_01287_, _26506_, \oc8051_golden_model_1.P2INREG [7]);
  or (_01288_, _01287_, _26632_);
  and (_25304_, _01288_, _25964_);
  and (_01289_, _26506_, \oc8051_golden_model_1.P1INREG [7]);
  or (_01290_, _01289_, _26753_);
  and (_25306_, _01290_, _25964_);
  and (_01291_, _26506_, \oc8051_golden_model_1.P0INREG [7]);
  or (_01292_, _01291_, _26541_);
  and (_25307_, _01292_, _25964_);
  nand (_01293_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_01294_, \oc8051_golden_model_1.PC [3]);
  or (_01295_, \oc8051_golden_model_1.PC [2], _01294_);
  or (_01296_, _01295_, _01293_);
  or (_01297_, _01296_, _26041_);
  not (_01298_, \oc8051_golden_model_1.PC [1]);
  or (_01299_, _01298_, \oc8051_golden_model_1.PC [0]);
  or (_01300_, _01299_, _01295_);
  or (_01301_, _01300_, _25993_);
  and (_01302_, _01301_, _01297_);
  not (_01303_, \oc8051_golden_model_1.PC [2]);
  or (_01304_, _01303_, \oc8051_golden_model_1.PC [3]);
  or (_01305_, _01304_, _01293_);
  or (_01306_, _01305_, _25862_);
  or (_01307_, _01304_, _01299_);
  or (_01308_, _01307_, _25821_);
  and (_01309_, _01308_, _01306_);
  and (_01310_, _01309_, _01302_);
  nand (_01311_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_01312_, _01311_, _01293_);
  or (_01313_, _01312_, _26205_);
  or (_01314_, _01311_, _01299_);
  or (_01315_, _01314_, _26164_);
  and (_01316_, _01315_, _01313_);
  or (_01317_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_01318_, _01317_, _01293_);
  or (_01319_, _01318_, _25698_);
  or (_01320_, _01317_, _01299_);
  or (_01321_, _01320_, _25657_);
  and (_01322_, _01321_, _01319_);
  and (_01323_, _01322_, _01316_);
  and (_01324_, _01323_, _01310_);
  not (_01325_, \oc8051_golden_model_1.PC [0]);
  or (_01326_, \oc8051_golden_model_1.PC [1], _01325_);
  or (_01327_, _01326_, _01311_);
  or (_01328_, _01327_, _26123_);
  or (_01329_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_01330_, _01329_, _01311_);
  or (_01331_, _01330_, _26082_);
  and (_01332_, _01331_, _01328_);
  or (_01333_, _01317_, _01329_);
  or (_01334_, _01333_, _25575_);
  or (_01335_, _01317_, _01326_);
  or (_01336_, _01335_, _25616_);
  and (_01337_, _01336_, _01334_);
  and (_01338_, _01337_, _01332_);
  or (_01339_, _01326_, _01295_);
  or (_01340_, _01339_, _25944_);
  or (_01341_, _01329_, _01295_);
  or (_01342_, _01341_, _25903_);
  and (_01343_, _01342_, _01340_);
  or (_01344_, _01326_, _01304_);
  or (_01345_, _01344_, _25780_);
  or (_01346_, _01329_, _01304_);
  or (_01347_, _01346_, _25739_);
  and (_01348_, _01347_, _01345_);
  and (_01349_, _01348_, _01343_);
  and (_01350_, _01349_, _01338_);
  nand (_01351_, _01350_, _01324_);
  or (_01352_, _01296_, _26046_);
  or (_01353_, _01300_, _25998_);
  and (_01354_, _01353_, _01352_);
  or (_01355_, _01305_, _25867_);
  or (_01356_, _01307_, _25826_);
  and (_01357_, _01356_, _01355_);
  and (_01358_, _01357_, _01354_);
  or (_01359_, _01312_, _26210_);
  or (_01360_, _01314_, _26169_);
  and (_01361_, _01360_, _01359_);
  or (_01362_, _01318_, _25703_);
  or (_01363_, _01320_, _25662_);
  and (_01364_, _01363_, _01362_);
  and (_01365_, _01364_, _01361_);
  and (_01366_, _01365_, _01358_);
  or (_01367_, _01327_, _26128_);
  or (_01368_, _01330_, _26087_);
  and (_01369_, _01368_, _01367_);
  or (_01370_, _01333_, _25580_);
  or (_01371_, _01335_, _25621_);
  and (_01372_, _01371_, _01370_);
  and (_01373_, _01372_, _01369_);
  or (_01374_, _01339_, _25949_);
  or (_01375_, _01341_, _25908_);
  and (_01376_, _01375_, _01374_);
  or (_01377_, _01344_, _25785_);
  or (_01378_, _01346_, _25744_);
  and (_01379_, _01378_, _01377_);
  and (_01380_, _01379_, _01376_);
  and (_01381_, _01380_, _01373_);
  nand (_01382_, _01381_, _01366_);
  or (_01383_, _01382_, _01351_);
  or (_01384_, _01296_, _26031_);
  or (_01385_, _01300_, _25983_);
  and (_01386_, _01385_, _01384_);
  or (_01387_, _01305_, _25852_);
  or (_01388_, _01307_, _25811_);
  and (_01389_, _01388_, _01387_);
  and (_01390_, _01389_, _01386_);
  or (_01391_, _01312_, _26195_);
  or (_01392_, _01314_, _26154_);
  and (_01393_, _01392_, _01391_);
  or (_01394_, _01318_, _25688_);
  or (_01395_, _01320_, _25647_);
  and (_01396_, _01395_, _01394_);
  and (_01397_, _01396_, _01393_);
  and (_01398_, _01397_, _01390_);
  or (_01399_, _01327_, _26113_);
  or (_01400_, _01330_, _26072_);
  and (_01401_, _01400_, _01399_);
  or (_01402_, _01333_, _25563_);
  or (_01403_, _01335_, _25606_);
  and (_01404_, _01403_, _01402_);
  and (_01405_, _01404_, _01401_);
  or (_01406_, _01339_, _25934_);
  or (_01407_, _01341_, _25893_);
  and (_01408_, _01407_, _01406_);
  or (_01409_, _01344_, _25770_);
  or (_01410_, _01346_, _25729_);
  and (_01411_, _01410_, _01409_);
  and (_01412_, _01411_, _01408_);
  and (_01413_, _01412_, _01405_);
  and (_01414_, _01413_, _01398_);
  or (_01415_, _01296_, _26036_);
  or (_01416_, _01300_, _25988_);
  and (_01417_, _01416_, _01415_);
  or (_01418_, _01305_, _25857_);
  or (_01419_, _01307_, _25816_);
  and (_01420_, _01419_, _01418_);
  and (_01421_, _01420_, _01417_);
  or (_01422_, _01312_, _26200_);
  or (_01423_, _01314_, _26159_);
  and (_01424_, _01423_, _01422_);
  or (_01425_, _01318_, _25693_);
  or (_01426_, _01320_, _25652_);
  and (_01427_, _01426_, _01425_);
  and (_01428_, _01427_, _01424_);
  and (_01429_, _01428_, _01421_);
  or (_01430_, _01327_, _26118_);
  or (_01431_, _01330_, _26077_);
  and (_01432_, _01431_, _01430_);
  or (_01433_, _01333_, _25568_);
  or (_01434_, _01335_, _25611_);
  and (_01435_, _01434_, _01433_);
  and (_01436_, _01435_, _01432_);
  or (_01437_, _01339_, _25939_);
  or (_01438_, _01341_, _25898_);
  and (_01439_, _01438_, _01437_);
  or (_01440_, _01344_, _25775_);
  or (_01441_, _01346_, _25734_);
  and (_01442_, _01441_, _01440_);
  and (_01443_, _01442_, _01439_);
  and (_01444_, _01443_, _01436_);
  nand (_01445_, _01444_, _01429_);
  or (_01446_, _01445_, _01414_);
  or (_01447_, _01446_, _01383_);
  not (_01448_, _01447_);
  or (_01449_, _01296_, _26061_);
  or (_01450_, _01300_, _26013_);
  and (_01451_, _01450_, _01449_);
  or (_01452_, _01305_, _25882_);
  or (_01453_, _01307_, _25841_);
  and (_01454_, _01453_, _01452_);
  and (_01455_, _01454_, _01451_);
  or (_01456_, _01312_, _26225_);
  or (_01457_, _01314_, _26184_);
  and (_01458_, _01457_, _01456_);
  or (_01459_, _01318_, _25718_);
  or (_01460_, _01320_, _25677_);
  and (_01461_, _01460_, _01459_);
  and (_01462_, _01461_, _01458_);
  and (_01463_, _01462_, _01455_);
  or (_01464_, _01327_, _26143_);
  or (_01465_, _01330_, _26102_);
  and (_01466_, _01465_, _01464_);
  or (_01467_, _01333_, _25595_);
  or (_01468_, _01335_, _25636_);
  and (_01469_, _01468_, _01467_);
  and (_01470_, _01469_, _01466_);
  or (_01471_, _01339_, _25965_);
  or (_01472_, _01341_, _25923_);
  and (_01473_, _01472_, _01471_);
  or (_01474_, _01344_, _25800_);
  or (_01475_, _01346_, _25759_);
  and (_01476_, _01475_, _01474_);
  and (_01477_, _01476_, _01473_);
  and (_01478_, _01477_, _01470_);
  and (_01479_, _01478_, _01463_);
  or (_01480_, _01296_, _26023_);
  or (_01481_, _01300_, _25974_);
  and (_01482_, _01481_, _01480_);
  or (_01483_, _01305_, _25847_);
  or (_01484_, _01307_, _25806_);
  and (_01485_, _01484_, _01483_);
  and (_01486_, _01485_, _01482_);
  or (_01487_, _01312_, _26190_);
  or (_01488_, _01314_, _26149_);
  and (_01489_, _01488_, _01487_);
  or (_01490_, _01318_, _25683_);
  or (_01491_, _01320_, _25642_);
  and (_01492_, _01491_, _01490_);
  and (_01493_, _01492_, _01489_);
  and (_01494_, _01493_, _01486_);
  or (_01495_, _01327_, _26108_);
  or (_01496_, _01330_, _26067_);
  and (_01497_, _01496_, _01495_);
  or (_01498_, _01333_, _25558_);
  or (_01499_, _01335_, _25601_);
  and (_01500_, _01499_, _01498_);
  and (_01501_, _01500_, _01497_);
  or (_01502_, _01339_, _25929_);
  or (_01503_, _01341_, _25888_);
  and (_01504_, _01503_, _01502_);
  or (_01505_, _01344_, _25765_);
  or (_01506_, _01346_, _25724_);
  and (_01507_, _01506_, _01505_);
  and (_01508_, _01507_, _01504_);
  and (_01509_, _01508_, _01501_);
  and (_01510_, _01509_, _01494_);
  and (_01511_, _01510_, _01479_);
  or (_01512_, _01296_, _26051_);
  or (_01513_, _01300_, _26003_);
  and (_01514_, _01513_, _01512_);
  or (_01515_, _01305_, _25872_);
  or (_01516_, _01307_, _25831_);
  and (_01517_, _01516_, _01515_);
  and (_01518_, _01517_, _01514_);
  or (_01519_, _01312_, _26215_);
  or (_01521_, _01314_, _26174_);
  and (_01523_, _01521_, _01519_);
  or (_01525_, _01318_, _25708_);
  or (_01526_, _01320_, _25667_);
  and (_01528_, _01526_, _01525_);
  and (_01529_, _01528_, _01523_);
  and (_01530_, _01529_, _01518_);
  or (_01531_, _01327_, _26133_);
  or (_01532_, _01330_, _26092_);
  and (_01533_, _01532_, _01531_);
  or (_01534_, _01333_, _25585_);
  or (_01535_, _01335_, _25626_);
  and (_01536_, _01535_, _01534_);
  and (_01537_, _01536_, _01533_);
  or (_01538_, _01339_, _25954_);
  or (_01539_, _01341_, _25913_);
  and (_01540_, _01539_, _01538_);
  or (_01541_, _01344_, _25790_);
  or (_01542_, _01346_, _25749_);
  and (_01543_, _01542_, _01541_);
  and (_01544_, _01543_, _01540_);
  and (_01545_, _01544_, _01537_);
  nand (_01546_, _01545_, _01530_);
  or (_01547_, _01296_, _26056_);
  or (_01548_, _01300_, _26008_);
  and (_01549_, _01548_, _01547_);
  or (_01550_, _01305_, _25877_);
  or (_01551_, _01307_, _25836_);
  and (_01552_, _01551_, _01550_);
  and (_01553_, _01552_, _01549_);
  or (_01554_, _01312_, _26220_);
  or (_01555_, _01314_, _26179_);
  and (_01556_, _01555_, _01554_);
  or (_01557_, _01318_, _25713_);
  or (_01558_, _01320_, _25672_);
  and (_01559_, _01558_, _01557_);
  and (_01560_, _01559_, _01556_);
  and (_01561_, _01560_, _01553_);
  or (_01562_, _01327_, _26138_);
  or (_01563_, _01330_, _26097_);
  and (_01564_, _01563_, _01562_);
  or (_01565_, _01333_, _25590_);
  or (_01566_, _01335_, _25631_);
  and (_01567_, _01566_, _01565_);
  and (_01568_, _01567_, _01564_);
  or (_01569_, _01339_, _25959_);
  or (_01570_, _01341_, _25918_);
  and (_01571_, _01570_, _01569_);
  or (_01572_, _01344_, _25795_);
  or (_01573_, _01346_, _25754_);
  and (_01574_, _01573_, _01572_);
  and (_01575_, _01574_, _01571_);
  and (_01576_, _01575_, _01568_);
  and (_01577_, _01576_, _01561_);
  or (_01578_, _01577_, _01546_);
  not (_01579_, _01578_);
  and (_01580_, _01579_, _01511_);
  and (_01581_, _01580_, _01448_);
  not (_01582_, _01383_);
  and (_01583_, _01445_, _01414_);
  and (_01584_, _01583_, _01582_);
  and (_01585_, _01584_, _01580_);
  nand (_01586_, _01576_, _01561_);
  or (_01587_, _01586_, _01546_);
  not (_01588_, _01587_);
  and (_01589_, _01511_, _01588_);
  not (_01590_, _01446_);
  not (_01591_, _01382_);
  and (_01592_, _01591_, _01351_);
  and (_01593_, _01592_, _01590_);
  and (_01594_, _01593_, _01589_);
  not (_01595_, _01594_);
  not (_01596_, _01585_);
  and (_01597_, _01593_, _01580_);
  nand (_01598_, _01478_, _01463_);
  or (_01599_, _01510_, _01598_);
  nor (_01601_, _01599_, _01587_);
  and (_01602_, _01601_, _01593_);
  and (_01603_, _01545_, _01530_);
  or (_01604_, _01586_, _01603_);
  nor (_01605_, _01604_, _01599_);
  and (_01606_, _01605_, _01448_);
  nor (_01607_, _01606_, _01602_);
  not (_01608_, _01414_);
  and (_01609_, _01445_, _01608_);
  and (_01610_, _01609_, _01582_);
  and (_01611_, _01605_, _01610_);
  and (_01612_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_01613_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_01614_, _01613_, _01612_);
  and (_01615_, _01614_, _01611_);
  not (_01616_, _01611_);
  or (_01617_, _01599_, _01578_);
  or (_01618_, _01617_, _01447_);
  or (_01619_, _01510_, _01479_);
  or (_01620_, _01619_, _01604_);
  or (_01621_, _01620_, _01447_);
  and (_01622_, _01621_, _01618_);
  or (_01623_, _01577_, _01603_);
  or (_01624_, _01623_, _01619_);
  or (_01625_, _01624_, _01447_);
  or (_01626_, _01619_, _01578_);
  or (_01627_, _01626_, _01447_);
  and (_01628_, _01627_, _01625_);
  or (_01629_, _01619_, _01587_);
  or (_01630_, _01629_, _01447_);
  or (_01631_, _01623_, _01599_);
  or (_01632_, _01631_, _01447_);
  and (_01633_, _01632_, _01630_);
  and (_01634_, _01633_, _01628_);
  nand (_01635_, _01634_, _01622_);
  or (_01636_, _01635_, _01325_);
  and (_01637_, _01634_, _01622_);
  or (_01638_, _01637_, \oc8051_golden_model_1.PC [0]);
  and (_01639_, _01638_, _01636_);
  and (_01640_, _01639_, _01616_);
  nor (_01641_, _01640_, _01615_);
  nand (_01642_, _01641_, _01607_);
  and (_01643_, _01601_, _01610_);
  nor (_01644_, _01607_, \oc8051_golden_model_1.PC [0]);
  nor (_01645_, _01644_, _01643_);
  nand (_01646_, _01645_, _01642_);
  not (_01647_, _01623_);
  and (_01648_, _01510_, _01598_);
  and (_01649_, _01648_, _01647_);
  and (_01650_, _01649_, _01448_);
  not (_01651_, _01650_);
  and (_01652_, _01648_, _01579_);
  and (_01653_, _01652_, _01448_);
  and (_01654_, _01601_, _01448_);
  nor (_01655_, _01654_, _01653_);
  and (_01656_, _01655_, _01651_);
  and (_01657_, _01448_, _01589_);
  not (_01658_, _01657_);
  and (_01659_, _01647_, _01511_);
  and (_01660_, _01659_, _01448_);
  nor (_01661_, _01660_, _01581_);
  and (_01662_, _01648_, _01588_);
  and (_01663_, _01662_, _01448_);
  not (_01664_, _01604_);
  and (_01665_, _01648_, _01664_);
  and (_01666_, _01665_, _01448_);
  nor (_01667_, _01666_, _01663_);
  and (_01668_, _01667_, _01661_);
  and (_01669_, _01664_, _01511_);
  and (_01670_, _01669_, _01448_);
  not (_01671_, _01670_);
  and (_01672_, _01671_, _01668_);
  and (_01673_, _01672_, _01658_);
  and (_01674_, _01673_, _01656_);
  not (_01675_, _01674_);
  and (_01676_, \oc8051_golden_model_1.ACC [0], _01325_);
  not (_01677_, _01676_);
  not (_01678_, _01643_);
  not (_01679_, \oc8051_golden_model_1.ACC [0]);
  and (_01680_, _01679_, \oc8051_golden_model_1.PC [0]);
  nor (_01681_, _01680_, _01678_);
  and (_01682_, _01681_, _01677_);
  nor (_01683_, _01682_, _01675_);
  and (_01684_, _01683_, _01646_);
  nor (_01685_, _01674_, \oc8051_golden_model_1.PC [0]);
  or (_01686_, _01685_, _01684_);
  and (_01687_, _01607_, _01637_);
  nand (_01688_, _01687_, _01674_);
  nand (_01689_, _01688_, _01298_);
  and (_01690_, _01326_, _01299_);
  or (_01691_, _01690_, _01635_);
  nand (_01692_, _01691_, _01616_);
  not (_01693_, _01607_);
  and (_01694_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_01695_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_01696_, _01695_, _01694_);
  and (_01697_, _01696_, _01612_);
  nor (_01698_, _01696_, _01612_);
  nor (_01699_, _01698_, _01697_);
  not (_01700_, _01699_);
  and (_01701_, _01700_, _01611_);
  nor (_01702_, _01701_, _01693_);
  nand (_01703_, _01702_, _01692_);
  nand (_01704_, _01703_, _01678_);
  not (_01705_, \oc8051_golden_model_1.ACC [1]);
  nor (_01706_, _01690_, _01705_);
  and (_01707_, _01690_, _01705_);
  nor (_01708_, _01707_, _01706_);
  and (_01709_, _01708_, _01676_);
  nor (_01710_, _01708_, _01676_);
  nor (_01711_, _01710_, _01709_);
  nor (_01712_, _01711_, _01678_);
  nor (_01713_, _01712_, _01675_);
  nand (_01714_, _01713_, _01704_);
  and (_01715_, _01714_, _01689_);
  or (_01716_, _01715_, _01686_);
  and (_01717_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  and (_01718_, _01717_, \oc8051_golden_model_1.PC [3]);
  nor (_01719_, _01717_, \oc8051_golden_model_1.PC [3]);
  nor (_01720_, _01719_, _01718_);
  or (_01721_, _01720_, _01674_);
  nor (_01722_, _01293_, _01303_);
  and (_01723_, _01293_, _01303_);
  nor (_01724_, _01723_, _01722_);
  and (_01725_, _01724_, \oc8051_golden_model_1.ACC [2]);
  nor (_01726_, _01709_, _01706_);
  nor (_01727_, _01724_, \oc8051_golden_model_1.ACC [2]);
  nor (_01728_, _01727_, _01725_);
  not (_01729_, _01728_);
  nor (_01730_, _01729_, _01726_);
  nor (_01731_, _01730_, _01725_);
  not (_01732_, \oc8051_golden_model_1.ACC [3]);
  not (_01733_, _01305_);
  nor (_01734_, _01722_, _01294_);
  nor (_01735_, _01734_, _01733_);
  nor (_01736_, _01735_, _01732_);
  and (_01737_, _01735_, _01732_);
  nor (_01738_, _01737_, _01736_);
  and (_01739_, _01738_, _01731_);
  nor (_01740_, _01738_, _01731_);
  nor (_01741_, _01740_, _01739_);
  nor (_01742_, _01741_, _01678_);
  or (_01743_, _01720_, _01687_);
  and (_01744_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_01745_, _01697_, _01694_);
  nor (_01746_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_01747_, _01746_, _01744_);
  not (_01748_, _01747_);
  nor (_01749_, _01748_, _01745_);
  nor (_01750_, _01749_, _01744_);
  and (_01751_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_01752_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_01753_, _01752_, _01751_);
  not (_01754_, _01753_);
  nor (_01755_, _01754_, _01750_);
  and (_01756_, _01754_, _01750_);
  nor (_01757_, _01756_, _01755_);
  nand (_01758_, _01757_, _01611_);
  and (_01759_, _01758_, _01607_);
  not (_01760_, _01735_);
  or (_01761_, _01635_, _01760_);
  nand (_01762_, _01761_, _01616_);
  nand (_01763_, _01762_, _01759_);
  and (_01764_, _01763_, _01678_);
  or (_01765_, _01764_, _01675_);
  and (_01766_, _01765_, _01743_);
  or (_01767_, _01766_, _01742_);
  nand (_01768_, _01767_, _01721_);
  nor (_01769_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_01770_, _01769_, _01717_);
  nor (_01771_, _01770_, _01687_);
  nor (_01772_, _01724_, _01611_);
  and (_01773_, _01772_, _01637_);
  and (_01774_, _01748_, _01745_);
  nor (_01775_, _01774_, _01749_);
  not (_01776_, _01775_);
  and (_01777_, _01776_, _01611_);
  or (_01778_, _01777_, _01773_);
  and (_01779_, _01778_, _01607_);
  or (_01780_, _01779_, _01643_);
  or (_01781_, _01780_, _01771_);
  and (_01782_, _01729_, _01726_);
  nor (_01783_, _01782_, _01730_);
  and (_01784_, _01783_, _01643_);
  not (_01785_, _01784_);
  and (_01786_, _01785_, _01656_);
  nand (_01787_, _01786_, _01781_);
  not (_01788_, _01673_);
  nor (_01789_, _01770_, _01656_);
  nor (_01790_, _01789_, _01788_);
  nand (_01791_, _01790_, _01787_);
  not (_01792_, _01770_);
  nor (_01793_, _01792_, _01673_);
  not (_01794_, _01793_);
  and (_01795_, _01794_, _01791_);
  or (_01796_, _01795_, _01768_);
  nor (_01797_, _01796_, _01716_);
  nand (_01798_, _01797_, _00063_);
  and (_01799_, _01767_, _01721_);
  nand (_01800_, _01794_, _01791_);
  or (_01801_, _01800_, _01799_);
  nand (_01802_, _01714_, _01689_);
  or (_01803_, _01802_, _01686_);
  or (_01804_, _01803_, _01801_);
  or (_01805_, _01804_, _25601_);
  and (_01806_, _01805_, _01798_);
  or (_01807_, _01800_, _01768_);
  or (_01808_, _01807_, _01716_);
  or (_01809_, _01808_, _26023_);
  or (_01810_, _01801_, _01716_);
  or (_01811_, _01810_, _25683_);
  and (_01812_, _01811_, _01809_);
  and (_01813_, _01812_, _01806_);
  or (_01814_, _01807_, _01803_);
  or (_01815_, _01814_, _25929_);
  nor (_01816_, _01685_, _01684_);
  or (_01817_, _01715_, _01816_);
  or (_01818_, _01817_, _01801_);
  or (_01819_, _01818_, _25642_);
  and (_01820_, _01819_, _01815_);
  or (_01821_, _01795_, _01799_);
  or (_01822_, _01821_, _01716_);
  or (_01823_, _01822_, _25847_);
  or (_01824_, _01803_, _01821_);
  or (_01825_, _01824_, _25765_);
  and (_01826_, _01825_, _01823_);
  and (_01827_, _01826_, _01820_);
  and (_01828_, _01827_, _01813_);
  or (_01829_, _01802_, _01816_);
  or (_01830_, _01829_, _01821_);
  or (_01831_, _01830_, _25724_);
  or (_01832_, _01829_, _01801_);
  or (_01833_, _01832_, _25558_);
  and (_01834_, _01833_, _01831_);
  or (_01835_, _01796_, _01803_);
  or (_01836_, _01835_, _26108_);
  or (_01837_, _01817_, _01807_);
  or (_01838_, _01837_, _25974_);
  and (_01839_, _01838_, _01836_);
  and (_01840_, _01839_, _01834_);
  or (_01841_, _01817_, _01796_);
  or (_01842_, _01841_, _26149_);
  or (_01843_, _01829_, _01807_);
  or (_01844_, _01843_, _25888_);
  and (_01845_, _01844_, _01842_);
  or (_01846_, _01829_, _01796_);
  or (_01847_, _01846_, _26067_);
  or (_01848_, _01817_, _01821_);
  or (_01849_, _01848_, _25806_);
  and (_01850_, _01849_, _01847_);
  and (_01851_, _01850_, _01845_);
  and (_01852_, _01851_, _01840_);
  and (_01853_, _01852_, _01828_);
  nor (_01854_, _01822_, _25882_);
  nor (_01855_, _01804_, _25636_);
  nor (_01856_, _01855_, _01854_);
  nor (_01857_, _01841_, _26184_);
  nor (_01858_, _01810_, _25718_);
  nor (_01859_, _01858_, _01857_);
  and (_01860_, _01859_, _01856_);
  nor (_01861_, _01835_, _26143_);
  nor (_01862_, _01846_, _26102_);
  nor (_01863_, _01862_, _01861_);
  nor (_01864_, _01848_, _25841_);
  nor (_01865_, _01830_, _25759_);
  nor (_01866_, _01865_, _01864_);
  and (_01867_, _01866_, _01863_);
  and (_01868_, _01867_, _01860_);
  nor (_01869_, _01837_, _26013_);
  nor (_01870_, _01843_, _25923_);
  nor (_01871_, _01870_, _01869_);
  nor (_01872_, _01832_, _25595_);
  nor (_01873_, _01818_, _25677_);
  nor (_01874_, _01873_, _01872_);
  and (_01875_, _01874_, _01871_);
  and (_01876_, _01797_, _00522_);
  nor (_01877_, _01824_, _25800_);
  nor (_01878_, _01877_, _01876_);
  nor (_01879_, _01808_, _26061_);
  nor (_01880_, _01814_, _25965_);
  nor (_01881_, _01880_, _01879_);
  and (_01882_, _01881_, _01878_);
  and (_01883_, _01882_, _01875_);
  and (_01884_, _01883_, _01868_);
  and (_01885_, _01884_, _01853_);
  or (_01886_, _01822_, _25867_);
  or (_01887_, _01810_, _25703_);
  and (_01888_, _01887_, _01886_);
  or (_01889_, _01835_, _26128_);
  or (_01890_, _01843_, _25908_);
  and (_01891_, _01890_, _01889_);
  and (_01892_, _01891_, _01888_);
  or (_01893_, _01818_, _25662_);
  or (_01894_, _01804_, _25621_);
  and (_01895_, _01894_, _01893_);
  or (_01896_, _01824_, _25785_);
  or (_01897_, _01830_, _25744_);
  and (_01898_, _01897_, _01896_);
  and (_01899_, _01898_, _01895_);
  and (_01900_, _01899_, _01892_);
  or (_01901_, _01808_, _26046_);
  or (_01902_, _01837_, _25998_);
  and (_01903_, _01902_, _01901_);
  or (_01904_, _01841_, _26169_);
  or (_01905_, _01814_, _25949_);
  and (_01906_, _01905_, _01904_);
  and (_01907_, _01906_, _01903_);
  or (_01908_, _01848_, _25826_);
  or (_01909_, _01832_, _25580_);
  and (_01910_, _01909_, _01908_);
  nand (_01911_, _01797_, _00350_);
  or (_01912_, _01846_, _26087_);
  and (_01913_, _01912_, _01911_);
  and (_01914_, _01913_, _01910_);
  and (_01915_, _01914_, _01907_);
  nand (_01916_, _01915_, _01900_);
  nor (_01917_, _01853_, _01916_);
  nor (_01918_, _01917_, _01885_);
  and (_01919_, _01649_, _01584_);
  and (_01920_, _01601_, _01584_);
  nor (_01921_, _01920_, _01919_);
  nor (_01922_, _01921_, _01918_);
  not (_01923_, _01602_);
  and (_01924_, _01605_, _01584_);
  not (_01925_, _01924_);
  not (_01926_, _01445_);
  and (_01927_, _01926_, _01414_);
  and (_01928_, _01927_, _01582_);
  not (_01929_, _01617_);
  and (_01930_, _01929_, _01928_);
  and (_01931_, _01929_, _01584_);
  nor (_01932_, _01931_, _01930_);
  nor (_01933_, _01932_, _01918_);
  and (_01934_, _01382_, _01351_);
  not (_01935_, _01934_);
  nor (_01936_, _01935_, _01617_);
  not (_01937_, _01351_);
  and (_01938_, _01382_, _01937_);
  not (_01939_, _01938_);
  or (_01940_, _01939_, _01617_);
  not (_01941_, _01940_);
  nor (_01942_, _01941_, _01936_);
  nor (_01943_, _01942_, _01916_);
  not (_01944_, _01631_);
  and (_01945_, _01944_, _01928_);
  and (_01946_, _01944_, _01584_);
  nor (_01947_, _01946_, _01945_);
  not (_01948_, _01947_);
  and (_01949_, _01948_, _01918_);
  not (_01950_, _01942_);
  and (_01951_, _01944_, _01593_);
  not (_01952_, _01629_);
  and (_01953_, _01952_, _01928_);
  nor (_01954_, _01953_, _01951_);
  nor (_01955_, _01954_, _01916_);
  not (_01956_, _01955_);
  and (_01957_, _01952_, _01584_);
  not (_01958_, _01620_);
  and (_01959_, _01958_, _01584_);
  or (_01960_, _01959_, _01957_);
  and (_01961_, _01960_, _01918_);
  not (_01962_, _01954_);
  and (_01963_, _01952_, _01593_);
  not (_01964_, _01963_);
  nor (_01965_, _01964_, _01916_);
  nor (_01966_, _01965_, _01957_);
  and (_01967_, _01958_, _01928_);
  nor (_01968_, _01967_, _01959_);
  and (_01969_, _01958_, _01593_);
  not (_01970_, _01626_);
  and (_01971_, _01970_, _01593_);
  nor (_01972_, _01971_, _01969_);
  nor (_01973_, _01972_, _01916_);
  not (_01974_, \oc8051_golden_model_1.PSW [3]);
  and (_01975_, _01972_, _01974_);
  nor (_01976_, _01975_, _01973_);
  and (_01977_, _01976_, _01968_);
  and (_01978_, _01967_, \oc8051_golden_model_1.SP [3]);
  or (_01979_, _01978_, _01963_);
  or (_01980_, _01979_, _01977_);
  and (_01981_, _01980_, _01966_);
  or (_01982_, _01981_, _01962_);
  and (_01983_, _01982_, _01947_);
  or (_01984_, _01983_, _01961_);
  and (_01985_, _01984_, _01956_);
  or (_01986_, _01985_, _01950_);
  nor (_01987_, _01986_, _01949_);
  nor (_01988_, _01987_, _01943_);
  not (_01989_, _01932_);
  nor (_01990_, _01989_, _01988_);
  and (_01991_, _01605_, _01593_);
  or (_01992_, _01991_, _01990_);
  nor (_01993_, _01992_, _01933_);
  and (_01994_, _01991_, _01916_);
  or (_01995_, _01994_, _01993_);
  and (_01996_, _01995_, _01925_);
  and (_01997_, _01924_, _01918_);
  or (_01998_, _01997_, _01996_);
  and (_01999_, _01998_, _01923_);
  not (_02000_, _01921_);
  and (_02001_, _01605_, _01928_);
  not (_02002_, _02001_);
  and (_02003_, _01926_, _01382_);
  and (_02004_, _02003_, _01351_);
  not (_02005_, _02004_);
  and (_02006_, _01938_, _01609_);
  and (_02007_, _01934_, _01583_);
  nor (_02008_, _02007_, _02006_);
  and (_02009_, _02008_, _02005_);
  and (_02010_, _01938_, _01927_);
  nor (_02011_, _02010_, _01592_);
  and (_02012_, _02011_, _02009_);
  nor (_02013_, _02012_, _01631_);
  not (_02014_, _02013_);
  and (_02015_, _01659_, _01928_);
  and (_02016_, _01662_, _01610_);
  nor (_02017_, _02016_, _02015_);
  and (_02018_, _01652_, _01610_);
  and (_02019_, _01649_, _01593_);
  nor (_02020_, _02019_, _02018_);
  and (_02021_, _02020_, _02017_);
  and (_02022_, _01580_, _01928_);
  and (_02023_, _01669_, _01584_);
  nor (_02024_, _02023_, _02022_);
  and (_02025_, _01669_, _01928_);
  and (_02026_, _01584_, _01589_);
  nor (_02027_, _02026_, _02025_);
  and (_02028_, _02027_, _02024_);
  and (_02029_, _02028_, _02021_);
  and (_02030_, _01938_, _01590_);
  and (_02031_, _02030_, _01944_);
  and (_02032_, _01934_, _01609_);
  and (_02033_, _02032_, _01944_);
  nor (_02034_, _02033_, _02031_);
  and (_02035_, _01938_, _01583_);
  and (_02036_, _02035_, _01944_);
  nor (_02037_, _02036_, _01969_);
  and (_02038_, _02037_, _02034_);
  and (_02039_, _01665_, _01610_);
  nor (_02040_, _02039_, \oc8051_golden_model_1.PC [0]);
  and (_02041_, _02040_, _02038_);
  and (_02042_, _02041_, _02029_);
  and (_02043_, _02042_, _02014_);
  and (_02044_, _02043_, _02002_);
  nor (_02045_, _02044_, _01298_);
  and (_02046_, _02044_, _01298_);
  nor (_02047_, _02046_, _02045_);
  nor (_02048_, _02001_, _02039_);
  and (_02049_, _02038_, _02048_);
  and (_02050_, _02049_, _02014_);
  and (_02051_, _02050_, _02029_);
  nor (_02052_, _02051_, \oc8051_golden_model_1.PC [0]);
  and (_02053_, _02051_, \oc8051_golden_model_1.PC [0]);
  nor (_02054_, _02053_, _02052_);
  nor (_02055_, _02054_, _02047_);
  nor (_02056_, _02051_, _01770_);
  not (_02057_, _01724_);
  and (_02058_, _02051_, _02057_);
  nor (_02059_, _02058_, _02056_);
  not (_02060_, _01720_);
  nor (_02061_, _02051_, _02060_);
  and (_02062_, _02051_, _01760_);
  nor (_02063_, _02062_, _02061_);
  not (_02064_, _02063_);
  nor (_02065_, _02064_, _02059_);
  and (_02066_, _02065_, _02055_);
  and (_02067_, _02066_, _00354_);
  not (_02068_, _02047_);
  nor (_02069_, _02054_, _02068_);
  and (_02070_, _02069_, _02065_);
  and (_02071_, _02070_, _00374_);
  nor (_02072_, _02071_, _02067_);
  and (_02073_, _02064_, _02059_);
  and (_02074_, _02073_, _02055_);
  and (_02075_, _02074_, _00360_);
  and (_02076_, _02063_, _02059_);
  and (_02077_, _02076_, _02069_);
  and (_02078_, _02077_, _00372_);
  nor (_02079_, _02078_, _02075_);
  and (_02080_, _02079_, _02072_);
  nor (_02081_, _02063_, _02059_);
  and (_02082_, _02054_, _02047_);
  and (_02083_, _02082_, _02081_);
  and (_02084_, _02083_, _00364_);
  and (_02085_, _02081_, _02055_);
  and (_02086_, _02085_, _00400_);
  nor (_02087_, _02086_, _02084_);
  and (_02088_, _02076_, _02055_);
  and (_02089_, _02088_, _00393_);
  and (_02090_, _02054_, _02068_);
  and (_02091_, _02090_, _02065_);
  and (_02092_, _02091_, _00387_);
  nor (_02093_, _02092_, _02089_);
  and (_02094_, _02093_, _02087_);
  and (_02095_, _02094_, _02080_);
  and (_02096_, _02082_, _02073_);
  and (_02097_, _02096_, _00350_);
  and (_02098_, _02073_, _02069_);
  and (_02099_, _02098_, _00378_);
  nor (_02100_, _02099_, _02097_);
  and (_02101_, _02090_, _02073_);
  and (_02102_, _02101_, _00370_);
  and (_02103_, _02090_, _02081_);
  and (_02104_, _02103_, _00398_);
  nor (_02105_, _02104_, _02102_);
  and (_02106_, _02105_, _02100_);
  and (_02107_, _02081_, _02069_);
  and (_02108_, _02107_, _00381_);
  and (_02109_, _02082_, _02065_);
  and (_02110_, _02109_, _00389_);
  nor (_02111_, _02110_, _02108_);
  and (_02112_, _02082_, _02076_);
  and (_02113_, _02112_, _00352_);
  and (_02114_, _02090_, _02076_);
  and (_02115_, _02114_, _00391_);
  nor (_02116_, _02115_, _02113_);
  and (_02117_, _02116_, _02111_);
  and (_02118_, _02117_, _02106_);
  and (_02119_, _02118_, _02095_);
  nor (_02120_, _02119_, _01923_);
  nor (_02121_, _02120_, _02000_);
  not (_02122_, _02121_);
  nor (_02123_, _02122_, _01999_);
  or (_02124_, _02123_, _01922_);
  and (_02125_, _01662_, _01593_);
  and (_02126_, _01662_, _01584_);
  nor (_02127_, _02126_, _02016_);
  not (_02128_, _02127_);
  nor (_02129_, _02128_, _02125_);
  and (_02130_, _01665_, _01584_);
  not (_02131_, _02130_);
  and (_02132_, _01665_, _01593_);
  nor (_02133_, _02132_, _02039_);
  and (_02134_, _02133_, _02131_);
  and (_02135_, _01652_, _01584_);
  not (_02136_, _02135_);
  and (_02137_, _01652_, _01593_);
  nor (_02138_, _02137_, _02018_);
  and (_02139_, _02138_, _02136_);
  and (_02140_, _02139_, _02134_);
  and (_02141_, _02140_, _02129_);
  and (_02142_, _01659_, _01593_);
  not (_02143_, _02142_);
  and (_02144_, _02143_, _02141_);
  nand (_02145_, _02144_, _02124_);
  and (_02146_, _01659_, _01584_);
  nor (_02147_, _02144_, _01916_);
  nor (_02148_, _02147_, _02146_);
  and (_02149_, _02148_, _02145_);
  and (_02150_, _02146_, \oc8051_golden_model_1.SP [3]);
  or (_02151_, _02150_, _02015_);
  nor (_02152_, _02151_, _02149_);
  not (_02153_, _02015_);
  nor (_02154_, _01918_, _02153_);
  or (_02155_, _02154_, _02152_);
  or (_02156_, _02155_, _01597_);
  nand (_02157_, _01916_, _01597_);
  and (_02158_, _02157_, _02156_);
  nand (_02159_, _02158_, _01596_);
  not (_02160_, \oc8051_golden_model_1.SP [3]);
  and (_02161_, _01585_, _02160_);
  nor (_02162_, _02161_, _02022_);
  nand (_02163_, _02162_, _02159_);
  and (_02164_, _01669_, _01593_);
  and (_02165_, _02022_, _01918_);
  nor (_02166_, _02165_, _02164_);
  nand (_02167_, _02166_, _02163_);
  not (_02168_, _02164_);
  nor (_02169_, _02168_, _01916_);
  nor (_02170_, _02169_, _02025_);
  and (_02171_, _02170_, _02167_);
  and (_02172_, _02025_, _01918_);
  or (_02173_, _02172_, _02171_);
  nand (_02174_, _02173_, _01595_);
  and (_02175_, _01916_, _01594_);
  not (_02176_, _02175_);
  and (_02177_, _02176_, _02174_);
  nor (_02178_, _01835_, _26138_);
  nor (_02179_, _01832_, _25590_);
  nor (_02180_, _02179_, _02178_);
  nor (_02181_, _01846_, _26097_);
  nor (_02182_, _01822_, _25877_);
  nor (_02183_, _02182_, _02181_);
  and (_02184_, _02183_, _02180_);
  nor (_02185_, _01818_, _25672_);
  nor (_02186_, _01804_, _25631_);
  nor (_02187_, _02186_, _02185_);
  nor (_02188_, _01841_, _26179_);
  nor (_02189_, _01837_, _26008_);
  nor (_02190_, _02189_, _02188_);
  and (_02191_, _02190_, _02187_);
  and (_02192_, _02191_, _02184_);
  nor (_02193_, _01843_, _25918_);
  nor (_02194_, _01830_, _25754_);
  nor (_02195_, _02194_, _02193_);
  and (_02196_, _01797_, _00460_);
  nor (_02197_, _01808_, _26056_);
  nor (_02198_, _02197_, _02196_);
  and (_02199_, _02198_, _02195_);
  nor (_02200_, _01814_, _25959_);
  nor (_02201_, _01848_, _25836_);
  nor (_02202_, _02201_, _02200_);
  nor (_02204_, _01824_, _25795_);
  nor (_02206_, _01810_, _25713_);
  nor (_02208_, _02206_, _02204_);
  and (_02210_, _02208_, _02202_);
  and (_02212_, _02210_, _02199_);
  and (_02214_, _02212_, _02192_);
  not (_02216_, _02214_);
  and (_02217_, _01924_, _01853_);
  and (_02218_, _02217_, _02216_);
  not (_02219_, _02218_);
  not (_02220_, _01853_);
  nor (_02221_, _02214_, _02220_);
  and (_02222_, _01932_, _01947_);
  not (_02223_, _01959_);
  nor (_02224_, _01957_, _02015_);
  and (_02225_, _02224_, _02223_);
  nor (_02226_, _02022_, _02025_);
  and (_02227_, _02226_, _01921_);
  and (_02228_, _02227_, _02225_);
  and (_02229_, _02228_, _02222_);
  not (_02230_, _02229_);
  and (_02231_, _02230_, _02221_);
  not (_02232_, _02231_);
  nor (_02233_, _01843_, _25903_);
  nor (_02234_, _01830_, _25739_);
  nor (_02235_, _02234_, _02233_);
  and (_02236_, _01797_, _00343_);
  nor (_02237_, _01822_, _25862_);
  nor (_02238_, _02237_, _02236_);
  and (_02239_, _02238_, _02235_);
  nor (_02240_, _01814_, _25944_);
  nor (_02241_, _01824_, _25780_);
  nor (_02242_, _02241_, _02240_);
  nor (_02243_, _01810_, _25698_);
  nor (_02244_, _01832_, _25575_);
  nor (_02245_, _02244_, _02243_);
  and (_02246_, _02245_, _02242_);
  and (_02247_, _02246_, _02239_);
  nor (_02248_, _01835_, _26123_);
  nor (_02249_, _01808_, _26041_);
  nor (_02250_, _02249_, _02248_);
  nor (_02251_, _01848_, _25821_);
  nor (_02252_, _01818_, _25657_);
  nor (_02253_, _02252_, _02251_);
  and (_02254_, _02253_, _02250_);
  nor (_02255_, _01846_, _26082_);
  nor (_02256_, _01837_, _25993_);
  nor (_02257_, _02256_, _02255_);
  nor (_02258_, _01841_, _26164_);
  nor (_02259_, _01804_, _25616_);
  nor (_02260_, _02259_, _02258_);
  and (_02261_, _02260_, _02257_);
  and (_02262_, _02261_, _02254_);
  and (_02263_, _02262_, _02247_);
  not (_02264_, _02263_);
  nor (_02265_, _02164_, _01594_);
  not (_02266_, _02265_);
  nand (_02267_, _01972_, _01954_);
  or (_02268_, _02267_, _01963_);
  or (_02269_, _02268_, _01991_);
  or (_02270_, _02269_, _01950_);
  or (_02271_, _02270_, _02266_);
  and (_02272_, _01592_, _01926_);
  and (_02273_, _01659_, _02272_);
  and (_02274_, _02273_, _01608_);
  nor (_02275_, _02274_, _01597_);
  nand (_02276_, _02275_, _02141_);
  or (_02277_, _02276_, _02271_);
  and (_02278_, _02277_, _02264_);
  and (_02279_, _02096_, _00343_);
  and (_02280_, _02114_, _00336_);
  nor (_02281_, _02280_, _02279_);
  and (_02282_, _02098_, _00306_);
  and (_02283_, _02103_, _00295_);
  nor (_02284_, _02283_, _02282_);
  and (_02285_, _02284_, _02281_);
  and (_02286_, _02091_, _00299_);
  and (_02287_, _02070_, _00319_);
  nor (_02288_, _02287_, _02286_);
  and (_02289_, _02083_, _00303_);
  and (_02290_, _02109_, _00338_);
  nor (_02291_, _02290_, _02289_);
  and (_02292_, _02291_, _02288_);
  and (_02293_, _02292_, _02285_);
  and (_02294_, _02101_, _00327_);
  and (_02295_, _02074_, _00324_);
  nor (_02296_, _02295_, _02294_);
  and (_02297_, _02085_, _00332_);
  and (_02298_, _02077_, _00310_);
  nor (_02299_, _02298_, _02297_);
  and (_02300_, _02299_, _02296_);
  and (_02301_, _02107_, _00316_);
  and (_02302_, _02112_, _00297_);
  nor (_02303_, _02302_, _02301_);
  and (_02304_, _02088_, _00334_);
  and (_02305_, _02066_, _00345_);
  nor (_02306_, _02305_, _02304_);
  and (_02307_, _02306_, _02303_);
  and (_02308_, _02307_, _02300_);
  and (_02309_, _02308_, _02293_);
  nor (_02310_, _02309_, _01923_);
  and (_02311_, _01934_, _01652_);
  nand (_02312_, _01648_, _01577_);
  not (_02313_, _01605_);
  and (_02314_, _01629_, _02313_);
  and (_02315_, _02314_, _01631_);
  and (_02316_, _02315_, _02312_);
  nor (_02317_, _02316_, _01935_);
  nor (_02318_, _02317_, _02311_);
  nor (_02319_, _02318_, _01445_);
  not (_02320_, _02319_);
  and (_02321_, _01934_, _01927_);
  or (_02322_, _01659_, _01580_);
  or (_02323_, _02322_, _01601_);
  and (_02324_, _02323_, _02321_);
  and (_02325_, _01934_, _01445_);
  nor (_02326_, _01599_, _01603_);
  and (_02327_, _02326_, _02325_);
  not (_02328_, _02325_);
  nor (_02329_, _01659_, _01652_);
  nor (_02330_, _02329_, _02328_);
  nor (_02331_, _02330_, _02327_);
  not (_02332_, _02331_);
  nor (_02333_, _02332_, _02324_);
  not (_02334_, \oc8051_golden_model_1.SP [2]);
  nor (_02335_, _01967_, _01585_);
  nor (_02336_, _02335_, _02334_);
  and (_02337_, _01934_, _01590_);
  not (_02338_, _02337_);
  not (_02339_, _01601_);
  nor (_02340_, _01669_, _01580_);
  and (_02341_, _02340_, _02339_);
  nor (_02342_, _02341_, _02338_);
  nor (_02343_, _02342_, _02336_);
  and (_02344_, _02343_, _02333_);
  and (_02345_, _02146_, \oc8051_golden_model_1.SP [2]);
  not (_02346_, _02345_);
  and (_02347_, _01934_, _01669_);
  and (_02348_, _02347_, _01927_);
  nor (_02349_, _01669_, _01952_);
  nor (_02350_, _02349_, _02328_);
  nor (_02351_, _02350_, _02348_);
  and (_02352_, _02351_, _02346_);
  nor (_02353_, _01935_, _01620_);
  not (_02354_, _02353_);
  nor (_02355_, _02312_, _02328_);
  and (_02356_, _02325_, _01601_);
  nor (_02357_, _02356_, _02355_);
  and (_02358_, _02357_, _02354_);
  and (_02359_, _01934_, _01589_);
  nor (_02360_, _01935_, _01626_);
  nor (_02361_, _02360_, _02359_);
  and (_02362_, _02337_, _01659_);
  and (_02363_, _02325_, _01580_);
  nor (_02364_, _02363_, _02362_);
  and (_02365_, _02364_, _02361_);
  and (_02366_, _02365_, _02358_);
  and (_02367_, _02366_, _02352_);
  and (_02368_, _02367_, _02344_);
  and (_02369_, _02368_, _02320_);
  not (_02370_, _02369_);
  nor (_02371_, _02370_, _02310_);
  not (_02372_, _02371_);
  nor (_02373_, _02372_, _02278_);
  and (_02374_, _02373_, _02232_);
  and (_02375_, _02374_, _02219_);
  not (_02376_, \oc8051_golden_model_1.IRAM[0] [7]);
  not (_02377_, _02025_);
  not (_02378_, _01951_);
  or (_02379_, _01808_, _26031_);
  or (_02380_, _01837_, _25983_);
  and (_02381_, _02380_, _02379_);
  or (_02382_, _01822_, _25852_);
  or (_02383_, _01848_, _25811_);
  and (_02384_, _02383_, _02382_);
  and (_02385_, _02384_, _02381_);
  nand (_02386_, _01797_, _00233_);
  or (_02387_, _01841_, _26154_);
  and (_02388_, _02387_, _02386_);
  or (_02389_, _01810_, _25688_);
  or (_02390_, _01818_, _25647_);
  and (_02391_, _02390_, _02389_);
  and (_02392_, _02391_, _02388_);
  and (_02393_, _02392_, _02385_);
  or (_02394_, _01835_, _26113_);
  or (_02395_, _01846_, _26072_);
  and (_02396_, _02395_, _02394_);
  or (_02397_, _01832_, _25563_);
  or (_02398_, _01804_, _25606_);
  and (_02399_, _02398_, _02397_);
  and (_02400_, _02399_, _02396_);
  or (_02401_, _01814_, _25934_);
  or (_02402_, _01843_, _25893_);
  and (_02403_, _02402_, _02401_);
  or (_02404_, _01824_, _25770_);
  or (_02405_, _01830_, _25729_);
  and (_02406_, _02405_, _02404_);
  and (_02407_, _02406_, _02403_);
  and (_02408_, _02407_, _02400_);
  and (_02409_, _02408_, _02393_);
  nor (_02410_, _02409_, _02378_);
  or (_02411_, _02409_, _01964_);
  not (_02412_, _01624_);
  and (_02413_, _01592_, _01583_);
  or (_02414_, _02413_, _01584_);
  and (_02415_, _02414_, _02412_);
  and (_02416_, _01934_, _01414_);
  nor (_02417_, _02416_, _01593_);
  not (_02418_, _02413_);
  nor (_02419_, _02035_, _02010_);
  and (_02420_, _02419_, _02418_);
  and (_02421_, _02420_, _02417_);
  nor (_02422_, _02421_, _01626_);
  nor (_02423_, _02422_, _02415_);
  not (_02424_, _01971_);
  nor (_02425_, _02409_, _02424_);
  or (_02426_, _02425_, _02423_);
  and (_02427_, _02417_, _02418_);
  nor (_02428_, _02427_, _01620_);
  not (_02429_, _02428_);
  and (_02430_, _01970_, _01584_);
  not (_02431_, _02430_);
  and (_02432_, _02010_, _01958_);
  and (_02433_, _02035_, _01958_);
  nor (_02434_, _02433_, _02432_);
  and (_02435_, _02434_, _02431_);
  and (_02436_, _02435_, _02429_);
  nand (_02437_, _02436_, _02426_);
  not (_02438_, _01969_);
  or (_02439_, _02409_, _02438_);
  nand (_02440_, _02439_, _02437_);
  not (_02441_, \oc8051_golden_model_1.SP [0]);
  and (_02442_, _01967_, _02441_);
  or (_02443_, _02442_, _01963_);
  and (_02444_, _02413_, _01952_);
  not (_02445_, _02416_);
  and (_02446_, _02419_, _02445_);
  nor (_02447_, _02446_, _01629_);
  or (_02448_, _02447_, _02444_);
  nor (_02449_, _02448_, _02443_);
  and (_02450_, _01853_, _01916_);
  or (_02451_, _02450_, _02223_);
  and (_02452_, _02451_, _02449_);
  nand (_02453_, _02452_, _02440_);
  nand (_02454_, _02453_, _02411_);
  nor (_02455_, _01957_, _01953_);
  nand (_02456_, _02455_, _02454_);
  not (_02457_, _01953_);
  nor (_02458_, _02409_, _02457_);
  and (_02459_, _02450_, _01957_);
  nor (_02460_, _02459_, _02458_);
  and (_02461_, _02460_, _02456_);
  nor (_02462_, _02421_, _01631_);
  nor (_02463_, _02462_, _02461_);
  or (_02464_, _02463_, _02410_);
  and (_02465_, _02464_, _01947_);
  and (_02466_, _02450_, _01948_);
  or (_02467_, _02466_, _02465_);
  and (_02468_, _02409_, _01950_);
  and (_02469_, _02413_, _01929_);
  nor (_02470_, _02469_, _01989_);
  not (_02471_, _02470_);
  nor (_02472_, _02471_, _02468_);
  and (_02473_, _02472_, _02467_);
  and (_02474_, _02450_, _01989_);
  nor (_02475_, _02474_, _02473_);
  nor (_02476_, _02421_, _02313_);
  nor (_02477_, _02476_, _02475_);
  not (_02478_, _02409_);
  and (_02479_, _02478_, _01991_);
  or (_02480_, _02479_, _02477_);
  and (_02481_, _02480_, _01925_);
  and (_02482_, _02450_, _01924_);
  nor (_02483_, _02482_, _02481_);
  nor (_02484_, _02421_, _02339_);
  nor (_02485_, _02484_, _02483_);
  and (_02486_, _02112_, _00187_);
  and (_02487_, _02091_, _00235_);
  nor (_02488_, _02487_, _02486_);
  and (_02489_, _02098_, _00210_);
  and (_02490_, _02109_, _00226_);
  nor (_02491_, _02490_, _02489_);
  and (_02492_, _02491_, _02488_);
  and (_02493_, _02077_, _00214_);
  and (_02494_, _02114_, _00229_);
  nor (_02495_, _02494_, _02493_);
  and (_02496_, _02101_, _00198_);
  and (_02497_, _02074_, _00193_);
  nor (_02498_, _02497_, _02496_);
  and (_02499_, _02498_, _02495_);
  and (_02500_, _02499_, _02492_);
  and (_02501_, _02107_, _00200_);
  and (_02502_, _02085_, _00185_);
  nor (_02503_, _02502_, _02501_);
  and (_02504_, _02066_, _00189_);
  and (_02505_, _02070_, _00204_);
  nor (_02506_, _02505_, _02504_);
  and (_02507_, _02506_, _02503_);
  and (_02508_, _02096_, _00233_);
  and (_02509_, _02088_, _00223_);
  nor (_02510_, _02509_, _02508_);
  and (_02511_, _02083_, _00195_);
  and (_02512_, _02103_, _00220_);
  nor (_02513_, _02512_, _02511_);
  and (_02514_, _02513_, _02510_);
  and (_02515_, _02514_, _02507_);
  and (_02516_, _02515_, _02500_);
  nor (_02517_, _02516_, _01923_);
  or (_02518_, _02517_, _02485_);
  not (_02519_, _01920_);
  nor (_02520_, _02450_, _02519_);
  and (_02521_, _02414_, _01649_);
  nor (_02522_, _02521_, _02520_);
  and (_02523_, _02522_, _02518_);
  and (_02524_, _02450_, _01919_);
  nor (_02525_, _02524_, _02523_);
  not (_02526_, _01652_);
  and (_02527_, _02420_, _02445_);
  nor (_02528_, _02527_, _02526_);
  nor (_02529_, _02528_, _02525_);
  nor (_02530_, _02478_, _02139_);
  not (_02531_, _01665_);
  nor (_02532_, _02527_, _02531_);
  nor (_02533_, _02532_, _02530_);
  and (_02534_, _02533_, _02529_);
  nor (_02535_, _02478_, _02134_);
  not (_02536_, _01662_);
  nor (_02537_, _02527_, _02536_);
  nor (_02538_, _02537_, _02535_);
  and (_02539_, _02538_, _02534_);
  nor (_02540_, _02478_, _02129_);
  not (_02541_, _01659_);
  nor (_02542_, _02421_, _02541_);
  nor (_02543_, _02542_, _02540_);
  and (_02544_, _02543_, _02539_);
  nor (_02545_, _02409_, _02143_);
  nor (_02546_, _02545_, _02544_);
  and (_02547_, _02146_, _02441_);
  nor (_02548_, _02547_, _02546_);
  nor (_02549_, _02450_, _02153_);
  not (_02550_, _01580_);
  nor (_02551_, _02421_, _02550_);
  nor (_02552_, _02551_, _02549_);
  and (_02553_, _02552_, _02548_);
  and (_02554_, _02478_, _01597_);
  nor (_02555_, _02554_, _02553_);
  and (_02556_, _01585_, _02441_);
  nor (_02557_, _02556_, _02555_);
  not (_02558_, _02022_);
  nor (_02559_, _02450_, _02558_);
  not (_02560_, _01669_);
  nor (_02561_, _02421_, _02560_);
  nor (_02562_, _02561_, _02559_);
  and (_02563_, _02562_, _02557_);
  nor (_02564_, _02409_, _02168_);
  or (_02565_, _02564_, _02563_);
  and (_02566_, _02565_, _02377_);
  and (_02567_, _02450_, _02025_);
  nor (_02568_, _02567_, _02566_);
  not (_02569_, _01589_);
  nor (_02570_, _02421_, _02569_);
  or (_02571_, _02570_, _02568_);
  nor (_02572_, _02409_, _01595_);
  not (_02573_, _02572_);
  nand (_02574_, _02573_, _02571_);
  or (_02575_, _02574_, _02376_);
  nor (_02576_, _01832_, _25585_);
  nor (_02577_, _01818_, _25667_);
  nor (_02578_, _02577_, _02576_);
  nor (_02579_, _01846_, _26092_);
  nor (_02580_, _01822_, _25872_);
  nor (_02581_, _02580_, _02579_);
  and (_02582_, _02581_, _02578_);
  nor (_02583_, _01808_, _26051_);
  nor (_02584_, _01843_, _25913_);
  nor (_02585_, _02584_, _02583_);
  nor (_02586_, _01824_, _25790_);
  nor (_02587_, _01810_, _25708_);
  nor (_02588_, _02587_, _02586_);
  and (_02589_, _02588_, _02585_);
  and (_02590_, _02589_, _02582_);
  and (_02591_, _01797_, _00442_);
  nor (_02592_, _01841_, _26174_);
  nor (_02593_, _02592_, _02591_);
  nor (_02594_, _01835_, _26133_);
  nor (_02595_, _01814_, _25954_);
  nor (_02596_, _02595_, _02594_);
  and (_02597_, _02596_, _02593_);
  nor (_02598_, _01837_, _26003_);
  nor (_02599_, _01804_, _25626_);
  nor (_02600_, _02599_, _02598_);
  nor (_02601_, _01848_, _25831_);
  nor (_02602_, _01830_, _25749_);
  nor (_02603_, _02602_, _02601_);
  and (_02604_, _02603_, _02600_);
  and (_02605_, _02604_, _02597_);
  and (_02606_, _02605_, _02590_);
  not (_02607_, _02606_);
  and (_02608_, _02607_, _02217_);
  not (_02609_, _02608_);
  nor (_02610_, _02606_, _02220_);
  and (_02611_, _02610_, _02230_);
  not (_02612_, _02611_);
  and (_02613_, _01797_, _00240_);
  nor (_02614_, _01824_, _25775_);
  nor (_02615_, _02614_, _02613_);
  nor (_02616_, _01841_, _26159_);
  nor (_02617_, _01843_, _25898_);
  nor (_02618_, _02617_, _02616_);
  and (_02619_, _02618_, _02615_);
  nor (_02620_, _01804_, _25611_);
  nor (_02621_, _01818_, _25652_);
  nor (_02622_, _02621_, _02620_);
  nor (_02623_, _01808_, _26036_);
  nor (_02624_, _01810_, _25693_);
  nor (_02625_, _02624_, _02623_);
  and (_02626_, _02625_, _02622_);
  and (_02627_, _02626_, _02619_);
  nor (_02628_, _01835_, _26118_);
  nor (_02629_, _01846_, _26077_);
  nor (_02630_, _02629_, _02628_);
  nor (_02631_, _01814_, _25939_);
  nor (_02632_, _01848_, _25816_);
  nor (_02633_, _02632_, _02631_);
  and (_02634_, _02633_, _02630_);
  nor (_02635_, _01837_, _25988_);
  nor (_02636_, _01822_, _25857_);
  nor (_02637_, _02636_, _02635_);
  nor (_02638_, _01830_, _25734_);
  nor (_02639_, _01832_, _25568_);
  nor (_02640_, _02639_, _02638_);
  and (_02641_, _02640_, _02637_);
  and (_02642_, _02641_, _02634_);
  and (_02643_, _02642_, _02627_);
  not (_02644_, _02643_);
  and (_02645_, _02644_, _02277_);
  and (_02646_, _02083_, _00247_);
  and (_02647_, _02112_, _00278_);
  nor (_02648_, _02647_, _02646_);
  and (_02649_, _02077_, _00260_);
  and (_02650_, _02091_, _00269_);
  nor (_02651_, _02650_, _02649_);
  and (_02652_, _02651_, _02648_);
  and (_02653_, _02101_, _00245_);
  and (_02654_, _02098_, _00286_);
  nor (_02655_, _02654_, _02653_);
  and (_02656_, _02096_, _00240_);
  and (_02657_, _02109_, _00271_);
  nor (_02658_, _02657_, _02656_);
  and (_02659_, _02658_, _02655_);
  and (_02660_, _02659_, _02652_);
  and (_02661_, _02114_, _00264_);
  and (_02662_, _02088_, _00256_);
  nor (_02663_, _02662_, _02661_);
  and (_02664_, _02107_, _00282_);
  and (_02665_, _02066_, _00288_);
  nor (_02666_, _02665_, _02664_);
  and (_02667_, _02666_, _02663_);
  and (_02668_, _02074_, _00249_);
  and (_02669_, _02070_, _00290_);
  nor (_02670_, _02669_, _02668_);
  and (_02671_, _02103_, _00280_);
  and (_02672_, _02085_, _00242_);
  nor (_02673_, _02672_, _02671_);
  and (_02674_, _02673_, _02670_);
  and (_02675_, _02674_, _02667_);
  and (_02676_, _02675_, _02660_);
  nor (_02677_, _02676_, _01923_);
  and (_02678_, _02325_, _01970_);
  not (_02679_, _02678_);
  and (_02680_, _02325_, _01589_);
  and (_02681_, _02035_, _01659_);
  nor (_02682_, _02681_, _02680_);
  and (_02683_, _02682_, _02679_);
  nor (_02684_, _02363_, _02355_);
  and (_02685_, _02035_, _01580_);
  nor (_02686_, _02685_, _02356_);
  and (_02687_, _02686_, _02684_);
  and (_02688_, _02687_, _02683_);
  not (_02689_, _02006_);
  nor (_02690_, _01659_, _01601_);
  and (_02691_, _02690_, _02313_);
  nor (_02692_, _02691_, _02689_);
  nor (_02693_, _02692_, _02332_);
  and (_02694_, _02693_, _02688_);
  not (_02695_, _02035_);
  nor (_02696_, _01605_, _01601_);
  nor (_02697_, _02696_, _02695_);
  not (_02698_, _02697_);
  and (_02699_, _02325_, _01958_);
  and (_02700_, _02035_, _01669_);
  nor (_02701_, _02700_, _02699_);
  and (_02702_, _02701_, _02698_);
  nor (_02703_, _02006_, _02035_);
  nor (_02704_, _02703_, _02536_);
  nor (_02705_, _02704_, _02350_);
  nor (_02706_, _02703_, _02526_);
  nor (_02707_, _02340_, _02689_);
  nor (_02708_, _02707_, _02706_);
  and (_02709_, _02708_, _02705_);
  and (_02710_, _02709_, _02702_);
  nor (_02711_, _01665_, _01589_);
  and (_02712_, _01620_, _01629_);
  and (_02713_, _01626_, _01631_);
  and (_02714_, _02713_, _02712_);
  and (_02715_, _02714_, _02711_);
  nor (_02716_, _02715_, _02703_);
  not (_02717_, \oc8051_golden_model_1.SP [1]);
  not (_02718_, _02146_);
  and (_02719_, _02335_, _02718_);
  nor (_02720_, _02719_, _02717_);
  nor (_02721_, _02720_, _02716_);
  and (_02722_, _02721_, _02710_);
  and (_02723_, _02722_, _02694_);
  not (_02724_, _02723_);
  nor (_02725_, _02724_, _02677_);
  not (_02726_, _02725_);
  nor (_02727_, _02726_, _02645_);
  and (_02728_, _02727_, _02612_);
  and (_02729_, _02728_, _02609_);
  not (_02730_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_02731_, _02573_, _02571_);
  or (_02732_, _02731_, _02730_);
  and (_02733_, _02732_, _02729_);
  nand (_02734_, _02733_, _02575_);
  not (_02735_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_02736_, _02731_, _02735_);
  not (_02737_, _02729_);
  not (_02738_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_02739_, _02574_, _02738_);
  and (_02740_, _02739_, _02737_);
  nand (_02741_, _02740_, _02736_);
  nand (_02742_, _02741_, _02734_);
  nand (_02743_, _02742_, _02375_);
  not (_02744_, _02375_);
  not (_02745_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_02746_, _02731_, _02745_);
  not (_02747_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_02748_, _02574_, _02747_);
  and (_02749_, _02748_, _02737_);
  nand (_02750_, _02749_, _02746_);
  not (_02751_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_02752_, _02574_, _02751_);
  not (_02753_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_02754_, _02731_, _02753_);
  and (_02755_, _02754_, _02729_);
  nand (_02756_, _02755_, _02752_);
  nand (_02757_, _02756_, _02750_);
  nand (_02758_, _02757_, _02744_);
  nand (_02759_, _02758_, _02743_);
  nand (_02760_, _02759_, _02177_);
  not (_02761_, _02177_);
  nand (_02762_, _02574_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand (_02763_, _02731_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_02764_, _02763_, _02737_);
  nand (_02765_, _02764_, _02762_);
  nand (_02766_, _02731_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_02767_, _02574_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_02768_, _02767_, _02729_);
  nand (_02769_, _02768_, _02766_);
  nand (_02770_, _02769_, _02765_);
  nand (_02772_, _02770_, _02375_);
  nand (_02773_, _02574_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_02774_, _02731_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_02776_, _02774_, _02737_);
  nand (_02777_, _02776_, _02773_);
  nand (_02778_, _02731_, \oc8051_golden_model_1.IRAM[12] [7]);
  nand (_02779_, _02574_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_02780_, _02779_, _02729_);
  nand (_02781_, _02780_, _02778_);
  nand (_02782_, _02781_, _02777_);
  nand (_02783_, _02782_, _02744_);
  nand (_02784_, _02783_, _02772_);
  nand (_02785_, _02784_, _02761_);
  nand (_02786_, _02785_, _02760_);
  nand (_02787_, _02786_, _01585_);
  and (_02788_, _02272_, _01580_);
  not (_02789_, _01312_);
  and (_02790_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_02791_, _02790_, _02789_);
  and (_02792_, _02791_, \oc8051_golden_model_1.PC [6]);
  and (_02793_, _02792_, \oc8051_golden_model_1.PC [7]);
  and (_02794_, _02793_, \oc8051_golden_model_1.PC [8]);
  and (_02795_, _02794_, \oc8051_golden_model_1.PC [9]);
  and (_02796_, _02795_, \oc8051_golden_model_1.PC [10]);
  and (_02797_, _02796_, \oc8051_golden_model_1.PC [11]);
  and (_02798_, _02797_, \oc8051_golden_model_1.PC [12]);
  and (_02799_, _02798_, \oc8051_golden_model_1.PC [13]);
  and (_02800_, _02799_, \oc8051_golden_model_1.PC [14]);
  or (_02801_, _02800_, \oc8051_golden_model_1.PC [15]);
  nand (_02802_, _02800_, \oc8051_golden_model_1.PC [15]);
  and (_02803_, _02802_, _02801_);
  and (_02804_, _01609_, _01592_);
  and (_02805_, _02804_, _01580_);
  and (_02806_, _02003_, _01608_);
  nor (_02807_, _02806_, _02006_);
  nor (_02808_, _02807_, _02550_);
  nor (_02809_, _02808_, _02805_);
  and (_02810_, _02321_, _01580_);
  nor (_02811_, _02685_, _02810_);
  not (_02812_, _02363_);
  and (_02813_, _02413_, _01580_);
  and (_02814_, _02010_, _01580_);
  nor (_02815_, _02814_, _02813_);
  and (_02816_, _02815_, _02812_);
  and (_02817_, _02816_, _02811_);
  and (_02818_, _02817_, _02809_);
  or (_02819_, _02818_, _02803_);
  nor (_02820_, _02706_, _02311_);
  and (_02821_, _02030_, _01652_);
  not (_02822_, _02821_);
  and (_02823_, _02413_, _01652_);
  and (_02824_, _02010_, _01652_);
  nor (_02825_, _02824_, _02823_);
  and (_02826_, _02804_, _01652_);
  not (_02827_, _02826_);
  and (_02828_, _02827_, _02825_);
  and (_02829_, _02828_, _02822_);
  and (_02830_, _02829_, _02820_);
  or (_02831_, _02830_, _02803_);
  and (_02832_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_02833_, _02832_, \oc8051_golden_model_1.PC [10]);
  and (_02834_, \oc8051_golden_model_1.PC [7], \oc8051_golden_model_1.PC [6]);
  and (_02835_, _02834_, _02790_);
  and (_02836_, _02835_, _01718_);
  and (_02837_, _02836_, _02833_);
  and (_02838_, _02837_, \oc8051_golden_model_1.PC [11]);
  and (_02839_, _02838_, \oc8051_golden_model_1.PC [12]);
  and (_02840_, _02839_, \oc8051_golden_model_1.PC [13]);
  and (_02841_, _02840_, \oc8051_golden_model_1.PC [14]);
  nor (_02842_, _02841_, \oc8051_golden_model_1.PC [15]);
  and (_02843_, _02836_, \oc8051_golden_model_1.PC [8]);
  and (_02844_, _02843_, \oc8051_golden_model_1.PC [9]);
  and (_02845_, _02844_, \oc8051_golden_model_1.PC [10]);
  and (_02846_, _02845_, \oc8051_golden_model_1.PC [11]);
  and (_02847_, _02846_, \oc8051_golden_model_1.PC [12]);
  and (_02848_, _02847_, \oc8051_golden_model_1.PC [13]);
  and (_02849_, _02848_, \oc8051_golden_model_1.PC [14]);
  and (_02850_, _02849_, \oc8051_golden_model_1.PC [15]);
  nor (_02851_, _02850_, _02842_);
  and (_02852_, _01592_, _01927_);
  and (_02853_, _02852_, _01649_);
  and (_02854_, _02853_, _02851_);
  not (_02855_, _02851_);
  not (_02856_, _01649_);
  and (_02857_, _01592_, _01445_);
  nor (_02858_, _02857_, _01382_);
  nor (_02859_, _02858_, _02856_);
  nand (_02860_, _02859_, _02855_);
  and (_02861_, _01329_, \oc8051_golden_model_1.PC [2]);
  and (_02862_, _02861_, \oc8051_golden_model_1.PC [3]);
  and (_02863_, _02862_, _02835_);
  and (_02864_, _02863_, _02833_);
  and (_02865_, _02864_, \oc8051_golden_model_1.PC [11]);
  and (_02866_, _02865_, \oc8051_golden_model_1.PC [12]);
  and (_02867_, _02866_, \oc8051_golden_model_1.PC [13]);
  and (_02868_, _02867_, \oc8051_golden_model_1.PC [14]);
  nor (_02869_, _02868_, \oc8051_golden_model_1.PC [15]);
  and (_02870_, _02863_, \oc8051_golden_model_1.PC [8]);
  and (_02871_, _02870_, \oc8051_golden_model_1.PC [9]);
  and (_02872_, _02871_, \oc8051_golden_model_1.PC [10]);
  and (_02873_, _02872_, \oc8051_golden_model_1.PC [11]);
  and (_02874_, _02873_, \oc8051_golden_model_1.PC [12]);
  and (_02875_, _02874_, \oc8051_golden_model_1.PC [13]);
  and (_02876_, _02875_, \oc8051_golden_model_1.PC [14]);
  and (_02877_, _02876_, \oc8051_golden_model_1.PC [15]);
  nor (_02878_, _02877_, _02869_);
  and (_02879_, _02878_, _01602_);
  and (_02880_, _01944_, _01610_);
  not (_02881_, _02880_);
  nor (_02882_, _02409_, \oc8051_golden_model_1.ACC [0]);
  and (_02883_, _02409_, \oc8051_golden_model_1.ACC [0]);
  nor (_02884_, _02883_, _02882_);
  nor (_02885_, _02643_, \oc8051_golden_model_1.ACC [1]);
  and (_02886_, _02643_, \oc8051_golden_model_1.ACC [1]);
  nor (_02887_, _02886_, _02885_);
  and (_02888_, _02887_, _02884_);
  and (_02889_, _01916_, _01732_);
  nor (_02890_, _01916_, _01732_);
  nor (_02891_, _02890_, _02889_);
  nor (_02892_, _02263_, \oc8051_golden_model_1.ACC [2]);
  and (_02893_, _02263_, \oc8051_golden_model_1.ACC [2]);
  nor (_02894_, _02893_, _02892_);
  and (_02895_, _02894_, _02891_);
  and (_02896_, _02895_, _02888_);
  nor (_02897_, _01884_, \oc8051_golden_model_1.ACC [6]);
  and (_02898_, _01884_, \oc8051_golden_model_1.ACC [6]);
  nor (_02899_, _02898_, _02897_);
  nor (_02900_, _01853_, \oc8051_golden_model_1.ACC [7]);
  and (_02901_, _01853_, \oc8051_golden_model_1.ACC [7]);
  nor (_02902_, _02901_, _02900_);
  and (_02903_, _02902_, _02899_);
  nor (_02904_, _02606_, \oc8051_golden_model_1.ACC [4]);
  and (_02905_, _02606_, \oc8051_golden_model_1.ACC [4]);
  nor (_02906_, _02905_, _02904_);
  nor (_02907_, _02214_, \oc8051_golden_model_1.ACC [5]);
  and (_02908_, _02214_, \oc8051_golden_model_1.ACC [5]);
  nor (_02909_, _02908_, _02907_);
  and (_02910_, _02909_, _02906_);
  and (_02911_, _02910_, _02903_);
  and (_02912_, _02911_, _02896_);
  and (_02913_, _02096_, _00063_);
  and (_02914_, _02083_, _00027_);
  nor (_02915_, _02914_, _02913_);
  and (_02916_, _02077_, _00043_);
  and (_02917_, _02066_, _00067_);
  nor (_02918_, _02917_, _02916_);
  and (_02919_, _02918_, _02915_);
  and (_02920_, _02098_, _00019_);
  and (_02921_, _02074_, _00014_);
  nor (_02922_, _02921_, _02920_);
  and (_02923_, _02101_, _00022_);
  and (_02924_, _02085_, _00030_);
  nor (_02925_, _02924_, _02923_);
  and (_02926_, _02925_, _02922_);
  and (_02927_, _02926_, _02919_);
  and (_02928_, _02088_, _00055_);
  and (_02929_, _02109_, _00049_);
  nor (_02930_, _02929_, _02928_);
  and (_02931_, _02112_, _29605_);
  and (_02932_, _02114_, _00040_);
  nor (_02933_, _02932_, _02931_);
  and (_02934_, _02933_, _02930_);
  and (_02935_, _02107_, _29623_);
  and (_02936_, _02103_, _00007_);
  nor (_02937_, _02936_, _02935_);
  and (_02938_, _02070_, _00071_);
  and (_02939_, _02091_, _00036_);
  nor (_02940_, _02939_, _02938_);
  and (_02941_, _02940_, _02937_);
  and (_02942_, _02941_, _02934_);
  and (_02943_, _02942_, _02927_);
  nor (_02944_, _02867_, \oc8051_golden_model_1.PC [14]);
  nor (_02945_, _02944_, _02868_);
  not (_02946_, _02945_);
  nor (_02947_, _02946_, _02943_);
  and (_02948_, _02946_, _02943_);
  nor (_02949_, _02948_, _02947_);
  not (_02950_, _02949_);
  not (_02951_, \oc8051_golden_model_1.PC [13]);
  and (_02952_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and (_02953_, _02952_, _02832_);
  and (_02954_, _02863_, _02953_);
  and (_02955_, _02954_, \oc8051_golden_model_1.PC [12]);
  nor (_02956_, _02955_, _02951_);
  and (_02957_, _02955_, _02951_);
  or (_02958_, _02957_, _02956_);
  not (_02959_, _02958_);
  nor (_02960_, _02959_, _02943_);
  and (_02961_, _02959_, _02943_);
  not (_02962_, _02943_);
  nor (_02963_, _02865_, \oc8051_golden_model_1.PC [12]);
  nor (_02964_, _02963_, _02866_);
  and (_02965_, _02964_, _02962_);
  nor (_02966_, _02871_, \oc8051_golden_model_1.PC [10]);
  nor (_02967_, _02966_, _02864_);
  not (_02968_, _02967_);
  nor (_02969_, _02968_, _02943_);
  not (_02970_, _02969_);
  not (_02971_, \oc8051_golden_model_1.PC [11]);
  nor (_02972_, _02864_, _02971_);
  and (_02973_, _02864_, _02971_);
  or (_02974_, _02973_, _02972_);
  not (_02975_, _02974_);
  nor (_02976_, _02975_, _02943_);
  and (_02977_, _02975_, _02943_);
  nor (_02978_, _02977_, _02976_);
  and (_02979_, _02968_, _02943_);
  nor (_02980_, _02979_, _02969_);
  and (_02981_, _02980_, _02978_);
  nor (_02982_, _02870_, \oc8051_golden_model_1.PC [9]);
  nor (_02983_, _02982_, _02871_);
  not (_02984_, _02983_);
  nor (_02985_, _02984_, _02943_);
  and (_02986_, _02984_, _02943_);
  nor (_02987_, _02986_, _02985_);
  and (_02988_, _02790_, \oc8051_golden_model_1.PC [6]);
  and (_02989_, _02862_, _02988_);
  nor (_02990_, _02989_, \oc8051_golden_model_1.PC [7]);
  nor (_02991_, _02990_, _02863_);
  not (_02992_, _02991_);
  nor (_02993_, _02992_, _02943_);
  and (_02994_, _02992_, _02943_);
  and (_02995_, _02083_, _00530_);
  and (_02996_, _02112_, _00565_);
  nor (_02997_, _02996_, _02995_);
  and (_02998_, _02077_, _00544_);
  and (_02999_, _02091_, _00552_);
  nor (_03000_, _02999_, _02998_);
  and (_03001_, _03000_, _02997_);
  and (_03002_, _02096_, _00522_);
  and (_03003_, _02109_, _00554_);
  nor (_03004_, _03003_, _03002_);
  and (_03005_, _02098_, _00541_);
  and (_03006_, _02074_, _00532_);
  nor (_03007_, _03006_, _03005_);
  and (_03008_, _03007_, _03004_);
  and (_03009_, _03008_, _03001_);
  and (_03010_, _02114_, _00556_);
  and (_03011_, _02088_, _00558_);
  nor (_03012_, _03011_, _03010_);
  and (_03013_, _02107_, _00546_);
  and (_03014_, _02066_, _00563_);
  nor (_03015_, _03014_, _03013_);
  and (_03016_, _03015_, _03012_);
  and (_03017_, _02101_, _00537_);
  and (_03018_, _02070_, _00539_);
  nor (_03019_, _03018_, _03017_);
  and (_03020_, _02103_, _00518_);
  and (_03021_, _02085_, _00526_);
  nor (_03022_, _03021_, _03020_);
  and (_03023_, _03022_, _03019_);
  and (_03024_, _03023_, _03016_);
  and (_03025_, _03024_, _03009_);
  and (_03026_, _02862_, _02790_);
  nor (_03027_, _03026_, \oc8051_golden_model_1.PC [6]);
  nor (_03028_, _03027_, _02989_);
  not (_03029_, _03028_);
  nor (_03030_, _03029_, _03025_);
  and (_03031_, _03029_, _03025_);
  nor (_03032_, _03031_, _03030_);
  not (_03033_, _03032_);
  and (_03034_, _02096_, _00460_);
  and (_03035_, _02103_, _00500_);
  nor (_03036_, _03035_, _03034_);
  and (_03037_, _02107_, _00502_);
  and (_03038_, _02109_, _00493_);
  nor (_03039_, _03038_, _03037_);
  and (_03040_, _03039_, _03036_);
  and (_03041_, _02112_, _00498_);
  and (_03042_, _02088_, _00482_);
  nor (_03043_, _03042_, _03041_);
  and (_03044_, _02101_, _00470_);
  and (_03045_, _02074_, _00476_);
  nor (_03046_, _03045_, _03044_);
  and (_03047_, _03046_, _03043_);
  and (_03048_, _03047_, _03040_);
  and (_03049_, _02114_, _00487_);
  and (_03050_, _02070_, _00510_);
  nor (_03051_, _03050_, _03049_);
  and (_03052_, _02066_, _00508_);
  and (_03053_, _02091_, _00491_);
  nor (_03054_, _03053_, _03052_);
  and (_03055_, _03054_, _03051_);
  and (_03056_, _02098_, _00506_);
  and (_03057_, _02077_, _00485_);
  nor (_03058_, _03057_, _03056_);
  and (_03059_, _02083_, _00474_);
  and (_03060_, _02085_, _00464_);
  nor (_03061_, _03060_, _03059_);
  and (_03062_, _03061_, _03058_);
  and (_03063_, _03062_, _03055_);
  and (_03064_, _03063_, _03048_);
  and (_03065_, _02862_, \oc8051_golden_model_1.PC [4]);
  nor (_03066_, _03065_, \oc8051_golden_model_1.PC [5]);
  nor (_03067_, _03066_, _03026_);
  not (_03068_, _03067_);
  nor (_03069_, _03068_, _03064_);
  and (_03070_, _03068_, _03064_);
  and (_03071_, _02109_, _00444_);
  and (_03072_, _02070_, _00422_);
  nor (_03073_, _03072_, _03071_);
  and (_03074_, _02088_, _00446_);
  and (_03075_, _02091_, _00453_);
  nor (_03076_, _03075_, _03074_);
  and (_03077_, _03076_, _03073_);
  and (_03078_, _02096_, _00442_);
  and (_03079_, _02098_, _00430_);
  nor (_03080_, _03079_, _03078_);
  and (_03081_, _02074_, _00436_);
  and (_03082_, _02107_, _00424_);
  nor (_03083_, _03082_, _03081_);
  and (_03084_, _03083_, _03080_);
  and (_03085_, _03084_, _03077_);
  and (_03086_, _02103_, _00410_);
  and (_03087_, _02114_, _00449_);
  nor (_03088_, _03087_, _03086_);
  and (_03089_, _02083_, _00418_);
  and (_03090_, _02066_, _00407_);
  nor (_03091_, _03090_, _03089_);
  and (_03092_, _03091_, _03088_);
  and (_03093_, _02085_, _00455_);
  and (_03094_, _02112_, _00405_);
  nor (_03095_, _03094_, _03093_);
  and (_03096_, _02101_, _00438_);
  and (_03097_, _02077_, _00427_);
  nor (_03098_, _03097_, _03096_);
  and (_03099_, _03098_, _03095_);
  and (_03100_, _03099_, _03092_);
  and (_03101_, _03100_, _03085_);
  nor (_03102_, _02862_, \oc8051_golden_model_1.PC [4]);
  nor (_03103_, _03102_, _03065_);
  not (_03104_, _03103_);
  nor (_03105_, _03104_, _03101_);
  nor (_03106_, _02861_, \oc8051_golden_model_1.PC [3]);
  nor (_03107_, _03106_, _02862_);
  not (_03108_, _03107_);
  nor (_03109_, _03108_, _02119_);
  and (_03110_, _03108_, _02119_);
  nor (_03111_, _01329_, \oc8051_golden_model_1.PC [2]);
  nor (_03112_, _03111_, _02861_);
  not (_03113_, _03112_);
  nor (_03114_, _03113_, _02309_);
  not (_03115_, _01690_);
  nor (_03116_, _02676_, _03115_);
  nor (_03117_, _02516_, \oc8051_golden_model_1.PC [0]);
  and (_03118_, _02676_, _03115_);
  nor (_03119_, _03118_, _03116_);
  and (_03120_, _03119_, _03117_);
  nor (_03121_, _03120_, _03116_);
  and (_03122_, _03113_, _02309_);
  nor (_03123_, _03122_, _03114_);
  not (_03124_, _03123_);
  nor (_03125_, _03124_, _03121_);
  nor (_03126_, _03125_, _03114_);
  nor (_03127_, _03126_, _03110_);
  nor (_03128_, _03127_, _03109_);
  and (_03129_, _03104_, _03101_);
  nor (_03130_, _03129_, _03105_);
  not (_03131_, _03130_);
  nor (_03132_, _03131_, _03128_);
  nor (_03133_, _03132_, _03105_);
  nor (_03134_, _03133_, _03070_);
  nor (_03135_, _03134_, _03069_);
  nor (_03136_, _03135_, _03033_);
  nor (_03137_, _03136_, _03030_);
  nor (_03138_, _03137_, _02994_);
  or (_03139_, _03138_, _02993_);
  nor (_03140_, _02863_, \oc8051_golden_model_1.PC [8]);
  nor (_03141_, _03140_, _02870_);
  not (_03142_, _03141_);
  nor (_03143_, _03142_, _02943_);
  and (_03144_, _03142_, _02943_);
  nor (_03145_, _03144_, _03143_);
  and (_03146_, _03145_, _03139_);
  and (_03147_, _03146_, _02987_);
  and (_03148_, _03147_, _02981_);
  nor (_03149_, _03143_, _02985_);
  not (_03150_, _03149_);
  and (_03151_, _03150_, _02981_);
  or (_03152_, _03151_, _02976_);
  nor (_03154_, _03152_, _03148_);
  and (_03155_, _03154_, _02970_);
  not (_03156_, _03155_);
  nor (_03157_, _02964_, _02962_);
  nor (_03158_, _03157_, _02965_);
  and (_03159_, _03158_, _03156_);
  nor (_03161_, _03159_, _02965_);
  nor (_03162_, _03161_, _02961_);
  nor (_03163_, _03162_, _02960_);
  nor (_03165_, _03163_, _02950_);
  nor (_03166_, _03165_, _02947_);
  not (_03168_, _02878_);
  and (_03169_, _02943_, _03168_);
  nor (_03171_, _02943_, _03168_);
  nor (_03172_, _03171_, _03169_);
  and (_03174_, _03172_, _03166_);
  nor (_03175_, _03172_, _03166_);
  or (_03176_, _03175_, _03174_);
  or (_03178_, _03176_, _02912_);
  and (_03179_, _02852_, _01944_);
  nand (_03181_, _02912_, _03168_);
  and (_03182_, _03181_, _03179_);
  and (_03184_, _03182_, _03178_);
  and (_03185_, _02857_, _01944_);
  not (_03187_, _03185_);
  not (_03188_, _01916_);
  or (_03189_, _02146_, _01585_);
  nor (_03190_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_03192_, _03190_, _02334_);
  nor (_03193_, _03190_, _02334_);
  nor (_03195_, _03193_, _03192_);
  not (_03196_, _03195_);
  and (_03198_, _03196_, _03189_);
  not (_03199_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_03201_, _02574_, _03199_);
  not (_03203_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_03205_, _02731_, _03203_);
  and (_03206_, _03205_, _02729_);
  nand (_03208_, _03206_, _03201_);
  not (_03209_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_03211_, _02731_, _03209_);
  not (_03213_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_03214_, _02574_, _03213_);
  and (_03216_, _03214_, _02737_);
  nand (_03217_, _03216_, _03211_);
  nand (_03219_, _03217_, _03208_);
  nand (_03220_, _03219_, _02375_);
  not (_03222_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_03223_, _02731_, _03222_);
  not (_03225_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_03227_, _02574_, _03225_);
  and (_03229_, _03227_, _02737_);
  nand (_03231_, _03229_, _03223_);
  not (_03233_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_03235_, _02574_, _03233_);
  not (_03237_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_03239_, _02731_, _03237_);
  and (_03241_, _03239_, _02729_);
  nand (_03243_, _03241_, _03235_);
  nand (_03245_, _03243_, _03231_);
  nand (_03246_, _03245_, _02744_);
  nand (_03247_, _03246_, _03220_);
  nand (_03248_, _03247_, _02177_);
  nand (_03249_, _02574_, \oc8051_golden_model_1.IRAM[11] [2]);
  not (_03250_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_03251_, _02574_, _03250_);
  and (_03252_, _03251_, _02737_);
  nand (_03253_, _03252_, _03249_);
  nand (_03254_, _02731_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_03255_, _02574_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_03256_, _03255_, _02729_);
  nand (_03257_, _03256_, _03254_);
  nand (_03258_, _03257_, _03253_);
  nand (_03259_, _03258_, _02375_);
  nand (_03260_, _02574_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_03261_, _02731_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_03262_, _03261_, _02737_);
  nand (_03263_, _03262_, _03260_);
  nand (_03264_, _02731_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_03265_, _02574_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_03266_, _03265_, _02729_);
  nand (_03267_, _03266_, _03264_);
  nand (_03268_, _03267_, _03263_);
  nand (_03269_, _03268_, _02744_);
  nand (_03270_, _03269_, _03259_);
  nand (_03271_, _03270_, _02761_);
  nand (_03272_, _03271_, _03248_);
  and (_03273_, _02857_, _01929_);
  not (_03274_, _03273_);
  and (_03275_, _03274_, _03272_);
  and (_03276_, _03273_, _02263_);
  or (_03277_, _03276_, _03189_);
  nor (_03278_, _03277_, _03275_);
  nor (_03279_, _03278_, _03198_);
  and (_03280_, _03189_, _02441_);
  not (_03281_, _03280_);
  nand (_03282_, _02375_, \oc8051_golden_model_1.IRAM[3] [0]);
  nand (_03283_, _02744_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_03284_, _03283_, _03282_);
  or (_03285_, _03284_, _02731_);
  nand (_03286_, _02375_, \oc8051_golden_model_1.IRAM[2] [0]);
  nand (_03287_, _02744_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_03288_, _03287_, _03286_);
  or (_03289_, _03288_, _02574_);
  and (_03290_, _03289_, _02737_);
  and (_03291_, _03290_, _03285_);
  nand (_03292_, _02375_, \oc8051_golden_model_1.IRAM[1] [0]);
  nand (_03293_, _02744_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_03294_, _03293_, _03292_);
  or (_03295_, _03294_, _02731_);
  nand (_03296_, _02375_, \oc8051_golden_model_1.IRAM[0] [0]);
  nand (_03297_, _02744_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_03298_, _03297_, _03296_);
  or (_03299_, _03298_, _02574_);
  and (_03300_, _03299_, _02729_);
  and (_03301_, _03300_, _03295_);
  or (_03302_, _03301_, _03291_);
  nand (_03303_, _03302_, _02177_);
  not (_03304_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_03305_, _02574_, _03304_);
  not (_03306_, \oc8051_golden_model_1.IRAM[9] [0]);
  or (_03307_, _02731_, _03306_);
  and (_03308_, _03307_, _02729_);
  nand (_03309_, _03308_, _03305_);
  not (_03310_, \oc8051_golden_model_1.IRAM[11] [0]);
  or (_03311_, _02731_, _03310_);
  not (_03312_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_03313_, _02574_, _03312_);
  and (_03314_, _03313_, _02737_);
  nand (_03315_, _03314_, _03311_);
  nand (_03316_, _03315_, _03309_);
  nand (_03317_, _03316_, _02375_);
  not (_03318_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_03319_, _02731_, _03318_);
  not (_03320_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_03321_, _02574_, _03320_);
  and (_03322_, _03321_, _02737_);
  nand (_03323_, _03322_, _03319_);
  not (_03324_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_03325_, _02574_, _03324_);
  not (_03326_, \oc8051_golden_model_1.IRAM[13] [0]);
  or (_03327_, _02731_, _03326_);
  and (_03328_, _03327_, _02729_);
  nand (_03329_, _03328_, _03325_);
  nand (_03330_, _03329_, _03323_);
  nand (_03331_, _03330_, _02744_);
  nand (_03332_, _03331_, _03317_);
  nand (_03333_, _03332_, _02761_);
  and (_03334_, _03333_, _03303_);
  or (_03335_, _03334_, _03273_);
  and (_03336_, _03273_, _02409_);
  nor (_03337_, _03336_, _03189_);
  nand (_03338_, _03337_, _03335_);
  and (_03339_, _03338_, _03281_);
  nand (_03340_, _03339_, \oc8051_golden_model_1.IRAM[0] [3]);
  not (_03341_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_03342_, _02574_, _03341_);
  not (_03343_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_03344_, _02731_, _03343_);
  and (_03345_, _03344_, _02729_);
  nand (_03346_, _03345_, _03342_);
  not (_03347_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_03348_, _02731_, _03347_);
  not (_03349_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_03350_, _02574_, _03349_);
  and (_03351_, _03350_, _02737_);
  nand (_03352_, _03351_, _03348_);
  nand (_03353_, _03352_, _03346_);
  nand (_03354_, _03353_, _02375_);
  not (_03355_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_03356_, _02731_, _03355_);
  not (_03357_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_03358_, _02574_, _03357_);
  and (_03359_, _03358_, _02737_);
  nand (_03360_, _03359_, _03356_);
  not (_03361_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_03362_, _02574_, _03361_);
  not (_03363_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_03364_, _02731_, _03363_);
  and (_03365_, _03364_, _02729_);
  nand (_03366_, _03365_, _03362_);
  nand (_03367_, _03366_, _03360_);
  nand (_03368_, _03367_, _02744_);
  nand (_03369_, _03368_, _03354_);
  nand (_03370_, _03369_, _02177_);
  nand (_03371_, _02574_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_03372_, _02731_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_03373_, _03372_, _02737_);
  nand (_03374_, _03373_, _03371_);
  nand (_03375_, _02731_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand (_03376_, _02574_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_03377_, _03376_, _02729_);
  nand (_03378_, _03377_, _03375_);
  nand (_03379_, _03378_, _03374_);
  nand (_03380_, _03379_, _02375_);
  nand (_03381_, _02574_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_03382_, _02731_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_03383_, _03382_, _02737_);
  nand (_03384_, _03383_, _03381_);
  nand (_03385_, _02731_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand (_03386_, _02574_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_03387_, _03386_, _02729_);
  nand (_03388_, _03387_, _03385_);
  nand (_03389_, _03388_, _03384_);
  nand (_03390_, _03389_, _02744_);
  nand (_03391_, _03390_, _03380_);
  nand (_03392_, _03391_, _02761_);
  nand (_03393_, _03392_, _03370_);
  nor (_03394_, _03393_, _03273_);
  nor (_03395_, _03274_, _02643_);
  nor (_03396_, _03395_, _03189_);
  not (_03397_, _03396_);
  or (_03398_, _03397_, _03394_);
  and (_03399_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  nor (_03400_, _03399_, _03190_);
  and (_03401_, _03400_, _03189_);
  not (_03402_, _03401_);
  and (_03403_, _03402_, _03398_);
  not (_03404_, _03403_);
  not (_03405_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_03406_, _03339_, _03405_);
  and (_03407_, _03406_, _03404_);
  nand (_03408_, _03407_, _03340_);
  nand (_03409_, _03339_, \oc8051_golden_model_1.IRAM[2] [3]);
  not (_03410_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_03411_, _03339_, _03410_);
  and (_03412_, _03411_, _03403_);
  nand (_03413_, _03412_, _03409_);
  nand (_03414_, _03413_, _03408_);
  nand (_03415_, _03414_, _03279_);
  nor (_03416_, _03192_, _02160_);
  nor (_03417_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_03418_, _03417_, _02160_);
  and (_03419_, _03418_, _02441_);
  nor (_03420_, _03419_, _03416_);
  not (_03421_, _03420_);
  and (_03422_, _03421_, _03189_);
  not (_03423_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_03424_, _02574_, _03423_);
  or (_03425_, _02731_, _03405_);
  and (_03426_, _03425_, _02729_);
  nand (_03427_, _03426_, _03424_);
  or (_03428_, _02731_, _03410_);
  not (_03429_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_03430_, _02574_, _03429_);
  and (_03431_, _03430_, _02737_);
  nand (_03432_, _03431_, _03428_);
  nand (_03433_, _03432_, _03427_);
  nand (_03434_, _03433_, _02375_);
  not (_03435_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_03436_, _02731_, _03435_);
  not (_03437_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_03438_, _02574_, _03437_);
  and (_03439_, _03438_, _02737_);
  nand (_03440_, _03439_, _03436_);
  not (_03441_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_03442_, _02574_, _03441_);
  not (_03443_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_03444_, _02731_, _03443_);
  and (_03445_, _03444_, _02729_);
  nand (_03446_, _03445_, _03442_);
  nand (_03447_, _03446_, _03440_);
  nand (_03448_, _03447_, _02744_);
  nand (_03449_, _03448_, _03434_);
  nand (_03450_, _03449_, _02177_);
  nand (_03451_, _02574_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_03452_, _02731_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_03453_, _03452_, _02737_);
  nand (_03454_, _03453_, _03451_);
  nand (_03455_, _02731_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_03456_, _02574_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_03457_, _03456_, _02729_);
  nand (_03458_, _03457_, _03455_);
  nand (_03459_, _03458_, _03454_);
  nand (_03460_, _03459_, _02375_);
  nand (_03461_, _02574_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_03462_, _02731_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_03463_, _03462_, _02737_);
  nand (_03464_, _03463_, _03461_);
  nand (_03465_, _02731_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_03466_, _02574_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_03467_, _03466_, _02729_);
  nand (_03468_, _03467_, _03465_);
  nand (_03469_, _03468_, _03464_);
  nand (_03470_, _03469_, _02744_);
  nand (_03471_, _03470_, _03460_);
  nand (_03472_, _03471_, _02761_);
  nand (_03473_, _03472_, _03450_);
  and (_03474_, _03473_, _03274_);
  nor (_03475_, _03274_, _01916_);
  or (_03476_, _03475_, _03189_);
  nor (_03477_, _03476_, _03474_);
  nor (_03478_, _03477_, _03422_);
  not (_03479_, _03279_);
  nand (_03480_, _03339_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_03481_, _03339_, _03443_);
  and (_03482_, _03481_, _03404_);
  nand (_03483_, _03482_, _03480_);
  nand (_03484_, _03339_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_03485_, _03339_, _03435_);
  and (_03486_, _03485_, _03403_);
  nand (_03487_, _03486_, _03484_);
  nand (_03488_, _03487_, _03483_);
  nand (_03489_, _03488_, _03479_);
  and (_03490_, _03489_, _03478_);
  and (_03491_, _03490_, _03415_);
  not (_03492_, _03339_);
  or (_03493_, _03492_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_03494_, _03339_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_03495_, _03494_, _03493_);
  nand (_03496_, _03495_, _03403_);
  or (_03497_, _03492_, \oc8051_golden_model_1.IRAM[8] [3]);
  or (_03498_, _03339_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand (_03499_, _03498_, _03497_);
  nand (_03500_, _03499_, _03404_);
  nand (_03501_, _03500_, _03496_);
  nand (_03502_, _03501_, _03279_);
  not (_03503_, _03478_);
  or (_03504_, _03492_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_03505_, _03339_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_03506_, _03505_, _03504_);
  nand (_03507_, _03506_, _03403_);
  or (_03508_, _03492_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_03509_, _03339_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand (_03510_, _03509_, _03508_);
  nand (_03511_, _03510_, _03404_);
  nand (_03512_, _03511_, _03507_);
  nand (_03513_, _03512_, _03479_);
  and (_03514_, _03513_, _03503_);
  and (_03515_, _03514_, _03502_);
  or (_03516_, _03515_, _03491_);
  nor (_03517_, _03516_, _03188_);
  and (_03518_, _03516_, _03188_);
  nor (_03519_, _03518_, _03517_);
  nand (_03520_, _03339_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_03521_, _03339_, _03203_);
  and (_03522_, _03521_, _03404_);
  nand (_03523_, _03522_, _03520_);
  nand (_03524_, _03339_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_03525_, _03339_, _03209_);
  and (_03526_, _03525_, _03403_);
  nand (_03527_, _03526_, _03524_);
  nand (_03528_, _03527_, _03523_);
  nand (_03529_, _03528_, _03279_);
  nand (_03530_, _03339_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_03531_, _03339_, _03237_);
  and (_03532_, _03531_, _03404_);
  nand (_03533_, _03532_, _03530_);
  nand (_03534_, _03339_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_03535_, _03339_, _03222_);
  and (_03536_, _03535_, _03403_);
  nand (_03537_, _03536_, _03534_);
  nand (_03538_, _03537_, _03533_);
  nand (_03539_, _03538_, _03479_);
  and (_03540_, _03539_, _03478_);
  and (_03541_, _03540_, _03529_);
  nand (_03542_, _03339_, _03250_);
  or (_03543_, _03339_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_03544_, _03543_, _03542_);
  nand (_03545_, _03544_, _03403_);
  or (_03546_, _03492_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_03547_, _03339_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_03548_, _03547_, _03546_);
  nand (_03549_, _03548_, _03404_);
  nand (_03550_, _03549_, _03545_);
  nand (_03551_, _03550_, _03279_);
  or (_03552_, _03492_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_03553_, _03339_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_03554_, _03553_, _03552_);
  nand (_03555_, _03554_, _03403_);
  or (_03556_, _03492_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_03557_, _03339_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand (_03558_, _03557_, _03556_);
  nand (_03559_, _03558_, _03404_);
  nand (_03560_, _03559_, _03555_);
  nand (_03561_, _03560_, _03479_);
  and (_03562_, _03561_, _03503_);
  and (_03563_, _03562_, _03551_);
  or (_03564_, _03563_, _03541_);
  nand (_03565_, _03564_, _02263_);
  or (_03566_, _03564_, _02263_);
  and (_03567_, _03566_, _03565_);
  and (_03568_, _03567_, _03519_);
  nand (_03569_, _03339_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_03570_, _03339_, _03343_);
  and (_03571_, _03570_, _03404_);
  nand (_03572_, _03571_, _03569_);
  nand (_03573_, _03339_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_03574_, _03339_, _03347_);
  and (_03575_, _03574_, _03403_);
  nand (_03576_, _03575_, _03573_);
  nand (_03577_, _03576_, _03572_);
  nand (_03578_, _03577_, _03279_);
  nand (_03579_, _03339_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_03580_, _03339_, _03363_);
  and (_03581_, _03580_, _03404_);
  nand (_03582_, _03581_, _03579_);
  nand (_03583_, _03339_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_03584_, _03339_, _03355_);
  and (_03585_, _03584_, _03403_);
  nand (_03586_, _03585_, _03583_);
  nand (_03587_, _03586_, _03582_);
  nand (_03588_, _03587_, _03479_);
  and (_03589_, _03588_, _03478_);
  and (_03590_, _03589_, _03578_);
  or (_03591_, _03492_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_03592_, _03339_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_03593_, _03592_, _03591_);
  nand (_03594_, _03593_, _03403_);
  or (_03595_, _03492_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_03596_, _03339_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_03597_, _03596_, _03595_);
  nand (_03598_, _03597_, _03404_);
  nand (_03599_, _03598_, _03594_);
  nand (_03600_, _03599_, _03279_);
  or (_03601_, _03492_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_03602_, _03339_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_03603_, _03602_, _03601_);
  nand (_03604_, _03603_, _03403_);
  or (_03605_, _03492_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_03606_, _03339_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand (_03607_, _03606_, _03605_);
  nand (_03608_, _03607_, _03404_);
  nand (_03609_, _03608_, _03604_);
  nand (_03610_, _03609_, _03479_);
  and (_03611_, _03610_, _03503_);
  and (_03612_, _03611_, _03600_);
  or (_03613_, _03612_, _03590_);
  or (_03614_, _03613_, _02644_);
  nand (_03615_, _03613_, _02644_);
  nand (_03616_, _03615_, _03614_);
  nand (_03617_, _03339_, \oc8051_golden_model_1.IRAM[0] [0]);
  not (_03618_, \oc8051_golden_model_1.IRAM[1] [0]);
  or (_03619_, _03339_, _03618_);
  and (_03620_, _03619_, _03404_);
  nand (_03621_, _03620_, _03617_);
  nand (_03622_, _03339_, \oc8051_golden_model_1.IRAM[2] [0]);
  nand (_03623_, _03492_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_03624_, _03623_, _03403_);
  nand (_03625_, _03624_, _03622_);
  nand (_03627_, _03625_, _03621_);
  nand (_03629_, _03627_, _03279_);
  nand (_03631_, _03339_, \oc8051_golden_model_1.IRAM[4] [0]);
  nand (_03633_, _03492_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_03635_, _03633_, _03404_);
  nand (_03637_, _03635_, _03631_);
  nand (_03639_, _03339_, \oc8051_golden_model_1.IRAM[6] [0]);
  nand (_03641_, _03492_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_03643_, _03641_, _03403_);
  nand (_03645_, _03643_, _03639_);
  nand (_03647_, _03645_, _03637_);
  nand (_03649_, _03647_, _03479_);
  nand (_03651_, _03649_, _03629_);
  nand (_03653_, _03651_, _03478_);
  nand (_03655_, _03339_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_03656_, _03339_, _03310_);
  and (_03657_, _03656_, _03403_);
  nand (_03658_, _03657_, _03655_);
  nand (_03659_, _03339_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_03660_, _03339_, _03306_);
  and (_03661_, _03660_, _03404_);
  nand (_03662_, _03661_, _03659_);
  nand (_03663_, _03662_, _03658_);
  nand (_03664_, _03663_, _03279_);
  nand (_03665_, _03339_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_03666_, _03339_, _03326_);
  and (_03667_, _03666_, _03404_);
  nand (_03668_, _03667_, _03665_);
  nand (_03669_, _03339_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_03670_, _03339_, _03318_);
  and (_03671_, _03670_, _03403_);
  nand (_03672_, _03671_, _03669_);
  nand (_03673_, _03672_, _03668_);
  nand (_03674_, _03673_, _03479_);
  nand (_03675_, _03674_, _03664_);
  nand (_03676_, _03675_, _03503_);
  and (_03677_, _03676_, _03653_);
  or (_03678_, _03677_, _02409_);
  nand (_03679_, _03677_, _02409_);
  and (_03680_, _03679_, _03678_);
  and (_03681_, _03680_, _03616_);
  and (_03682_, _03681_, _03568_);
  not (_03683_, _01884_);
  nand (_03684_, _03339_, \oc8051_golden_model_1.IRAM[0] [6]);
  not (_03685_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_03687_, _03339_, _03685_);
  and (_03689_, _03687_, _03404_);
  nand (_03691_, _03689_, _03684_);
  nand (_03693_, _03339_, \oc8051_golden_model_1.IRAM[2] [6]);
  not (_03695_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_03697_, _03339_, _03695_);
  and (_03699_, _03697_, _03403_);
  nand (_03701_, _03699_, _03693_);
  nand (_03703_, _03701_, _03691_);
  nand (_03705_, _03703_, _03279_);
  nand (_03707_, _03339_, \oc8051_golden_model_1.IRAM[4] [6]);
  not (_03709_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_03711_, _03339_, _03709_);
  and (_03713_, _03711_, _03404_);
  nand (_03715_, _03713_, _03707_);
  nand (_03716_, _03339_, \oc8051_golden_model_1.IRAM[6] [6]);
  not (_03717_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_03718_, _03339_, _03717_);
  and (_03719_, _03718_, _03403_);
  nand (_03720_, _03719_, _03716_);
  nand (_03721_, _03720_, _03715_);
  nand (_03722_, _03721_, _03479_);
  and (_03723_, _03722_, _03478_);
  and (_03724_, _03723_, _03705_);
  or (_03725_, _03492_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_03726_, _03339_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_03727_, _03726_, _03725_);
  nand (_03728_, _03727_, _03403_);
  or (_03729_, _03492_, \oc8051_golden_model_1.IRAM[8] [6]);
  or (_03730_, _03339_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand (_03731_, _03730_, _03729_);
  nand (_03732_, _03731_, _03404_);
  nand (_03733_, _03732_, _03728_);
  nand (_03734_, _03733_, _03279_);
  or (_03735_, _03492_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_03736_, _03339_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_03737_, _03736_, _03735_);
  nand (_03738_, _03737_, _03403_);
  nand (_03739_, _03339_, \oc8051_golden_model_1.IRAM[12] [6]);
  not (_03740_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_03741_, _03339_, _03740_);
  and (_03742_, _03741_, _03739_);
  nand (_03743_, _03742_, _03404_);
  nand (_03744_, _03743_, _03738_);
  nand (_03745_, _03744_, _03479_);
  and (_03746_, _03745_, _03503_);
  and (_03747_, _03746_, _03734_);
  or (_03748_, _03747_, _03724_);
  or (_03749_, _03748_, _03683_);
  nand (_03750_, _03748_, _03683_);
  nand (_03751_, _03750_, _03749_);
  nand (_03752_, _03339_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_03753_, _03339_, _02730_);
  and (_03754_, _03753_, _03404_);
  nand (_03755_, _03754_, _03752_);
  nand (_03756_, _03339_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_03757_, _03339_, _02735_);
  and (_03758_, _03757_, _03403_);
  nand (_03759_, _03758_, _03756_);
  nand (_03760_, _03759_, _03755_);
  nand (_03761_, _03760_, _03279_);
  nand (_03762_, _03339_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_03763_, _03339_, _02753_);
  and (_03764_, _03763_, _03404_);
  nand (_03765_, _03764_, _03762_);
  nand (_03766_, _03339_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_03767_, _03339_, _02745_);
  and (_03768_, _03767_, _03403_);
  nand (_03769_, _03768_, _03766_);
  nand (_03770_, _03769_, _03765_);
  nand (_03771_, _03770_, _03479_);
  and (_03772_, _03771_, _03478_);
  and (_03773_, _03772_, _03761_);
  or (_03774_, _03492_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_03775_, _03339_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand (_03776_, _03775_, _03774_);
  nand (_03777_, _03776_, _03403_);
  or (_03778_, _03492_, \oc8051_golden_model_1.IRAM[8] [7]);
  or (_03779_, _03339_, \oc8051_golden_model_1.IRAM[9] [7]);
  nand (_03780_, _03779_, _03778_);
  nand (_03781_, _03780_, _03404_);
  nand (_03782_, _03781_, _03777_);
  nand (_03783_, _03782_, _03279_);
  or (_03784_, _03492_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_03785_, _03339_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_03786_, _03785_, _03784_);
  nand (_03787_, _03786_, _03403_);
  or (_03788_, _03492_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_03789_, _03339_, \oc8051_golden_model_1.IRAM[13] [7]);
  nand (_03790_, _03789_, _03788_);
  nand (_03791_, _03790_, _03404_);
  nand (_03792_, _03791_, _03787_);
  nand (_03793_, _03792_, _03479_);
  and (_03794_, _03793_, _03503_);
  and (_03795_, _03794_, _03783_);
  or (_03796_, _03795_, _03773_);
  or (_03797_, _03796_, _01853_);
  nand (_03798_, _03796_, _01853_);
  and (_03799_, _03798_, _03797_);
  and (_03800_, _03799_, _03751_);
  nand (_03801_, _03339_, \oc8051_golden_model_1.IRAM[0] [5]);
  not (_03802_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_03803_, _03339_, _03802_);
  and (_03804_, _03803_, _03404_);
  nand (_03805_, _03804_, _03801_);
  nand (_03806_, _03339_, \oc8051_golden_model_1.IRAM[2] [5]);
  not (_03807_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_03808_, _03339_, _03807_);
  and (_03809_, _03808_, _03403_);
  nand (_03810_, _03809_, _03806_);
  nand (_03811_, _03810_, _03805_);
  nand (_03812_, _03811_, _03279_);
  nand (_03813_, _03339_, \oc8051_golden_model_1.IRAM[4] [5]);
  not (_03814_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_03815_, _03339_, _03814_);
  and (_03816_, _03815_, _03404_);
  nand (_03817_, _03816_, _03813_);
  nand (_03818_, _03339_, \oc8051_golden_model_1.IRAM[6] [5]);
  not (_03819_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_03820_, _03339_, _03819_);
  and (_03821_, _03820_, _03403_);
  nand (_03822_, _03821_, _03818_);
  nand (_03823_, _03822_, _03817_);
  nand (_03824_, _03823_, _03479_);
  and (_03825_, _03824_, _03478_);
  and (_03826_, _03825_, _03812_);
  or (_03827_, _03492_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_03828_, _03339_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_03829_, _03828_, _03827_);
  nand (_03830_, _03829_, _03403_);
  or (_03831_, _03492_, \oc8051_golden_model_1.IRAM[8] [5]);
  or (_03832_, _03339_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand (_03833_, _03832_, _03831_);
  nand (_03834_, _03833_, _03404_);
  nand (_03835_, _03834_, _03830_);
  nand (_03836_, _03835_, _03279_);
  or (_03837_, _03492_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_03838_, _03339_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_03839_, _03838_, _03837_);
  nand (_03840_, _03839_, _03403_);
  nand (_03841_, _03339_, \oc8051_golden_model_1.IRAM[12] [5]);
  not (_03842_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_03843_, _03339_, _03842_);
  and (_03844_, _03843_, _03841_);
  nand (_03845_, _03844_, _03404_);
  nand (_03846_, _03845_, _03840_);
  nand (_03847_, _03846_, _03479_);
  and (_03848_, _03847_, _03503_);
  and (_03849_, _03848_, _03836_);
  or (_03850_, _03849_, _03826_);
  nor (_03851_, _03850_, _02214_);
  and (_03852_, _03850_, _02214_);
  nor (_03853_, _03852_, _03851_);
  nand (_03854_, _03339_, \oc8051_golden_model_1.IRAM[0] [4]);
  not (_03855_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_03856_, _03339_, _03855_);
  and (_03857_, _03856_, _03404_);
  nand (_03858_, _03857_, _03854_);
  nand (_03859_, _03339_, \oc8051_golden_model_1.IRAM[2] [4]);
  not (_03860_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_03861_, _03339_, _03860_);
  and (_03862_, _03861_, _03403_);
  nand (_03863_, _03862_, _03859_);
  nand (_03864_, _03863_, _03858_);
  nand (_03865_, _03864_, _03279_);
  nand (_03866_, _03339_, \oc8051_golden_model_1.IRAM[4] [4]);
  not (_03867_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_03868_, _03339_, _03867_);
  and (_03869_, _03868_, _03404_);
  nand (_03870_, _03869_, _03866_);
  nand (_03871_, _03339_, \oc8051_golden_model_1.IRAM[6] [4]);
  not (_03872_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_03873_, _03339_, _03872_);
  and (_03874_, _03873_, _03403_);
  nand (_03875_, _03874_, _03871_);
  nand (_03876_, _03875_, _03870_);
  nand (_03877_, _03876_, _03479_);
  and (_03878_, _03877_, _03478_);
  and (_03879_, _03878_, _03865_);
  or (_03880_, _03492_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_03881_, _03339_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_03882_, _03881_, _03880_);
  nand (_03883_, _03882_, _03403_);
  or (_03884_, _03492_, \oc8051_golden_model_1.IRAM[8] [4]);
  or (_03885_, _03339_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand (_03886_, _03885_, _03884_);
  nand (_03887_, _03886_, _03404_);
  nand (_03888_, _03887_, _03883_);
  nand (_03889_, _03888_, _03279_);
  or (_03890_, _03492_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_03891_, _03339_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_03892_, _03891_, _03890_);
  nand (_03893_, _03892_, _03403_);
  nand (_03894_, _03339_, \oc8051_golden_model_1.IRAM[12] [4]);
  not (_03895_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_03896_, _03339_, _03895_);
  and (_03897_, _03896_, _03894_);
  nand (_03898_, _03897_, _03404_);
  nand (_03899_, _03898_, _03893_);
  nand (_03900_, _03899_, _03479_);
  and (_03901_, _03900_, _03503_);
  and (_03902_, _03901_, _03889_);
  or (_03903_, _03902_, _03879_);
  or (_03904_, _03903_, _02606_);
  nand (_03905_, _03903_, _02606_);
  and (_03906_, _03905_, _03904_);
  and (_03907_, _03906_, _03853_);
  and (_03908_, _03907_, _03800_);
  and (_03909_, _03908_, _03682_);
  or (_03910_, _03909_, _03176_);
  nand (_03911_, _03909_, _03168_);
  and (_03912_, _03911_, _03910_);
  or (_03913_, _03912_, _03187_);
  and (_03914_, _03393_, _02644_);
  nor (_03915_, _03393_, _02644_);
  nor (_03916_, _03915_, _03914_);
  nand (_03917_, _03333_, _03303_);
  and (_03918_, _03917_, _02478_);
  and (_03919_, _03334_, _02409_);
  or (_03920_, _03919_, _03918_);
  not (_03921_, _03920_);
  and (_03922_, _03921_, _03916_);
  and (_03923_, _03272_, _02264_);
  nor (_03924_, _03272_, _02264_);
  or (_03925_, _03924_, _03923_);
  not (_03926_, _03925_);
  and (_03927_, _03473_, _01916_);
  nor (_03928_, _03473_, _01916_);
  nor (_03929_, _03928_, _03927_);
  and (_03930_, _03929_, _03926_);
  and (_03931_, _03930_, _03922_);
  nand (_03932_, _02731_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_03933_, _02731_, _03802_);
  and (_03934_, _03933_, _02729_);
  nand (_03935_, _03934_, _03932_);
  or (_03936_, _02731_, _03807_);
  nand (_03937_, _02731_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_03938_, _03937_, _02737_);
  nand (_03939_, _03938_, _03936_);
  nand (_03940_, _03939_, _03935_);
  nand (_03941_, _03940_, _02375_);
  or (_03942_, _02731_, _03819_);
  nand (_03943_, _02731_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_03944_, _03943_, _02737_);
  nand (_03945_, _03944_, _03942_);
  nand (_03946_, _02731_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_03947_, _02731_, _03814_);
  and (_03948_, _03947_, _02729_);
  nand (_03949_, _03948_, _03946_);
  nand (_03950_, _03949_, _03945_);
  nand (_03951_, _03950_, _02744_);
  nand (_03952_, _03951_, _03941_);
  nand (_03953_, _03952_, _02177_);
  nand (_03954_, _02574_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_03955_, _02731_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_03956_, _03955_, _02737_);
  nand (_03957_, _03956_, _03954_);
  nand (_03958_, _02731_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand (_03959_, _02574_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_03960_, _03959_, _02729_);
  nand (_03961_, _03960_, _03958_);
  nand (_03962_, _03961_, _03957_);
  nand (_03963_, _03962_, _02375_);
  nand (_03964_, _02574_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_03965_, _02731_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_03966_, _03965_, _02737_);
  nand (_03967_, _03966_, _03964_);
  nand (_03968_, _02731_, \oc8051_golden_model_1.IRAM[12] [5]);
  or (_03969_, _02731_, _03842_);
  and (_03970_, _03969_, _02729_);
  nand (_03971_, _03970_, _03968_);
  nand (_03972_, _03971_, _03967_);
  nand (_03973_, _03972_, _02744_);
  nand (_03974_, _03973_, _03963_);
  nand (_03975_, _03974_, _02761_);
  nand (_03976_, _03975_, _03953_);
  and (_03977_, _03976_, _02216_);
  nor (_03978_, _03976_, _02216_);
  nor (_03979_, _03978_, _03977_);
  nand (_03980_, _02731_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_03981_, _02731_, _03855_);
  and (_03982_, _03981_, _02729_);
  nand (_03983_, _03982_, _03980_);
  or (_03984_, _02731_, _03860_);
  nand (_03985_, _02731_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_03986_, _03985_, _02737_);
  nand (_03987_, _03986_, _03984_);
  nand (_03988_, _03987_, _03983_);
  nand (_03989_, _03988_, _02375_);
  or (_03990_, _02731_, _03872_);
  nand (_03991_, _02731_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_03992_, _03991_, _02737_);
  nand (_03993_, _03992_, _03990_);
  nand (_03994_, _02731_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_03995_, _02731_, _03867_);
  and (_03996_, _03995_, _02729_);
  nand (_03997_, _03996_, _03994_);
  nand (_03998_, _03997_, _03993_);
  nand (_03999_, _03998_, _02744_);
  nand (_04000_, _03999_, _03989_);
  nand (_04001_, _04000_, _02177_);
  nand (_04002_, _02574_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_04003_, _02731_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_04004_, _04003_, _02737_);
  nand (_04005_, _04004_, _04002_);
  nand (_04006_, _02731_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand (_04007_, _02574_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_04008_, _04007_, _02729_);
  nand (_04009_, _04008_, _04006_);
  nand (_04010_, _04009_, _04005_);
  nand (_04011_, _04010_, _02375_);
  nand (_04012_, _02574_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_04013_, _02731_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_04014_, _04013_, _02737_);
  nand (_04015_, _04014_, _04012_);
  nand (_04016_, _02731_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_04017_, _02731_, _03895_);
  and (_04018_, _04017_, _02729_);
  nand (_04019_, _04018_, _04016_);
  nand (_04020_, _04019_, _04015_);
  nand (_04021_, _04020_, _02744_);
  nand (_04022_, _04021_, _04011_);
  nand (_04023_, _04022_, _02761_);
  nand (_04024_, _04023_, _04001_);
  and (_04025_, _04024_, _02607_);
  nor (_04026_, _04024_, _02607_);
  or (_04027_, _04026_, _04025_);
  not (_04028_, _04027_);
  and (_04029_, _04028_, _03979_);
  nand (_04030_, _02731_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_04031_, _02731_, _03685_);
  and (_04032_, _04031_, _02729_);
  nand (_04033_, _04032_, _04030_);
  or (_04034_, _02731_, _03695_);
  nand (_04035_, _02731_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_04036_, _04035_, _02737_);
  nand (_04037_, _04036_, _04034_);
  nand (_04038_, _04037_, _04033_);
  nand (_04039_, _04038_, _02375_);
  or (_04040_, _02731_, _03717_);
  nand (_04041_, _02731_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_04042_, _04041_, _02737_);
  nand (_04043_, _04042_, _04040_);
  nand (_04044_, _02731_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_04045_, _02731_, _03709_);
  and (_04046_, _04045_, _02729_);
  nand (_04047_, _04046_, _04044_);
  nand (_04048_, _04047_, _04043_);
  nand (_04049_, _04048_, _02744_);
  nand (_04050_, _04049_, _04039_);
  nand (_04051_, _04050_, _02177_);
  nand (_04052_, _02574_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_04053_, _02731_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_04054_, _04053_, _02737_);
  nand (_04055_, _04054_, _04052_);
  nand (_04056_, _02731_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_04057_, _02574_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_04058_, _04057_, _02729_);
  nand (_04059_, _04058_, _04056_);
  nand (_04060_, _04059_, _04055_);
  nand (_04061_, _04060_, _02375_);
  nand (_04062_, _02574_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_04063_, _02731_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_04064_, _04063_, _02737_);
  nand (_04065_, _04064_, _04062_);
  nand (_04066_, _02731_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_04067_, _02731_, _03740_);
  and (_04068_, _04067_, _02729_);
  nand (_04069_, _04068_, _04066_);
  nand (_04070_, _04069_, _04065_);
  nand (_04071_, _04070_, _02744_);
  nand (_04072_, _04071_, _04061_);
  nand (_04073_, _04072_, _02761_);
  nand (_04074_, _04073_, _04051_);
  nor (_04075_, _04074_, _03683_);
  and (_04076_, _04074_, _03683_);
  or (_04077_, _04076_, _04075_);
  not (_04078_, _04077_);
  or (_04079_, _02786_, _02220_);
  not (_04080_, _04079_);
  and (_04081_, _02786_, _02220_);
  nor (_04082_, _04081_, _04080_);
  and (_04083_, _04082_, _04078_);
  and (_04084_, _04083_, _04029_);
  and (_04085_, _04084_, _03931_);
  or (_04086_, _04085_, _03176_);
  nand (_04087_, _04085_, _03168_);
  and (_04088_, _04087_, _04086_);
  nor (_04089_, _01631_, _01591_);
  not (_04090_, _04089_);
  or (_04091_, _04090_, _04088_);
  and (_04092_, _02851_, _01963_);
  nor (_04093_, _02852_, _01610_);
  nor (_04094_, _04093_, _01620_);
  or (_04095_, _03473_, _02220_);
  and (_04096_, _01884_, _02220_);
  and (_04097_, _04096_, _02214_);
  and (_04098_, _04097_, _02606_);
  and (_04099_, _04098_, _03188_);
  nor (_04100_, _02643_, _02409_);
  and (_04101_, _04100_, _02263_);
  and (_04102_, _04101_, _04099_);
  and (_04103_, _04102_, \oc8051_golden_model_1.DPH [3]);
  not (_04104_, _04103_);
  nor (_04105_, _02643_, _02478_);
  and (_04106_, _04105_, _02263_);
  and (_04107_, _04106_, _04099_);
  and (_04108_, _04107_, \oc8051_golden_model_1.DPL [3]);
  and (_04109_, _02643_, _02478_);
  and (_04110_, _04109_, _02263_);
  and (_04111_, _04110_, _04099_);
  and (_04112_, _04111_, \oc8051_golden_model_1.SP [3]);
  nor (_04113_, _04112_, _04108_);
  and (_04114_, _04113_, _04104_);
  and (_04115_, _02643_, _02409_);
  not (_04116_, _04115_);
  nand (_04117_, _02263_, _01916_);
  nor (_04118_, _04117_, _04116_);
  and (_04119_, _04118_, _04098_);
  and (_04120_, _04119_, \oc8051_golden_model_1.TCON [3]);
  not (_04121_, _04120_);
  not (_04122_, _04098_);
  or (_04123_, _02263_, _03188_);
  or (_04124_, _04123_, _04116_);
  nor (_04125_, _04124_, _04122_);
  and (_04126_, _04125_, \oc8051_golden_model_1.TH0 [3]);
  and (_04127_, _02607_, _02214_);
  and (_04128_, _04127_, _04096_);
  and (_04129_, _04128_, _04118_);
  and (_04130_, _04129_, \oc8051_golden_model_1.SCON [3]);
  nor (_04131_, _04130_, _04126_);
  and (_04132_, _04131_, _04121_);
  and (_04133_, _04110_, _01916_);
  and (_04134_, _04133_, _04098_);
  and (_04135_, _04134_, \oc8051_golden_model_1.TMOD [3]);
  not (_04136_, _04109_);
  or (_04137_, _04123_, _04136_);
  nor (_04138_, _04137_, _04122_);
  and (_04139_, _04138_, \oc8051_golden_model_1.TH1 [3]);
  nor (_04140_, _04139_, _04135_);
  not (_04141_, _04105_);
  or (_04142_, _04117_, _04141_);
  nor (_04143_, _04142_, _04122_);
  and (_04144_, _04143_, \oc8051_golden_model_1.TL0 [3]);
  not (_04145_, _04100_);
  or (_04146_, _04117_, _04145_);
  nor (_04147_, _04146_, _04122_);
  and (_04148_, _04147_, \oc8051_golden_model_1.TL1 [3]);
  nor (_04149_, _04148_, _04144_);
  and (_04150_, _04149_, _04140_);
  and (_04151_, _04150_, _04132_);
  and (_04152_, _04151_, _04114_);
  nor (_04153_, _02606_, _02214_);
  and (_04154_, _04153_, _04096_);
  and (_04155_, _04154_, _04118_);
  and (_04156_, _04155_, \oc8051_golden_model_1.IP [3]);
  and (_04157_, _04115_, _02263_);
  nand (_04158_, _04157_, _03188_);
  and (_04159_, _02606_, _02216_);
  nor (_04160_, _01884_, _01853_);
  and (_04161_, _04160_, _04159_);
  not (_04162_, _04161_);
  nor (_04163_, _04162_, _04158_);
  and (_04164_, _04163_, \oc8051_golden_model_1.ACC [3]);
  nor (_04165_, _04164_, _04156_);
  and (_04166_, _04160_, _04127_);
  not (_04167_, _04166_);
  nor (_04168_, _04167_, _04158_);
  and (_04169_, _04168_, \oc8051_golden_model_1.PSW [3]);
  and (_04170_, _04160_, _04153_);
  not (_04171_, _04170_);
  nor (_04172_, _04171_, _04158_);
  and (_04173_, _04172_, \oc8051_golden_model_1.B [3]);
  nor (_04174_, _04173_, _04169_);
  and (_04175_, _04174_, _04165_);
  and (_04176_, _04100_, _02264_);
  and (_04177_, _04176_, _04099_);
  and (_04178_, _04177_, \oc8051_golden_model_1.PCON [3]);
  not (_04179_, _04178_);
  and (_04180_, _04133_, _04128_);
  and (_04181_, _04180_, \oc8051_golden_model_1.SBUF [3]);
  and (_04182_, _04159_, _04096_);
  and (_04183_, _04182_, _04118_);
  and (_04184_, _04183_, \oc8051_golden_model_1.IE [3]);
  nor (_04185_, _04184_, _04181_);
  and (_04186_, _04185_, _04179_);
  and (_04187_, _04186_, _04175_);
  and (_04188_, _04157_, _04099_);
  nand (_04189_, _04188_, \oc8051_golden_model_1.P0 [3]);
  not (_04190_, _04182_);
  nor (_04191_, _04190_, _04158_);
  and (_04192_, _04191_, \oc8051_golden_model_1.P2 [3]);
  not (_04193_, _04128_);
  nor (_04194_, _04158_, _04193_);
  and (_04195_, _04194_, \oc8051_golden_model_1.P1 [3]);
  not (_04196_, _04154_);
  nor (_04197_, _04158_, _04196_);
  and (_04198_, _04197_, \oc8051_golden_model_1.P3 [3]);
  or (_04199_, _04198_, _04195_);
  nor (_04200_, _04199_, _04192_);
  and (_04201_, _04200_, _04189_);
  and (_04202_, _04201_, _04187_);
  and (_04203_, _04202_, _04152_);
  and (_04204_, _04203_, _04095_);
  or (_04205_, _03272_, _02220_);
  and (_04206_, _04111_, \oc8051_golden_model_1.SP [2]);
  not (_04207_, _04206_);
  and (_04208_, _04107_, \oc8051_golden_model_1.DPL [2]);
  and (_04209_, _04102_, \oc8051_golden_model_1.DPH [2]);
  nor (_04210_, _04209_, _04208_);
  and (_04211_, _04210_, _04207_);
  and (_04212_, _04143_, \oc8051_golden_model_1.TL0 [2]);
  not (_04213_, _04212_);
  and (_04214_, _04147_, \oc8051_golden_model_1.TL1 [2]);
  and (_04215_, _04138_, \oc8051_golden_model_1.TH1 [2]);
  nor (_04216_, _04215_, _04214_);
  and (_04217_, _04216_, _04213_);
  and (_04218_, _04125_, \oc8051_golden_model_1.TH0 [2]);
  and (_04219_, _04163_, \oc8051_golden_model_1.ACC [2]);
  nor (_04220_, _04219_, _04218_);
  and (_04221_, _04119_, \oc8051_golden_model_1.TCON [2]);
  and (_04222_, _04134_, \oc8051_golden_model_1.TMOD [2]);
  nor (_04223_, _04222_, _04221_);
  and (_04224_, _04223_, _04220_);
  and (_04225_, _04129_, \oc8051_golden_model_1.SCON [2]);
  and (_04226_, _04155_, \oc8051_golden_model_1.IP [2]);
  nor (_04227_, _04226_, _04225_);
  and (_04228_, _04168_, \oc8051_golden_model_1.PSW [2]);
  and (_04229_, _04172_, \oc8051_golden_model_1.B [2]);
  nor (_04230_, _04229_, _04228_);
  and (_04231_, _04230_, _04227_);
  and (_04232_, _04231_, _04224_);
  and (_04233_, _04232_, _04217_);
  and (_04234_, _04233_, _04211_);
  and (_04235_, _04177_, \oc8051_golden_model_1.PCON [2]);
  not (_04236_, _04235_);
  and (_04237_, _04180_, \oc8051_golden_model_1.SBUF [2]);
  and (_04238_, _04183_, \oc8051_golden_model_1.IE [2]);
  nor (_04239_, _04238_, _04237_);
  and (_04240_, _04239_, _04236_);
  and (_04241_, _04188_, \oc8051_golden_model_1.P0 [2]);
  not (_04242_, _04241_);
  and (_04243_, _04194_, \oc8051_golden_model_1.P1 [2]);
  not (_04244_, _04243_);
  and (_04245_, _04191_, \oc8051_golden_model_1.P2 [2]);
  and (_04246_, _04197_, \oc8051_golden_model_1.P3 [2]);
  nor (_04247_, _04246_, _04245_);
  and (_04248_, _04247_, _04244_);
  and (_04249_, _04248_, _04242_);
  and (_04250_, _04249_, _04240_);
  and (_04251_, _04250_, _04234_);
  and (_04252_, _04251_, _04205_);
  and (_04253_, _04252_, _04204_);
  or (_04254_, _04024_, _02220_);
  and (_04255_, _04111_, \oc8051_golden_model_1.SP [4]);
  and (_04256_, _04102_, \oc8051_golden_model_1.DPH [4]);
  nor (_04257_, _04256_, _04255_);
  and (_04258_, _04177_, \oc8051_golden_model_1.PCON [4]);
  and (_04259_, _04107_, \oc8051_golden_model_1.DPL [4]);
  nor (_04260_, _04259_, _04258_);
  and (_04261_, _04260_, _04257_);
  and (_04262_, _04125_, \oc8051_golden_model_1.TH0 [4]);
  and (_04263_, _04138_, \oc8051_golden_model_1.TH1 [4]);
  nor (_04264_, _04263_, _04262_);
  and (_04265_, _04143_, \oc8051_golden_model_1.TL0 [4]);
  and (_04266_, _04147_, \oc8051_golden_model_1.TL1 [4]);
  nor (_04267_, _04266_, _04265_);
  and (_04268_, _04267_, _04264_);
  and (_04269_, _04129_, \oc8051_golden_model_1.SCON [4]);
  and (_04270_, _04183_, \oc8051_golden_model_1.IE [4]);
  nor (_04271_, _04270_, _04269_);
  and (_04272_, _04134_, \oc8051_golden_model_1.TMOD [4]);
  and (_04273_, _04180_, \oc8051_golden_model_1.SBUF [4]);
  nor (_04274_, _04273_, _04272_);
  and (_04275_, _04274_, _04271_);
  and (_04276_, _04275_, _04268_);
  and (_04277_, _04276_, _04261_);
  and (_04278_, _04155_, \oc8051_golden_model_1.IP [4]);
  and (_04279_, _04163_, \oc8051_golden_model_1.ACC [4]);
  nor (_04280_, _04279_, _04278_);
  and (_04281_, _04119_, \oc8051_golden_model_1.TCON [4]);
  not (_04282_, _04281_);
  and (_04283_, _04168_, \oc8051_golden_model_1.PSW [4]);
  and (_04284_, _04172_, \oc8051_golden_model_1.B [4]);
  nor (_04285_, _04284_, _04283_);
  and (_04286_, _04285_, _04282_);
  and (_04287_, _04286_, _04280_);
  and (_04288_, _04188_, \oc8051_golden_model_1.P0 [4]);
  not (_04289_, _04288_);
  and (_04290_, _04194_, \oc8051_golden_model_1.P1 [4]);
  not (_04291_, _04290_);
  and (_04292_, _04191_, \oc8051_golden_model_1.P2 [4]);
  and (_04293_, _04197_, \oc8051_golden_model_1.P3 [4]);
  nor (_04294_, _04293_, _04292_);
  and (_04295_, _04294_, _04291_);
  and (_04296_, _04295_, _04289_);
  and (_04297_, _04296_, _04287_);
  and (_04298_, _04297_, _04277_);
  and (_04299_, _04298_, _04254_);
  or (_04300_, _03976_, _02220_);
  and (_04301_, _04102_, \oc8051_golden_model_1.DPH [5]);
  not (_04302_, _04301_);
  and (_04303_, _04107_, \oc8051_golden_model_1.DPL [5]);
  and (_04304_, _04111_, \oc8051_golden_model_1.SP [5]);
  nor (_04305_, _04304_, _04303_);
  and (_04306_, _04305_, _04302_);
  and (_04307_, _04119_, \oc8051_golden_model_1.TCON [5]);
  not (_04308_, _04307_);
  and (_04309_, _04125_, \oc8051_golden_model_1.TH0 [5]);
  and (_04310_, _04129_, \oc8051_golden_model_1.SCON [5]);
  nor (_04311_, _04310_, _04309_);
  and (_04312_, _04311_, _04308_);
  and (_04313_, _04134_, \oc8051_golden_model_1.TMOD [5]);
  and (_04314_, _04138_, \oc8051_golden_model_1.TH1 [5]);
  nor (_04315_, _04314_, _04313_);
  and (_04316_, _04143_, \oc8051_golden_model_1.TL0 [5]);
  and (_04317_, _04147_, \oc8051_golden_model_1.TL1 [5]);
  nor (_04318_, _04317_, _04316_);
  and (_04319_, _04318_, _04315_);
  and (_04320_, _04319_, _04312_);
  and (_04321_, _04320_, _04306_);
  and (_04322_, _04155_, \oc8051_golden_model_1.IP [5]);
  and (_04323_, _04172_, \oc8051_golden_model_1.B [5]);
  nor (_04324_, _04323_, _04322_);
  and (_04325_, _04168_, \oc8051_golden_model_1.PSW [5]);
  and (_04326_, _04163_, \oc8051_golden_model_1.ACC [5]);
  nor (_04327_, _04326_, _04325_);
  and (_04328_, _04327_, _04324_);
  and (_04329_, _04177_, \oc8051_golden_model_1.PCON [5]);
  not (_04330_, _04329_);
  and (_04331_, _04180_, \oc8051_golden_model_1.SBUF [5]);
  and (_04332_, _04183_, \oc8051_golden_model_1.IE [5]);
  nor (_04333_, _04332_, _04331_);
  and (_04334_, _04333_, _04330_);
  and (_04335_, _04334_, _04328_);
  and (_04336_, _04188_, \oc8051_golden_model_1.P0 [5]);
  not (_04337_, _04336_);
  and (_04338_, _04194_, \oc8051_golden_model_1.P1 [5]);
  not (_04339_, _04338_);
  and (_04340_, _04191_, \oc8051_golden_model_1.P2 [5]);
  and (_04341_, _04197_, \oc8051_golden_model_1.P3 [5]);
  nor (_04342_, _04341_, _04340_);
  and (_04343_, _04342_, _04339_);
  and (_04344_, _04343_, _04337_);
  and (_04345_, _04344_, _04335_);
  and (_04346_, _04345_, _04321_);
  and (_04347_, _04346_, _04300_);
  and (_04348_, _04347_, _04299_);
  and (_04349_, _04348_, _04253_);
  or (_04350_, _03917_, _02220_);
  and (_04351_, _04191_, \oc8051_golden_model_1.P2 [0]);
  and (_04352_, _04197_, \oc8051_golden_model_1.P3 [0]);
  nor (_04353_, _04352_, _04351_);
  and (_04354_, _04177_, \oc8051_golden_model_1.PCON [0]);
  not (_04355_, _04354_);
  and (_04356_, _04180_, \oc8051_golden_model_1.SBUF [0]);
  and (_04357_, _04183_, \oc8051_golden_model_1.IE [0]);
  nor (_04358_, _04357_, _04356_);
  and (_04359_, _04358_, _04355_);
  and (_04360_, _04359_, _04353_);
  and (_04361_, _04168_, \oc8051_golden_model_1.PSW [0]);
  not (_04362_, _04361_);
  and (_04363_, _04163_, \oc8051_golden_model_1.ACC [0]);
  and (_04364_, _04172_, \oc8051_golden_model_1.B [0]);
  nor (_04365_, _04364_, _04363_);
  and (_04366_, _04155_, \oc8051_golden_model_1.IP [0]);
  not (_04367_, _04366_);
  and (_04368_, _04367_, _04365_);
  and (_04369_, _04368_, _04362_);
  and (_04370_, _04125_, \oc8051_golden_model_1.TH0 [0]);
  and (_04371_, _04119_, \oc8051_golden_model_1.TCON [0]);
  nor (_04372_, _04371_, _04370_);
  and (_04373_, _04147_, \oc8051_golden_model_1.TL1 [0]);
  and (_04374_, _04194_, \oc8051_golden_model_1.P1 [0]);
  nor (_04375_, _04374_, _04373_);
  and (_04376_, _04375_, _04372_);
  and (_04377_, _04134_, \oc8051_golden_model_1.TMOD [0]);
  and (_04378_, _04143_, \oc8051_golden_model_1.TL0 [0]);
  nor (_04379_, _04378_, _04377_);
  and (_04380_, _04129_, \oc8051_golden_model_1.SCON [0]);
  and (_04381_, _04138_, \oc8051_golden_model_1.TH1 [0]);
  nor (_04382_, _04381_, _04380_);
  and (_04383_, _04382_, _04379_);
  and (_04384_, _04383_, _04376_);
  and (_04385_, _04384_, _04369_);
  and (_04386_, _04385_, _04360_);
  nor (_04387_, _04158_, _04122_);
  and (_04388_, _04387_, \oc8051_golden_model_1.P0 [0]);
  not (_04389_, _04388_);
  nand (_04390_, _02263_, _03188_);
  nor (_04391_, _04390_, _04145_);
  and (_04392_, _04391_, _04098_);
  and (_04393_, _04392_, \oc8051_golden_model_1.DPH [0]);
  not (_04394_, _04393_);
  or (_04395_, _04390_, _04136_);
  nor (_04396_, _04395_, _04122_);
  and (_04397_, _04396_, \oc8051_golden_model_1.SP [0]);
  nor (_04398_, _04390_, _04141_);
  and (_04399_, _04398_, _04098_);
  and (_04400_, _04399_, \oc8051_golden_model_1.DPL [0]);
  nor (_04401_, _04400_, _04397_);
  and (_04402_, _04401_, _04394_);
  and (_04403_, _04402_, _04389_);
  and (_04404_, _04403_, _04386_);
  nand (_04405_, _04404_, _04350_);
  or (_04406_, _03393_, _02220_);
  and (_04407_, _04111_, \oc8051_golden_model_1.SP [1]);
  not (_04408_, _04407_);
  and (_04409_, _04102_, \oc8051_golden_model_1.DPH [1]);
  and (_04410_, _04107_, \oc8051_golden_model_1.DPL [1]);
  nor (_04411_, _04410_, _04409_);
  and (_04412_, _04411_, _04408_);
  and (_04413_, _04168_, \oc8051_golden_model_1.PSW [1]);
  not (_04414_, _04413_);
  and (_04415_, _04163_, \oc8051_golden_model_1.ACC [1]);
  and (_04416_, _04172_, \oc8051_golden_model_1.B [1]);
  nor (_04417_, _04416_, _04415_);
  and (_04418_, _04417_, _04414_);
  and (_04419_, _04119_, \oc8051_golden_model_1.TCON [1]);
  and (_04420_, _04138_, \oc8051_golden_model_1.TH1 [1]);
  nor (_04421_, _04420_, _04419_);
  and (_04422_, _04147_, \oc8051_golden_model_1.TL1 [1]);
  and (_04423_, _04129_, \oc8051_golden_model_1.SCON [1]);
  nor (_04424_, _04423_, _04422_);
  and (_04425_, _04424_, _04421_);
  and (_04426_, _04143_, \oc8051_golden_model_1.TL0 [1]);
  and (_04427_, _04155_, \oc8051_golden_model_1.IP [1]);
  nor (_04428_, _04427_, _04426_);
  and (_04429_, _04134_, \oc8051_golden_model_1.TMOD [1]);
  and (_04430_, _04125_, \oc8051_golden_model_1.TH0 [1]);
  nor (_04431_, _04430_, _04429_);
  and (_04432_, _04431_, _04428_);
  and (_04433_, _04432_, _04425_);
  and (_04434_, _04433_, _04418_);
  and (_04435_, _04434_, _04412_);
  not (_04436_, _04435_);
  and (_04437_, _04177_, \oc8051_golden_model_1.PCON [1]);
  not (_04438_, _04437_);
  and (_04439_, _04180_, \oc8051_golden_model_1.SBUF [1]);
  and (_04440_, _04183_, \oc8051_golden_model_1.IE [1]);
  nor (_04441_, _04440_, _04439_);
  and (_04442_, _04441_, _04438_);
  nand (_04443_, _04188_, \oc8051_golden_model_1.P0 [1]);
  and (_04444_, _04191_, \oc8051_golden_model_1.P2 [1]);
  and (_04445_, _04194_, \oc8051_golden_model_1.P1 [1]);
  and (_04446_, _04197_, \oc8051_golden_model_1.P3 [1]);
  or (_04447_, _04446_, _04445_);
  nor (_04448_, _04447_, _04444_);
  and (_04449_, _04448_, _04443_);
  nand (_04450_, _04449_, _04442_);
  nor (_04451_, _04450_, _04436_);
  and (_04452_, _04451_, _04406_);
  and (_04453_, _04452_, _04405_);
  or (_04454_, _04074_, _02220_);
  and (_04455_, _04177_, \oc8051_golden_model_1.PCON [6]);
  not (_04456_, _04455_);
  and (_04457_, _04180_, \oc8051_golden_model_1.SBUF [6]);
  and (_04458_, _04183_, \oc8051_golden_model_1.IE [6]);
  nor (_04459_, _04458_, _04457_);
  and (_04460_, _04459_, _04456_);
  and (_04461_, _04102_, \oc8051_golden_model_1.DPH [6]);
  not (_04462_, _04461_);
  and (_04463_, _04125_, \oc8051_golden_model_1.TH0 [6]);
  and (_04464_, _04147_, \oc8051_golden_model_1.TL1 [6]);
  nor (_04465_, _04464_, _04463_);
  and (_04466_, _04465_, _04462_);
  and (_04467_, _04466_, _04460_);
  and (_04468_, _04138_, \oc8051_golden_model_1.TH1 [6]);
  and (_04469_, _04129_, \oc8051_golden_model_1.SCON [6]);
  nor (_04470_, _04469_, _04468_);
  and (_04471_, _04134_, \oc8051_golden_model_1.TMOD [6]);
  and (_04472_, _04143_, \oc8051_golden_model_1.TL0 [6]);
  nor (_04473_, _04472_, _04471_);
  and (_04474_, _04473_, _04470_);
  and (_04475_, _04155_, \oc8051_golden_model_1.IP [6]);
  and (_04476_, _04172_, \oc8051_golden_model_1.B [6]);
  nor (_04477_, _04476_, _04475_);
  and (_04478_, _04168_, \oc8051_golden_model_1.PSW [6]);
  and (_04479_, _04163_, \oc8051_golden_model_1.ACC [6]);
  nor (_04480_, _04479_, _04478_);
  and (_04481_, _04480_, _04477_);
  and (_04482_, _04481_, _04474_);
  and (_04483_, _04482_, _04467_);
  and (_04484_, _04107_, \oc8051_golden_model_1.DPL [6]);
  not (_04485_, _04484_);
  and (_04486_, _04119_, \oc8051_golden_model_1.TCON [6]);
  and (_04487_, _04111_, \oc8051_golden_model_1.SP [6]);
  nor (_04488_, _04487_, _04486_);
  and (_04489_, _04488_, _04485_);
  and (_04490_, _04188_, \oc8051_golden_model_1.P0 [6]);
  not (_04491_, _04490_);
  and (_04492_, _04197_, \oc8051_golden_model_1.P3 [6]);
  not (_04493_, _04492_);
  and (_04494_, _04194_, \oc8051_golden_model_1.P1 [6]);
  and (_04495_, _04191_, \oc8051_golden_model_1.P2 [6]);
  nor (_04496_, _04495_, _04494_);
  and (_04497_, _04496_, _04493_);
  and (_04498_, _04497_, _04491_);
  and (_04499_, _04498_, _04489_);
  and (_04500_, _04499_, _04483_);
  and (_04501_, _04500_, _04454_);
  and (_04502_, _04155_, \oc8051_golden_model_1.IP [7]);
  not (_04503_, _04502_);
  and (_04504_, _04168_, \oc8051_golden_model_1.PSW [7]);
  not (_04505_, _04504_);
  and (_04506_, _04172_, \oc8051_golden_model_1.B [7]);
  and (_04507_, _04163_, \oc8051_golden_model_1.ACC [7]);
  nor (_04508_, _04507_, _04506_);
  and (_04509_, _04508_, _04505_);
  and (_04510_, _04509_, _04503_);
  and (_04511_, _04125_, \oc8051_golden_model_1.TH0 [7]);
  and (_04512_, _04119_, \oc8051_golden_model_1.TCON [7]);
  nor (_04513_, _04512_, _04511_);
  and (_04514_, _04147_, \oc8051_golden_model_1.TL1 [7]);
  and (_04515_, _04194_, \oc8051_golden_model_1.P1 [7]);
  nor (_04516_, _04515_, _04514_);
  and (_04517_, _04516_, _04513_);
  and (_04518_, _04134_, \oc8051_golden_model_1.TMOD [7]);
  and (_04519_, _04143_, \oc8051_golden_model_1.TL0 [7]);
  nor (_04520_, _04519_, _04518_);
  and (_04521_, _04129_, \oc8051_golden_model_1.SCON [7]);
  and (_04522_, _04138_, \oc8051_golden_model_1.TH1 [7]);
  nor (_04523_, _04522_, _04521_);
  and (_04524_, _04523_, _04520_);
  and (_04525_, _04524_, _04517_);
  and (_04526_, _04177_, \oc8051_golden_model_1.PCON [7]);
  not (_04527_, _04526_);
  and (_04528_, _04180_, \oc8051_golden_model_1.SBUF [7]);
  and (_04529_, _04183_, \oc8051_golden_model_1.IE [7]);
  nor (_04530_, _04529_, _04528_);
  and (_04531_, _04530_, _04527_);
  and (_04532_, _04197_, \oc8051_golden_model_1.P3 [7]);
  and (_04533_, _04191_, \oc8051_golden_model_1.P2 [7]);
  nor (_04534_, _04533_, _04532_);
  and (_04535_, _04534_, _04531_);
  and (_04536_, _04387_, \oc8051_golden_model_1.P0 [7]);
  not (_04537_, _04536_);
  and (_04538_, _04392_, \oc8051_golden_model_1.DPH [7]);
  not (_04539_, _04538_);
  and (_04540_, _04396_, \oc8051_golden_model_1.SP [7]);
  and (_04541_, _04399_, \oc8051_golden_model_1.DPL [7]);
  nor (_04542_, _04541_, _04540_);
  and (_04543_, _04542_, _04539_);
  and (_04544_, _04543_, _04537_);
  and (_04545_, _04544_, _04535_);
  and (_04546_, _04545_, _04525_);
  and (_04547_, _04546_, _04510_);
  and (_04548_, _04547_, _04079_);
  and (_04549_, _04548_, _04501_);
  and (_04550_, _04549_, _04453_);
  nand (_04551_, _04550_, _04349_);
  and (_04552_, _04551_, _03176_);
  and (_04553_, _04550_, _04349_);
  and (_04554_, _04553_, _02878_);
  or (_04555_, _04554_, _02438_);
  or (_04556_, _04555_, _04552_);
  nor (_04557_, _01620_, _01591_);
  not (_04558_, _01627_);
  and (_04559_, _02852_, _02412_);
  nor (_04560_, _02858_, _01624_);
  nor (_04561_, _04560_, _04559_);
  and (_04562_, _02852_, _01970_);
  nor (_04563_, _02858_, _01626_);
  nor (_04564_, _04563_, _04562_);
  and (_04565_, _04564_, _04561_);
  or (_04566_, _04565_, _02803_);
  not (_04567_, _04564_);
  not (_04568_, _01625_);
  or (_04569_, _04568_, \oc8051_golden_model_1.PC [15]);
  or (_04570_, _04569_, _01971_);
  and (_04571_, _02412_, _01593_);
  or (_04572_, _04571_, _04559_);
  or (_04573_, _04572_, _04570_);
  or (_04574_, _04573_, _04567_);
  or (_04575_, _04574_, _04560_);
  and (_04576_, _04575_, _04566_);
  or (_04577_, _04576_, _04558_);
  or (_04578_, _04571_, _04568_);
  nor (_04579_, _04578_, _01971_);
  and (_04580_, _04579_, _01627_);
  or (_04581_, _04580_, _02851_);
  and (_04582_, _04581_, _04577_);
  or (_04583_, _04582_, _04557_);
  nor (_04584_, _02840_, \oc8051_golden_model_1.PC [14]);
  nor (_04585_, _04584_, _02841_);
  not (_04586_, _04585_);
  nor (_04587_, _04586_, _01853_);
  and (_04588_, _04586_, _01853_);
  nor (_04589_, _04588_, _04587_);
  not (_04590_, _04589_);
  nor (_04591_, _02847_, \oc8051_golden_model_1.PC [13]);
  nor (_04592_, _04591_, _02848_);
  and (_04593_, _04592_, _02220_);
  nor (_04594_, _04592_, _02220_);
  nor (_04595_, _02838_, \oc8051_golden_model_1.PC [12]);
  nor (_04596_, _04595_, _02839_);
  not (_04597_, _04596_);
  nor (_04598_, _04597_, _01853_);
  nor (_04599_, _02844_, \oc8051_golden_model_1.PC [10]);
  nor (_04600_, _04599_, _02837_);
  not (_04601_, _04600_);
  nor (_04602_, _04601_, _01853_);
  not (_04603_, _04602_);
  nor (_04604_, _02837_, _02971_);
  and (_04605_, _02837_, _02971_);
  or (_04606_, _04605_, _04604_);
  not (_04607_, _04606_);
  nor (_04608_, _04607_, _01853_);
  and (_04609_, _04607_, _01853_);
  nor (_04610_, _04609_, _04608_);
  and (_04611_, _04601_, _01853_);
  nor (_04612_, _04611_, _04602_);
  and (_04613_, _04612_, _04610_);
  nor (_04614_, _02843_, \oc8051_golden_model_1.PC [9]);
  nor (_04615_, _04614_, _02844_);
  not (_04616_, _04615_);
  nor (_04617_, _04616_, _01853_);
  and (_04618_, _04616_, _01853_);
  nor (_04619_, _04618_, _04617_);
  and (_04620_, _02988_, _01718_);
  nor (_04621_, _04620_, \oc8051_golden_model_1.PC [7]);
  nor (_04622_, _04621_, _02836_);
  not (_04623_, _04622_);
  nor (_04624_, _04623_, _01853_);
  and (_04625_, _04623_, _01853_);
  and (_04626_, _02790_, _01718_);
  nor (_04627_, _04626_, \oc8051_golden_model_1.PC [6]);
  nor (_04628_, _04627_, _04620_);
  not (_04629_, _04628_);
  nor (_04630_, _04629_, _01884_);
  and (_04631_, _04629_, _01884_);
  nor (_04632_, _04631_, _04630_);
  not (_04633_, _04632_);
  and (_04634_, _01718_, \oc8051_golden_model_1.PC [4]);
  nor (_04635_, _04634_, \oc8051_golden_model_1.PC [5]);
  nor (_04636_, _04635_, _04626_);
  not (_04637_, _04636_);
  nor (_04638_, _04637_, _02214_);
  and (_04639_, _04637_, _02214_);
  nor (_04640_, _01718_, \oc8051_golden_model_1.PC [4]);
  nor (_04641_, _04640_, _04634_);
  not (_04642_, _04641_);
  nor (_04643_, _04642_, _02606_);
  and (_04644_, _01916_, _01720_);
  nor (_04645_, _01916_, _01720_);
  nor (_04646_, _02263_, _01792_);
  nor (_04647_, _02643_, \oc8051_golden_model_1.PC [1]);
  nor (_04648_, _02409_, _01325_);
  and (_04649_, _02643_, \oc8051_golden_model_1.PC [1]);
  nor (_04650_, _04649_, _04647_);
  and (_04651_, _04650_, _04648_);
  nor (_04652_, _04651_, _04647_);
  and (_04653_, _02263_, _01792_);
  nor (_04654_, _04653_, _04646_);
  not (_04655_, _04654_);
  nor (_04656_, _04655_, _04652_);
  nor (_04657_, _04656_, _04646_);
  nor (_04658_, _04657_, _04645_);
  nor (_04659_, _04658_, _04644_);
  and (_04660_, _04642_, _02606_);
  nor (_04661_, _04660_, _04643_);
  not (_04662_, _04661_);
  nor (_04663_, _04662_, _04659_);
  nor (_04664_, _04663_, _04643_);
  nor (_04665_, _04664_, _04639_);
  nor (_04666_, _04665_, _04638_);
  nor (_04667_, _04666_, _04633_);
  nor (_04668_, _04667_, _04630_);
  nor (_04669_, _04668_, _04625_);
  or (_04670_, _04669_, _04624_);
  nor (_04671_, _02836_, \oc8051_golden_model_1.PC [8]);
  nor (_04672_, _04671_, _02843_);
  not (_04673_, _04672_);
  nor (_04674_, _04673_, _01853_);
  and (_04675_, _04673_, _01853_);
  nor (_04676_, _04675_, _04674_);
  and (_04677_, _04676_, _04670_);
  and (_04678_, _04677_, _04619_);
  and (_04679_, _04678_, _04613_);
  nor (_04680_, _04674_, _04617_);
  not (_04681_, _04680_);
  and (_04682_, _04681_, _04613_);
  or (_04683_, _04682_, _04608_);
  nor (_04684_, _04683_, _04679_);
  and (_04685_, _04684_, _04603_);
  not (_04686_, _04685_);
  and (_04687_, _04597_, _01853_);
  nor (_04688_, _04687_, _04598_);
  and (_04689_, _04688_, _04686_);
  nor (_04690_, _04689_, _04598_);
  nor (_04691_, _04690_, _04594_);
  nor (_04692_, _04691_, _04593_);
  nor (_04693_, _04692_, _04590_);
  nor (_04694_, _04693_, _04587_);
  and (_04695_, _02855_, _01853_);
  nor (_04696_, _02855_, _01853_);
  nor (_04697_, _04696_, _04695_);
  and (_04698_, _04697_, _04694_);
  nor (_04699_, _04697_, _04694_);
  or (_04700_, _04699_, _04698_);
  and (_04701_, _03473_, _03272_);
  and (_04702_, _03976_, _04024_);
  and (_04703_, _04702_, _04701_);
  and (_04704_, _03393_, _03334_);
  and (_04705_, _04074_, _02786_);
  and (_04706_, _04705_, _04704_);
  nand (_04707_, _04706_, _04703_);
  and (_04708_, _04707_, _04700_);
  not (_04709_, _04557_);
  and (_04710_, _04706_, _04703_);
  and (_04711_, _04710_, _02851_);
  or (_04712_, _04711_, _04709_);
  or (_04713_, _04712_, _04708_);
  and (_04714_, _04713_, _04583_);
  and (_04715_, _02857_, _01958_);
  or (_04716_, _04715_, _01969_);
  or (_04717_, _04716_, _04714_);
  and (_04718_, _04717_, _04556_);
  or (_04719_, _04718_, _04094_);
  and (_04720_, _01968_, _01621_);
  nor (_04721_, _04715_, _04094_);
  or (_04722_, _04721_, _02803_);
  and (_04723_, _04722_, _04720_);
  and (_04724_, _04723_, _04719_);
  nor (_04725_, _02858_, _01629_);
  nor (_04726_, _04720_, _02855_);
  or (_04727_, _04726_, _04725_);
  or (_04728_, _04727_, _04724_);
  not (_04729_, _04725_);
  or (_04730_, _04729_, _02803_);
  and (_04731_, _04730_, _01964_);
  and (_04732_, _04731_, _04728_);
  or (_04733_, _04732_, _04092_);
  nor (_04734_, _04093_, _01629_);
  not (_04735_, _04734_);
  and (_04736_, _04735_, _04733_);
  and (_04737_, _04734_, _02803_);
  and (_04738_, _02455_, _01630_);
  not (_04739_, _04738_);
  or (_04740_, _04739_, _04737_);
  or (_04741_, _04740_, _04736_);
  or (_04742_, _04738_, _02851_);
  and (_04743_, _04742_, _04741_);
  or (_04744_, _04743_, _04089_);
  and (_04745_, _04744_, _04091_);
  or (_04746_, _04745_, _03185_);
  and (_04747_, _04746_, _03913_);
  or (_04748_, _04747_, _01951_);
  not (_04749_, _03179_);
  and (_04750_, _04191_, \oc8051_golden_model_1.P2INREG [1]);
  and (_04751_, _04197_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_04752_, _04751_, _04750_);
  and (_04753_, _04194_, \oc8051_golden_model_1.P1INREG [1]);
  and (_04754_, _04387_, \oc8051_golden_model_1.P0INREG [1]);
  nor (_04755_, _04754_, _04753_);
  and (_04756_, _04755_, _04752_);
  and (_04757_, _04756_, _04442_);
  and (_04758_, _04757_, _04435_);
  and (_04759_, _04758_, _04406_);
  nor (_04760_, _04759_, \oc8051_golden_model_1.ACC [1]);
  and (_04761_, _04759_, \oc8051_golden_model_1.ACC [1]);
  nor (_04762_, _04761_, _04760_);
  not (_04763_, _04511_);
  and (_04764_, _04520_, _04763_);
  nor (_04765_, _04512_, _04514_);
  and (_04766_, _04765_, _04764_);
  and (_04767_, _04197_, \oc8051_golden_model_1.P3INREG [7]);
  and (_04768_, _04191_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_04769_, _04768_, _04767_);
  and (_04770_, _04194_, \oc8051_golden_model_1.P1INREG [7]);
  and (_04771_, _04387_, \oc8051_golden_model_1.P0INREG [7]);
  nor (_04772_, _04771_, _04770_);
  and (_04773_, _04772_, _04769_);
  and (_04774_, _04773_, _04766_);
  and (_04775_, _04531_, _04523_);
  and (_04776_, _04775_, _04543_);
  and (_04777_, _04776_, _04510_);
  and (_04778_, _04777_, _04774_);
  and (_04779_, _04778_, _04079_);
  nor (_04780_, _04779_, \oc8051_golden_model_1.ACC [7]);
  and (_04781_, _04779_, \oc8051_golden_model_1.ACC [7]);
  nor (_04782_, _04781_, _04780_);
  and (_04783_, _04782_, _04762_);
  and (_04784_, _04191_, \oc8051_golden_model_1.P2INREG [2]);
  and (_04785_, _04197_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_04786_, _04785_, _04784_);
  and (_04787_, _04194_, \oc8051_golden_model_1.P1INREG [2]);
  and (_04788_, _04387_, \oc8051_golden_model_1.P0INREG [2]);
  nor (_04789_, _04788_, _04787_);
  and (_04790_, _04789_, _04786_);
  and (_04791_, _04790_, _04240_);
  and (_04792_, _04791_, _04234_);
  and (_04793_, _04792_, _04205_);
  nor (_04794_, _04793_, \oc8051_golden_model_1.ACC [2]);
  and (_04795_, _04793_, \oc8051_golden_model_1.ACC [2]);
  nor (_04796_, _04795_, _04794_);
  and (_04797_, _04191_, \oc8051_golden_model_1.P2INREG [6]);
  and (_04798_, _04197_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_04799_, _04798_, _04797_);
  and (_04800_, _04194_, \oc8051_golden_model_1.P1INREG [6]);
  and (_04801_, _04387_, \oc8051_golden_model_1.P0INREG [6]);
  nor (_04802_, _04801_, _04800_);
  and (_04803_, _04802_, _04799_);
  and (_04804_, _04803_, _04489_);
  and (_04805_, _04804_, _04483_);
  and (_04806_, _04805_, _04454_);
  nor (_04807_, _04806_, \oc8051_golden_model_1.ACC [6]);
  and (_04808_, _04806_, \oc8051_golden_model_1.ACC [6]);
  nor (_04809_, _04808_, _04807_);
  and (_04810_, _04809_, _04796_);
  and (_04811_, _04810_, _04783_);
  and (_04812_, _04197_, \oc8051_golden_model_1.P3INREG [0]);
  and (_04813_, _04191_, \oc8051_golden_model_1.P2INREG [0]);
  nor (_04814_, _04813_, _04812_);
  and (_04815_, _04194_, \oc8051_golden_model_1.P1INREG [0]);
  and (_04816_, _04387_, \oc8051_golden_model_1.P0INREG [0]);
  nor (_04817_, _04816_, _04815_);
  and (_04818_, _04817_, _04814_);
  not (_04819_, _04370_);
  and (_04820_, _04379_, _04819_);
  nor (_04821_, _04371_, _04373_);
  and (_04822_, _04821_, _04820_);
  and (_04823_, _04822_, _04818_);
  and (_04824_, _04382_, _04359_);
  and (_04825_, _04824_, _04402_);
  and (_04826_, _04825_, _04369_);
  and (_04827_, _04826_, _04823_);
  and (_04828_, _04827_, _04350_);
  nor (_04829_, _04828_, \oc8051_golden_model_1.ACC [0]);
  and (_04830_, _04828_, \oc8051_golden_model_1.ACC [0]);
  nor (_04831_, _04830_, _04829_);
  and (_04832_, _04191_, \oc8051_golden_model_1.P2INREG [4]);
  and (_04833_, _04197_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_04834_, _04833_, _04832_);
  and (_04835_, _04194_, \oc8051_golden_model_1.P1INREG [4]);
  and (_04836_, _04387_, \oc8051_golden_model_1.P0INREG [4]);
  nor (_04837_, _04836_, _04835_);
  and (_04838_, _04837_, _04834_);
  and (_04839_, _04838_, _04287_);
  and (_04840_, _04839_, _04277_);
  and (_04841_, _04840_, _04254_);
  nor (_04842_, _04841_, \oc8051_golden_model_1.ACC [4]);
  and (_04843_, _04841_, \oc8051_golden_model_1.ACC [4]);
  nor (_04844_, _04843_, _04842_);
  and (_04845_, _04844_, _04831_);
  and (_04846_, _04191_, \oc8051_golden_model_1.P2INREG [3]);
  and (_04847_, _04197_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_04848_, _04847_, _04846_);
  and (_04849_, _04194_, \oc8051_golden_model_1.P1INREG [3]);
  and (_04850_, _04387_, \oc8051_golden_model_1.P0INREG [3]);
  nor (_04851_, _04850_, _04849_);
  and (_04852_, _04851_, _04848_);
  and (_04853_, _04852_, _04187_);
  and (_04854_, _04853_, _04152_);
  and (_04855_, _04854_, _04095_);
  nor (_04856_, _04855_, \oc8051_golden_model_1.ACC [3]);
  and (_04857_, _04855_, \oc8051_golden_model_1.ACC [3]);
  nor (_04858_, _04857_, _04856_);
  and (_04859_, _04191_, \oc8051_golden_model_1.P2INREG [5]);
  and (_04860_, _04197_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_04861_, _04860_, _04859_);
  and (_04862_, _04194_, \oc8051_golden_model_1.P1INREG [5]);
  and (_04863_, _04387_, \oc8051_golden_model_1.P0INREG [5]);
  nor (_04864_, _04863_, _04862_);
  and (_04865_, _04864_, _04861_);
  and (_04866_, _04865_, _04335_);
  and (_04867_, _04866_, _04321_);
  and (_04868_, _04867_, _04300_);
  nor (_04869_, _04868_, \oc8051_golden_model_1.ACC [5]);
  and (_04870_, _04868_, \oc8051_golden_model_1.ACC [5]);
  nor (_04871_, _04870_, _04869_);
  and (_04872_, _04871_, _04858_);
  and (_04873_, _04872_, _04845_);
  and (_04874_, _04873_, _04811_);
  not (_04875_, _04874_);
  and (_04876_, _04875_, _03176_);
  and (_04877_, _04874_, _02878_);
  or (_04878_, _04877_, _02378_);
  or (_04879_, _04878_, _04876_);
  and (_04880_, _04879_, _04749_);
  and (_04881_, _04880_, _04748_);
  or (_04882_, _04881_, _03184_);
  and (_04883_, _04882_, _02881_);
  nand (_04884_, _02880_, _02803_);
  not (_04885_, _01946_);
  and (_04886_, _02003_, _01937_);
  and (_04887_, _04886_, _01929_);
  and (_04888_, _02035_, _01929_);
  nor (_04889_, _04888_, _04887_);
  not (_04890_, _02032_);
  and (_04891_, _02008_, _04890_);
  nor (_04892_, _04891_, _01617_);
  nor (_04893_, _04892_, _01945_);
  and (_04894_, _04893_, _04889_);
  and (_04895_, _02004_, _01929_);
  nor (_04896_, _04895_, _03273_);
  and (_04897_, _04896_, _04894_);
  and (_04898_, _04897_, _01632_);
  and (_04899_, _04898_, _04885_);
  nand (_04900_, _04899_, _04884_);
  or (_04901_, _04900_, _04883_);
  or (_04902_, _04899_, _02851_);
  and (_04903_, _01929_, _01593_);
  nor (_04904_, _04093_, _01617_);
  nor (_04905_, _04904_, _04903_);
  and (_04906_, _04905_, _04902_);
  and (_04907_, _04906_, _04901_);
  not (_04908_, _04905_);
  and (_04909_, _04908_, _02803_);
  and (_04910_, _01932_, _01618_);
  not (_04911_, _04910_);
  or (_04912_, _04911_, _04909_);
  or (_04913_, _04912_, _04907_);
  and (_04914_, _02010_, _01605_);
  and (_04915_, _02804_, _01605_);
  or (_04916_, _04915_, _04914_);
  not (_04917_, _04916_);
  not (_04918_, _01927_);
  nor (_04919_, _01939_, _01609_);
  and (_04920_, _04919_, _01605_);
  and (_04921_, _04920_, _04918_);
  not (_04922_, _04921_);
  and (_04923_, _02413_, _01605_);
  or (_04924_, _02006_, _01934_);
  and (_04925_, _04924_, _01605_);
  nor (_04926_, _04925_, _04923_);
  and (_04927_, _04926_, _04922_);
  and (_04928_, _04927_, _04917_);
  or (_04929_, _04910_, _02851_);
  and (_04930_, _04929_, _04928_);
  and (_04931_, _04930_, _04913_);
  and (_04932_, _01605_, _02272_);
  not (_04933_, _04928_);
  and (_04934_, _04933_, _02803_);
  or (_04935_, _04934_, _04932_);
  or (_04936_, _04935_, _04931_);
  not (_04937_, _04932_);
  or (_04938_, _02851_, _04937_);
  and (_04939_, _04938_, _01616_);
  and (_04940_, _04939_, _04936_);
  and (_04941_, _02803_, _01611_);
  nor (_04942_, _01924_, _01606_);
  not (_04943_, _04942_);
  or (_04944_, _04943_, _04941_);
  or (_04945_, _04944_, _04940_);
  or (_04946_, _04942_, _02851_);
  and (_04947_, _04946_, _02002_);
  and (_04948_, _04947_, _04945_);
  and (_04949_, _02878_, _02001_);
  and (_04950_, _01601_, _01382_);
  and (_04951_, _02857_, _01601_);
  nor (_04952_, _04951_, _04950_);
  not (_04953_, _04952_);
  or (_04954_, _04953_, _04949_);
  or (_04955_, _04954_, _04948_);
  or (_04956_, _04952_, _02851_);
  and (_04957_, _04956_, _01923_);
  and (_04958_, _04957_, _04955_);
  or (_04959_, _04958_, _02879_);
  nor (_04960_, _04093_, _02339_);
  not (_04961_, _04960_);
  and (_04962_, _04961_, _04959_);
  nor (_04963_, _01920_, _01654_);
  not (_04964_, _04963_);
  and (_04965_, _04960_, _02803_);
  or (_04966_, _04965_, _04964_);
  or (_04967_, _04966_, _04962_);
  and (_04968_, _01601_, _01928_);
  not (_04969_, _04968_);
  or (_04970_, _04963_, _02851_);
  and (_04971_, _04970_, _04969_);
  and (_04972_, _04971_, _04967_);
  and (_04973_, _04968_, _04700_);
  or (_04974_, _02859_, _04973_);
  or (_04975_, _04974_, _04972_);
  and (_04976_, _04975_, _02860_);
  or (_04977_, _04976_, _02019_);
  not (_04978_, _02853_);
  not (_04979_, _02019_);
  or (_04980_, _02878_, _04979_);
  and (_04981_, _04980_, _04978_);
  and (_04982_, _04981_, _04977_);
  or (_04983_, _04982_, _02854_);
  and (_04984_, _01649_, _01610_);
  not (_04985_, _04984_);
  and (_04986_, _04985_, _04983_);
  not (_04987_, \oc8051_golden_model_1.DPH [7]);
  and (_04988_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_04989_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_04990_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_04991_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_04992_, _04991_, _04990_);
  not (_04993_, _04992_);
  and (_04994_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_04995_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_04996_, _04995_, _04994_);
  not (_04997_, _04996_);
  and (_04998_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_04999_, _01755_, _01751_);
  nor (_05000_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_05001_, _05000_, _04998_);
  not (_05002_, _05001_);
  nor (_05003_, _05002_, _04999_);
  nor (_05004_, _05003_, _04998_);
  nor (_05005_, _05004_, _04997_);
  nor (_05006_, _05005_, _04994_);
  nor (_05007_, _05006_, _04993_);
  nor (_05008_, _05007_, _04990_);
  nor (_05009_, _05008_, _04989_);
  or (_05010_, _05009_, _04988_);
  and (_05011_, _05010_, \oc8051_golden_model_1.DPH [0]);
  and (_05012_, _05011_, \oc8051_golden_model_1.DPH [1]);
  and (_05013_, _05012_, \oc8051_golden_model_1.DPH [2]);
  and (_05014_, _05013_, \oc8051_golden_model_1.DPH [3]);
  and (_05015_, _05014_, \oc8051_golden_model_1.DPH [4]);
  and (_05016_, _05015_, \oc8051_golden_model_1.DPH [5]);
  and (_05017_, _05016_, \oc8051_golden_model_1.DPH [6]);
  nor (_05018_, _05017_, _04987_);
  and (_05019_, _05017_, _04987_);
  or (_05020_, _05019_, _05018_);
  and (_05021_, _05020_, _04984_);
  nor (_05022_, _01919_, _01650_);
  not (_05023_, _05022_);
  or (_05024_, _05023_, _05021_);
  or (_05025_, _05024_, _04986_);
  and (_05026_, _01649_, _01928_);
  not (_05027_, _05026_);
  or (_05028_, _05022_, _02851_);
  and (_05029_, _05028_, _05027_);
  and (_05030_, _05029_, _05025_);
  not (_05031_, _02830_);
  nor (_05032_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_05033_, \oc8051_golden_model_1.ACC [6], \oc8051_golden_model_1.ACC [3]);
  and (_05034_, _05033_, _05032_);
  nor (_05035_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [7]);
  nor (_05036_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  and (_05037_, _05036_, _05035_);
  and (_05038_, _05037_, _05034_);
  or (_05039_, _05038_, _04700_);
  not (_05040_, _05038_);
  or (_05041_, _05040_, _02851_);
  and (_05042_, _05041_, _05026_);
  and (_05043_, _05042_, _05039_);
  or (_05044_, _05043_, _05031_);
  or (_05045_, _05044_, _05030_);
  and (_05046_, _05045_, _02831_);
  and (_05047_, _01652_, _02272_);
  or (_05048_, _05047_, _05046_);
  not (_05049_, _02018_);
  not (_05050_, _05047_);
  or (_05051_, _05050_, _02851_);
  and (_05052_, _05051_, _05049_);
  and (_05053_, _05052_, _05048_);
  and (_05054_, _02878_, _02018_);
  nor (_05055_, _02135_, _01653_);
  not (_05056_, _05055_);
  or (_05057_, _05056_, _05054_);
  or (_05058_, _05057_, _05053_);
  and (_05059_, _01652_, _01928_);
  not (_05060_, _05059_);
  or (_05061_, _05055_, _02851_);
  and (_05062_, _05061_, _05060_);
  and (_05063_, _05062_, _05058_);
  or (_05064_, _05040_, _04700_);
  or (_05065_, _05038_, _02851_);
  and (_05066_, _05065_, _05059_);
  and (_05067_, _05066_, _05064_);
  or (_05068_, _05067_, _05063_);
  nor (_05069_, _02858_, _02531_);
  not (_05070_, _05069_);
  and (_05071_, _05070_, _05068_);
  and (_05072_, _01665_, _02272_);
  and (_05073_, _05069_, _02803_);
  or (_05074_, _05073_, _05072_);
  or (_05075_, _05074_, _05071_);
  not (_05076_, _02039_);
  not (_05077_, _05072_);
  or (_05078_, _02851_, _05077_);
  and (_05079_, _05078_, _05076_);
  and (_05080_, _05079_, _05075_);
  and (_05081_, _02878_, _02039_);
  nor (_05082_, _02130_, _01666_);
  not (_05083_, _05082_);
  or (_05084_, _05083_, _05081_);
  or (_05085_, _05084_, _05080_);
  and (_05086_, _01665_, _01928_);
  not (_05087_, _05086_);
  or (_05088_, _05082_, _02851_);
  and (_05089_, _05088_, _05087_);
  and (_05090_, _05089_, _05085_);
  or (_05091_, _04700_, \oc8051_golden_model_1.PSW [7]);
  not (_05092_, \oc8051_golden_model_1.PSW [7]);
  or (_05093_, _02851_, _05092_);
  and (_05094_, _05093_, _05086_);
  and (_05095_, _05094_, _05091_);
  or (_05096_, _05095_, _05090_);
  nor (_05097_, _02858_, _02536_);
  not (_05098_, _05097_);
  and (_05099_, _05098_, _05096_);
  and (_05100_, _05097_, _02803_);
  and (_05101_, _01662_, _02272_);
  or (_05102_, _05101_, _05100_);
  or (_05103_, _05102_, _05099_);
  not (_05104_, _02016_);
  not (_05105_, _05101_);
  or (_05106_, _05105_, _02851_);
  and (_05107_, _05106_, _05104_);
  and (_05108_, _05107_, _05103_);
  and (_05109_, _02878_, _02016_);
  nor (_05110_, _02126_, _01663_);
  not (_05111_, _05110_);
  or (_05112_, _05111_, _05109_);
  or (_05113_, _05112_, _05108_);
  and (_05114_, _01662_, _01928_);
  not (_05115_, _05114_);
  or (_05116_, _05110_, _02851_);
  and (_05117_, _05116_, _05115_);
  and (_05118_, _05117_, _05113_);
  or (_05119_, _04700_, _05092_);
  or (_05120_, _02851_, \oc8051_golden_model_1.PSW [7]);
  and (_05121_, _05120_, _05114_);
  and (_05122_, _05121_, _05119_);
  or (_05123_, _05122_, _05118_);
  and (_05124_, _02413_, _01659_);
  not (_05125_, _05124_);
  and (_05126_, _02321_, _01659_);
  nor (_05127_, _02681_, _05126_);
  and (_05128_, _05127_, _05125_);
  and (_05129_, _02804_, _01659_);
  nor (_05130_, _05129_, _02362_);
  and (_05131_, _02006_, _01659_);
  and (_05132_, _02030_, _01659_);
  nor (_05133_, _05132_, _05131_);
  and (_05134_, _05133_, _05130_);
  and (_05135_, _02325_, _01659_);
  and (_05136_, _02010_, _01659_);
  nor (_05137_, _05136_, _05135_);
  and (_05138_, _05137_, _05134_);
  and (_05139_, _05138_, _05128_);
  and (_05140_, _05139_, _05123_);
  not (_05141_, _05139_);
  and (_05142_, _05141_, _02803_);
  or (_05143_, _05142_, _02273_);
  or (_05144_, _05143_, _05140_);
  and (_05145_, _01659_, _01610_);
  not (_05146_, _05145_);
  not (_05147_, _02273_);
  or (_05148_, _02851_, _05147_);
  and (_05149_, _05148_, _05146_);
  and (_05150_, _05149_, _05144_);
  and (_05151_, _05145_, _02803_);
  or (_05152_, _05151_, _02146_);
  or (_05153_, _05152_, _05150_);
  nand (_05154_, _02786_, _02146_);
  and (_05155_, _05154_, _05153_);
  or (_05156_, _05155_, _01660_);
  not (_05157_, _01660_);
  or (_05158_, _02851_, _05157_);
  and (_05159_, _05158_, _02153_);
  and (_05160_, _05159_, _05156_);
  not (_05161_, _02818_);
  not (_05162_, _04106_);
  nor (_05163_, _02610_, _02450_);
  not (_05164_, _02221_);
  and (_05165_, _05164_, _01918_);
  and (_05166_, _05165_, _05163_);
  and (_05167_, _05166_, _04098_);
  and (_05168_, _05167_, \oc8051_golden_model_1.TCON [2]);
  nor (_05169_, _02221_, _01918_);
  and (_05170_, _05169_, _05163_);
  and (_05171_, _04170_, _05170_);
  and (_05172_, _05171_, \oc8051_golden_model_1.B [2]);
  nor (_05173_, _05172_, _05168_);
  and (_05174_, _05166_, _04154_);
  and (_05175_, _05174_, \oc8051_golden_model_1.IP [2]);
  not (_05176_, _05175_);
  and (_05177_, _04166_, _05170_);
  and (_05178_, _05177_, \oc8051_golden_model_1.PSW [2]);
  and (_05179_, _04161_, _05170_);
  and (_05180_, _05179_, \oc8051_golden_model_1.ACC [2]);
  nor (_05181_, _05180_, _05178_);
  and (_05182_, _05181_, _05176_);
  and (_05183_, _05182_, _05173_);
  and (_05184_, _05166_, _04128_);
  and (_05185_, _05184_, \oc8051_golden_model_1.SCON [2]);
  and (_05186_, _05166_, _04182_);
  and (_05187_, _05186_, \oc8051_golden_model_1.IE [2]);
  nor (_05188_, _05187_, _05185_);
  and (_05189_, _04182_, _05170_);
  and (_05190_, _05189_, \oc8051_golden_model_1.P2INREG [2]);
  and (_05191_, _04154_, _05170_);
  and (_05192_, _05191_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_05193_, _05192_, _05190_);
  and (_05194_, _04099_, \oc8051_golden_model_1.P0INREG [2]);
  and (_05195_, _04128_, _05170_);
  and (_05196_, _05195_, \oc8051_golden_model_1.P1INREG [2]);
  nor (_05197_, _05196_, _05194_);
  and (_05198_, _05197_, _05193_);
  and (_05199_, _05198_, _05188_);
  and (_05200_, _05199_, _05183_);
  and (_05201_, _05200_, _04205_);
  nor (_05202_, _05201_, _05162_);
  not (_05203_, _04110_);
  and (_05204_, _05167_, \oc8051_golden_model_1.TCON [1]);
  and (_05205_, _05179_, \oc8051_golden_model_1.ACC [1]);
  nor (_05206_, _05205_, _05204_);
  and (_05207_, _05177_, \oc8051_golden_model_1.PSW [1]);
  not (_05208_, _05207_);
  and (_05209_, _05174_, \oc8051_golden_model_1.IP [1]);
  and (_05210_, _05171_, \oc8051_golden_model_1.B [1]);
  nor (_05211_, _05210_, _05209_);
  and (_05212_, _05211_, _05208_);
  and (_05213_, _05212_, _05206_);
  and (_05214_, _05184_, \oc8051_golden_model_1.SCON [1]);
  and (_05215_, _05186_, \oc8051_golden_model_1.IE [1]);
  nor (_05216_, _05215_, _05214_);
  and (_05217_, _05189_, \oc8051_golden_model_1.P2INREG [1]);
  and (_05218_, _05191_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_05219_, _05218_, _05217_);
  and (_05220_, _04099_, \oc8051_golden_model_1.P0INREG [1]);
  and (_05221_, _05195_, \oc8051_golden_model_1.P1INREG [1]);
  nor (_05222_, _05221_, _05220_);
  and (_05223_, _05222_, _05219_);
  and (_05224_, _05223_, _05216_);
  and (_05225_, _05224_, _05213_);
  and (_05226_, _05225_, _04406_);
  nor (_05227_, _05226_, _05203_);
  nor (_05228_, _05227_, _05202_);
  and (_05229_, _05167_, \oc8051_golden_model_1.TCON [4]);
  and (_05230_, _05171_, \oc8051_golden_model_1.B [4]);
  nor (_05231_, _05230_, _05229_);
  and (_05232_, _05174_, \oc8051_golden_model_1.IP [4]);
  not (_05233_, _05232_);
  and (_05234_, _05177_, \oc8051_golden_model_1.PSW [4]);
  and (_05235_, _05179_, \oc8051_golden_model_1.ACC [4]);
  nor (_05236_, _05235_, _05234_);
  and (_05237_, _05236_, _05233_);
  and (_05238_, _05237_, _05231_);
  and (_05239_, _05184_, \oc8051_golden_model_1.SCON [4]);
  and (_05240_, _05186_, \oc8051_golden_model_1.IE [4]);
  nor (_05241_, _05240_, _05239_);
  and (_05242_, _05189_, \oc8051_golden_model_1.P2INREG [4]);
  and (_05243_, _05191_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_05244_, _05243_, _05242_);
  and (_05245_, _04099_, \oc8051_golden_model_1.P0INREG [4]);
  and (_05246_, _05195_, \oc8051_golden_model_1.P1INREG [4]);
  nor (_05247_, _05246_, _05245_);
  and (_05248_, _05247_, _05244_);
  and (_05249_, _05248_, _05241_);
  and (_05250_, _05249_, _05238_);
  and (_05251_, _05250_, _04254_);
  and (_05252_, _04115_, _02264_);
  not (_05253_, _05252_);
  nor (_05254_, _05253_, _05251_);
  not (_05255_, _04176_);
  and (_05256_, _05167_, \oc8051_golden_model_1.TCON [7]);
  and (_05257_, _05179_, \oc8051_golden_model_1.ACC [7]);
  nor (_05258_, _05257_, _05256_);
  and (_05259_, _05174_, \oc8051_golden_model_1.IP [7]);
  not (_05260_, _05259_);
  and (_05261_, _05177_, \oc8051_golden_model_1.PSW [7]);
  and (_05262_, _05171_, \oc8051_golden_model_1.B [7]);
  nor (_05263_, _05262_, _05261_);
  and (_05264_, _05263_, _05260_);
  and (_05265_, _05264_, _05258_);
  and (_05266_, _05184_, \oc8051_golden_model_1.SCON [7]);
  and (_05267_, _05186_, \oc8051_golden_model_1.IE [7]);
  nor (_05268_, _05267_, _05266_);
  and (_05269_, _05189_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05270_, _05191_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05271_, _05270_, _05269_);
  and (_05272_, _04099_, \oc8051_golden_model_1.P0INREG [7]);
  and (_05273_, _05195_, \oc8051_golden_model_1.P1INREG [7]);
  nor (_05274_, _05273_, _05272_);
  and (_05275_, _05274_, _05271_);
  and (_05276_, _05275_, _05268_);
  and (_05277_, _05276_, _05265_);
  and (_05278_, _05277_, _04079_);
  nor (_05279_, _05278_, _05255_);
  nor (_05280_, _05279_, _05254_);
  and (_05281_, _05280_, _05228_);
  not (_05282_, _04157_);
  and (_05283_, _05195_, \oc8051_golden_model_1.P1INREG [0]);
  and (_05284_, _04099_, \oc8051_golden_model_1.P0INREG [0]);
  nor (_05285_, _05284_, _05283_);
  and (_05286_, _05184_, \oc8051_golden_model_1.SCON [0]);
  and (_05287_, _05186_, \oc8051_golden_model_1.IE [0]);
  nor (_05288_, _05287_, _05286_);
  and (_05289_, _05174_, \oc8051_golden_model_1.IP [0]);
  and (_05290_, _05171_, \oc8051_golden_model_1.B [0]);
  nor (_05291_, _05290_, _05289_);
  and (_05292_, _05177_, \oc8051_golden_model_1.PSW [0]);
  and (_05293_, _05179_, \oc8051_golden_model_1.ACC [0]);
  nor (_05294_, _05293_, _05292_);
  and (_05295_, _05294_, _05291_);
  and (_05296_, _05167_, \oc8051_golden_model_1.TCON [0]);
  and (_05297_, _05191_, \oc8051_golden_model_1.P3INREG [0]);
  and (_05298_, _05189_, \oc8051_golden_model_1.P2INREG [0]);
  or (_05299_, _05298_, _05297_);
  nor (_05300_, _05299_, _05296_);
  and (_05301_, _05300_, _05295_);
  and (_05302_, _05301_, _05288_);
  and (_05303_, _05302_, _05285_);
  and (_05304_, _05303_, _04350_);
  nor (_05305_, _05304_, _05282_);
  and (_05306_, _05167_, \oc8051_golden_model_1.TCON [6]);
  and (_05307_, _05179_, \oc8051_golden_model_1.ACC [6]);
  nor (_05308_, _05307_, _05306_);
  and (_05309_, _05177_, \oc8051_golden_model_1.PSW [6]);
  not (_05310_, _05309_);
  and (_05311_, _05174_, \oc8051_golden_model_1.IP [6]);
  and (_05312_, _05171_, \oc8051_golden_model_1.B [6]);
  nor (_05313_, _05312_, _05311_);
  and (_05314_, _05313_, _05310_);
  and (_05315_, _05314_, _05308_);
  and (_05316_, _05184_, \oc8051_golden_model_1.SCON [6]);
  and (_05317_, _05186_, \oc8051_golden_model_1.IE [6]);
  nor (_05318_, _05317_, _05316_);
  and (_05319_, _05189_, \oc8051_golden_model_1.P2INREG [6]);
  and (_05320_, _05191_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_05321_, _05320_, _05319_);
  and (_05322_, _04099_, \oc8051_golden_model_1.P0INREG [6]);
  and (_05324_, _05195_, \oc8051_golden_model_1.P1INREG [6]);
  nor (_05325_, _05324_, _05322_);
  and (_05326_, _05325_, _05321_);
  and (_05327_, _05326_, _05318_);
  and (_05328_, _05327_, _05315_);
  and (_05329_, _05328_, _04454_);
  and (_05330_, _04105_, _02264_);
  not (_05331_, _05330_);
  nor (_05332_, _05331_, _05329_);
  nor (_05333_, _05332_, _05305_);
  not (_05334_, _04101_);
  and (_05335_, _05177_, \oc8051_golden_model_1.PSW [3]);
  and (_05336_, _05179_, \oc8051_golden_model_1.ACC [3]);
  nor (_05337_, _05336_, _05335_);
  and (_05338_, _05174_, \oc8051_golden_model_1.IP [3]);
  and (_05339_, _05171_, \oc8051_golden_model_1.B [3]);
  nor (_05340_, _05339_, _05338_);
  and (_05341_, _05340_, _05337_);
  and (_05342_, _05167_, \oc8051_golden_model_1.TCON [3]);
  not (_05343_, _05342_);
  and (_05344_, _05189_, \oc8051_golden_model_1.P2INREG [3]);
  and (_05345_, _05191_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_05346_, _05345_, _05344_);
  and (_05347_, _05346_, _05343_);
  and (_05348_, _05184_, \oc8051_golden_model_1.SCON [3]);
  and (_05349_, _05186_, \oc8051_golden_model_1.IE [3]);
  nor (_05350_, _05349_, _05348_);
  and (_05351_, _04099_, \oc8051_golden_model_1.P0INREG [3]);
  and (_05352_, _05195_, \oc8051_golden_model_1.P1INREG [3]);
  nor (_05353_, _05352_, _05351_);
  and (_05354_, _05353_, _05350_);
  and (_05355_, _05354_, _05347_);
  and (_05356_, _05355_, _05341_);
  and (_05357_, _05356_, _04095_);
  nor (_05358_, _05357_, _05334_);
  and (_05359_, _05195_, \oc8051_golden_model_1.P1INREG [5]);
  and (_05360_, _04099_, \oc8051_golden_model_1.P0INREG [5]);
  nor (_05361_, _05360_, _05359_);
  and (_05362_, _05184_, \oc8051_golden_model_1.SCON [5]);
  and (_05363_, _05186_, \oc8051_golden_model_1.IE [5]);
  nor (_05364_, _05363_, _05362_);
  and (_05365_, _05174_, \oc8051_golden_model_1.IP [5]);
  and (_05366_, _05171_, \oc8051_golden_model_1.B [5]);
  nor (_05367_, _05366_, _05365_);
  and (_05368_, _05177_, \oc8051_golden_model_1.PSW [5]);
  and (_05369_, _05179_, \oc8051_golden_model_1.ACC [5]);
  nor (_05370_, _05369_, _05368_);
  and (_05371_, _05370_, _05367_);
  and (_05372_, _05167_, \oc8051_golden_model_1.TCON [5]);
  and (_05373_, _05191_, \oc8051_golden_model_1.P3INREG [5]);
  and (_05374_, _05189_, \oc8051_golden_model_1.P2INREG [5]);
  or (_05375_, _05374_, _05373_);
  nor (_05376_, _05375_, _05372_);
  and (_05377_, _05376_, _05371_);
  and (_05378_, _05377_, _05364_);
  and (_05379_, _05378_, _05361_);
  and (_05380_, _05379_, _04300_);
  and (_05381_, _04109_, _02264_);
  not (_05382_, _05381_);
  nor (_05383_, _05382_, _05380_);
  nor (_05384_, _05383_, _05358_);
  and (_05385_, _05384_, _05333_);
  and (_05386_, _05385_, _05281_);
  not (_05387_, _05386_);
  or (_05388_, _05387_, _03176_);
  or (_05389_, _05386_, _02878_);
  and (_05390_, _05389_, _02015_);
  and (_05391_, _05390_, _05388_);
  or (_05392_, _05391_, _05161_);
  or (_05393_, _05392_, _05160_);
  and (_05394_, _05393_, _02819_);
  or (_05395_, _05394_, _02788_);
  and (_05396_, _01610_, _01580_);
  not (_05397_, _05396_);
  not (_05398_, _02788_);
  or (_05399_, _02851_, _05398_);
  and (_05400_, _05399_, _05397_);
  and (_05401_, _05400_, _05395_);
  and (_05402_, _05396_, _02803_);
  or (_05403_, _05402_, _01585_);
  or (_05404_, _05403_, _05401_);
  and (_05405_, _05404_, _02787_);
  or (_05406_, _05405_, _01581_);
  not (_05407_, _01581_);
  or (_05408_, _02851_, _05407_);
  and (_05409_, _05408_, _02558_);
  and (_05410_, _05409_, _05406_);
  or (_05411_, _05386_, _03176_);
  nand (_05412_, _05386_, _03168_);
  and (_05413_, _05412_, _05411_);
  and (_05414_, _05413_, _02022_);
  nand (_05415_, _01669_, _01382_);
  not (_05416_, _05415_);
  and (_05417_, _02857_, _01669_);
  nor (_05418_, _05417_, _05416_);
  not (_05419_, _05418_);
  or (_05420_, _05419_, _05414_);
  or (_05421_, _05420_, _05410_);
  or (_05422_, _05418_, _02803_);
  and (_05423_, _05422_, _02168_);
  and (_05424_, _05423_, _05421_);
  and (_05425_, _02851_, _02164_);
  nor (_05426_, _04093_, _02560_);
  or (_05427_, _05426_, _05425_);
  or (_05428_, _05427_, _05424_);
  not (_05429_, _02023_);
  not (_05430_, _05426_);
  or (_05431_, _05430_, _02803_);
  and (_05432_, _05431_, _05429_);
  and (_05433_, _05432_, _05428_);
  nor (_05434_, _05429_, _01853_);
  or (_05435_, _05434_, _01670_);
  or (_05436_, _05435_, _05433_);
  or (_05437_, _02851_, _01671_);
  and (_05438_, _05437_, _02377_);
  and (_05439_, _05438_, _05436_);
  and (_05440_, _05413_, _02025_);
  and (_05441_, _02857_, _01589_);
  not (_05442_, _05441_);
  and (_05443_, _01938_, _01589_);
  nor (_05444_, _05443_, _02359_);
  and (_05445_, _05444_, _05442_);
  not (_05446_, _05445_);
  or (_05447_, _05446_, _05440_);
  or (_05448_, _05447_, _05439_);
  or (_05449_, _05445_, _02803_);
  and (_05450_, _05449_, _01595_);
  and (_05451_, _05450_, _05448_);
  and (_05452_, _02851_, _01594_);
  nor (_05453_, _04093_, _02569_);
  or (_05454_, _05453_, _05452_);
  or (_05455_, _05454_, _05451_);
  not (_05456_, _02026_);
  not (_05457_, _05453_);
  or (_05458_, _05457_, _02803_);
  and (_05459_, _05458_, _05456_);
  and (_05460_, _05459_, _05455_);
  nor (_05461_, _05456_, _01853_);
  or (_05462_, _05461_, _01657_);
  or (_05463_, _05462_, _05460_);
  and (_05464_, _01928_, _01589_);
  not (_05465_, _05464_);
  or (_05466_, _02851_, _01658_);
  and (_05467_, _05466_, _05465_);
  and (_05468_, _05467_, _05463_);
  and (_05469_, _02803_, _05464_);
  or (_05470_, _05469_, _05468_);
  or (_05471_, _05470_, _26506_);
  or (_05472_, _26505_, \oc8051_golden_model_1.PC [15]);
  and (_05473_, _05472_, _25964_);
  and (_25309_, _05473_, _05471_);
  not (_05474_, _02126_);
  not (_05475_, \oc8051_golden_model_1.TMOD [7]);
  nor (_05476_, _04134_, _05475_);
  and (_05477_, _04134_, _02962_);
  nor (_05478_, _05477_, _05476_);
  and (_05479_, _05478_, _02019_);
  not (_05480_, _04134_);
  nor (_05481_, _05480_, _02786_);
  nor (_05482_, _05481_, _05476_);
  and (_05483_, _05482_, _04950_);
  and (_05484_, _04134_, \oc8051_golden_model_1.ACC [7]);
  nor (_05485_, _05484_, _05476_);
  nor (_05486_, _05485_, _01964_);
  not (_05487_, _01967_);
  not (_05488_, _04571_);
  nor (_05489_, _05485_, _05488_);
  nor (_05490_, _04571_, _05475_);
  or (_05491_, _05490_, _05489_);
  and (_05492_, _05491_, _02438_);
  not (_05493_, _04405_);
  and (_05494_, _04452_, _05493_);
  and (_05495_, _05494_, _04349_);
  and (_05496_, _05495_, _04501_);
  nor (_05497_, _05496_, _04548_);
  and (_05498_, _05496_, _04548_);
  nor (_05499_, _05498_, _05497_);
  nor (_05500_, _05499_, _05480_);
  nor (_05501_, _05500_, _05476_);
  nor (_05502_, _05501_, _02438_);
  or (_05503_, _05502_, _05492_);
  and (_05504_, _05503_, _05487_);
  nor (_05505_, _05482_, _05487_);
  nor (_05506_, _05505_, _05504_);
  nor (_05507_, _05506_, _01963_);
  or (_05508_, _05507_, _04950_);
  nor (_05509_, _05508_, _05486_);
  nor (_05510_, _05509_, _05483_);
  nor (_05511_, _05510_, _04951_);
  and (_05512_, _04134_, _03796_);
  not (_05513_, _04951_);
  nor (_05514_, _05476_, _05513_);
  not (_05515_, _05514_);
  nor (_05516_, _05515_, _05512_);
  or (_05517_, _05516_, _01602_);
  nor (_05518_, _05517_, _05511_);
  nor (_05519_, _02962_, _02786_);
  and (_05520_, _02309_, _02119_);
  and (_05521_, _02676_, _02516_);
  and (_05522_, _05521_, _05520_);
  and (_05523_, _03025_, _02962_);
  not (_05524_, _03101_);
  and (_05525_, _05524_, _03064_);
  and (_05526_, _05525_, _05523_);
  and (_05527_, _05526_, _05522_);
  and (_05528_, _05527_, \oc8051_golden_model_1.P1INREG [7]);
  not (_05529_, _02119_);
  and (_05530_, _02309_, _05529_);
  not (_05531_, _02516_);
  and (_05532_, _02676_, _05531_);
  and (_05533_, _05532_, _05530_);
  and (_05534_, _05533_, _05526_);
  and (_05535_, _05534_, \oc8051_golden_model_1.SBUF [7]);
  nor (_05536_, _05535_, _05528_);
  and (_05537_, _03101_, _03064_);
  and (_05538_, _05537_, _05523_);
  and (_05539_, _05530_, _05521_);
  and (_05540_, _05539_, _05538_);
  and (_05541_, _05540_, \oc8051_golden_model_1.TCON [7]);
  nor (_05542_, _03025_, _02943_);
  and (_05543_, _05542_, _05522_);
  and (_05544_, _05543_, _05525_);
  and (_05545_, _05544_, \oc8051_golden_model_1.PSW [7]);
  nor (_05546_, _05545_, _05541_);
  and (_05547_, _05546_, _05536_);
  not (_05548_, _03064_);
  and (_05549_, _03101_, _05548_);
  and (_05550_, _05549_, _05543_);
  and (_05551_, _05550_, \oc8051_golden_model_1.ACC [7]);
  nor (_05552_, _03101_, _03064_);
  and (_05553_, _05552_, _05543_);
  and (_05554_, _05553_, \oc8051_golden_model_1.B [7]);
  nor (_05555_, _05554_, _05551_);
  and (_05556_, _05538_, _05522_);
  and (_05557_, _05556_, \oc8051_golden_model_1.P0INREG [7]);
  and (_05558_, _05539_, _05526_);
  and (_05559_, _05558_, \oc8051_golden_model_1.SCON [7]);
  nor (_05560_, _05559_, _05557_);
  and (_05561_, _05560_, _05555_);
  and (_05562_, _05561_, _05547_);
  not (_05563_, _02309_);
  nor (_05564_, _02676_, _02516_);
  and (_05565_, _05564_, _05538_);
  and (_05566_, _05565_, _02119_);
  and (_05567_, _05566_, _05563_);
  and (_05568_, _05567_, \oc8051_golden_model_1.PCON [7]);
  and (_05569_, _05566_, _02309_);
  and (_05570_, _05569_, \oc8051_golden_model_1.DPH [7]);
  nor (_05571_, _05570_, _05568_);
  and (_05572_, _05571_, _05562_);
  not (_05573_, _02676_);
  and (_05574_, _05573_, _02516_);
  and (_05575_, _05538_, _05520_);
  and (_05576_, _05575_, _05574_);
  and (_05577_, _05576_, \oc8051_golden_model_1.DPL [7]);
  and (_05578_, _05565_, _05530_);
  and (_05579_, _05578_, \oc8051_golden_model_1.TL1 [7]);
  nor (_05580_, _05579_, _05577_);
  and (_05581_, _05538_, _05530_);
  and (_05582_, _05574_, _05581_);
  and (_05583_, _05582_, \oc8051_golden_model_1.TL0 [7]);
  nor (_05584_, _02309_, _02119_);
  and (_05585_, _05584_, _05538_);
  and (_05587_, _05585_, _05521_);
  and (_05589_, _05587_, \oc8051_golden_model_1.TH0 [7]);
  nor (_05591_, _05589_, _05583_);
  and (_05593_, _05591_, _05580_);
  and (_05595_, _05585_, _05532_);
  and (_05597_, _05595_, \oc8051_golden_model_1.TH1 [7]);
  not (_05599_, _05597_);
  and (_05601_, _05549_, _05523_);
  and (_05603_, _05601_, _05539_);
  and (_05605_, _05603_, \oc8051_golden_model_1.IE [7]);
  and (_05607_, _05552_, _05523_);
  and (_05609_, _05607_, _05522_);
  and (_05611_, _05609_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05613_, _05611_, _05605_);
  and (_05615_, _05601_, _05522_);
  and (_05617_, _05615_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05619_, _05607_, _05539_);
  and (_05621_, _05619_, \oc8051_golden_model_1.IP [7]);
  nor (_05623_, _05621_, _05617_);
  and (_05625_, _05623_, _05613_);
  and (_05627_, _05625_, _05599_);
  and (_05629_, _05581_, _05532_);
  and (_05631_, _05629_, \oc8051_golden_model_1.TMOD [7]);
  and (_05633_, _05575_, _05532_);
  and (_05635_, _05633_, \oc8051_golden_model_1.SP [7]);
  nor (_05637_, _05635_, _05631_);
  and (_05639_, _05637_, _05627_);
  and (_05641_, _05639_, _05593_);
  and (_05643_, _05641_, _05572_);
  not (_05645_, _05643_);
  nor (_05647_, _05645_, _05519_);
  nor (_05648_, _05647_, _05480_);
  nor (_05650_, _05648_, _05476_);
  nor (_05651_, _05650_, _01923_);
  or (_05653_, _05651_, _02019_);
  nor (_05654_, _05653_, _05518_);
  nor (_05656_, _05654_, _05479_);
  or (_05658_, _05656_, _02018_);
  and (_05659_, _04548_, _02943_);
  nor (_05661_, _04548_, _02943_);
  nor (_05662_, _05661_, _05659_);
  and (_05664_, _05662_, _04134_);
  or (_05665_, _05664_, _05476_);
  or (_05667_, _05665_, _05049_);
  and (_05668_, _05667_, _02136_);
  and (_05670_, _05668_, _05658_);
  not (_05671_, \oc8051_golden_model_1.ACC [7]);
  and (_05673_, _04548_, _05671_);
  nor (_05674_, _04548_, _05671_);
  nor (_05676_, _05674_, _05673_);
  and (_05677_, _05676_, _04134_);
  nor (_05679_, _05677_, _05476_);
  nor (_05681_, _05679_, _02136_);
  nor (_05683_, _05681_, _05670_);
  nor (_05685_, _05683_, _02039_);
  not (_05687_, _04548_);
  nor (_05689_, _05476_, _05687_);
  not (_05691_, _05689_);
  nor (_05693_, _05478_, _05076_);
  and (_05695_, _05693_, _05691_);
  nor (_05697_, _05695_, _05685_);
  nor (_05699_, _05697_, _02130_);
  or (_05701_, _05689_, _02131_);
  nor (_05703_, _05701_, _05485_);
  or (_05705_, _05703_, _02016_);
  nor (_05707_, _05705_, _05699_);
  nor (_05709_, _05659_, _05480_);
  nor (_05711_, _05709_, _05476_);
  and (_05713_, _05711_, _02016_);
  nor (_05715_, _05713_, _05707_);
  and (_05717_, _05715_, _05474_);
  nor (_05719_, _05673_, _05480_);
  nor (_05721_, _05719_, _05476_);
  nor (_05723_, _05721_, _05474_);
  or (_05725_, _05723_, _05717_);
  and (_05727_, _05725_, _02168_);
  nor (_05729_, _05501_, _02168_);
  or (_05731_, _05729_, _01594_);
  nor (_05733_, _05731_, _05727_);
  not (_05735_, _04501_);
  not (_05737_, _04204_);
  not (_05739_, _04252_);
  not (_05741_, _04452_);
  and (_05743_, _05741_, _04405_);
  and (_05745_, _05743_, _05739_);
  and (_05747_, _05745_, _05737_);
  nor (_05749_, _04347_, _04299_);
  and (_05751_, _05749_, _05747_);
  and (_05753_, _05751_, _05735_);
  and (_05755_, _05753_, _04548_);
  nor (_05757_, _05753_, _04548_);
  or (_05759_, _05757_, _05755_);
  and (_05761_, _05759_, _04134_);
  nor (_05763_, _05761_, _05476_);
  and (_05765_, _05763_, _01594_);
  nor (_05767_, _05765_, _05733_);
  or (_05769_, _05767_, _26506_);
  or (_05771_, _26505_, \oc8051_golden_model_1.TMOD [7]);
  and (_05773_, _05771_, _25964_);
  and (_25310_, _05773_, _05769_);
  not (_05776_, \oc8051_golden_model_1.TL1 [7]);
  nor (_05778_, _04147_, _05776_);
  and (_05780_, _04147_, _02962_);
  nor (_05782_, _05780_, _05778_);
  and (_05784_, _05782_, _02019_);
  and (_05786_, _04147_, \oc8051_golden_model_1.ACC [7]);
  nor (_05788_, _05786_, _05778_);
  nor (_05790_, _05788_, _01964_);
  nor (_05792_, _05788_, _05488_);
  nor (_05794_, _04571_, _05776_);
  or (_05796_, _05794_, _05792_);
  and (_05798_, _05796_, _02438_);
  not (_05800_, _04147_);
  nor (_05802_, _05499_, _05800_);
  nor (_05804_, _05802_, _05778_);
  nor (_05806_, _05804_, _02438_);
  or (_05808_, _05806_, _05798_);
  and (_05810_, _05808_, _05487_);
  nor (_05812_, _05800_, _02786_);
  nor (_05814_, _05812_, _05778_);
  nor (_05816_, _05814_, _05487_);
  nor (_05818_, _05816_, _05810_);
  nor (_05820_, _05818_, _01963_);
  or (_05822_, _05820_, _04950_);
  nor (_05824_, _05822_, _05790_);
  and (_05826_, _05814_, _04950_);
  nor (_05828_, _05826_, _05824_);
  nor (_05830_, _05828_, _04951_);
  and (_05832_, _04147_, _03796_);
  nor (_05834_, _05778_, _05513_);
  not (_05836_, _05834_);
  nor (_05838_, _05836_, _05832_);
  or (_05840_, _05838_, _01602_);
  nor (_05842_, _05840_, _05830_);
  nor (_05844_, _05647_, _05800_);
  nor (_05846_, _05844_, _05778_);
  nor (_05848_, _05846_, _01923_);
  or (_05850_, _05848_, _02019_);
  nor (_05852_, _05850_, _05842_);
  nor (_05854_, _05852_, _05784_);
  or (_05856_, _05854_, _02018_);
  and (_05858_, _05662_, _04147_);
  or (_05860_, _05858_, _05778_);
  or (_05862_, _05860_, _05049_);
  and (_05864_, _05862_, _02136_);
  and (_05866_, _05864_, _05856_);
  and (_05868_, _05676_, _04147_);
  nor (_05870_, _05868_, _05778_);
  nor (_05872_, _05870_, _02136_);
  nor (_05874_, _05872_, _05866_);
  nor (_05876_, _05874_, _02039_);
  nor (_05878_, _05778_, _05687_);
  not (_05880_, _05878_);
  nor (_05882_, _05782_, _05076_);
  and (_05884_, _05882_, _05880_);
  nor (_05886_, _05884_, _05876_);
  nor (_05888_, _05886_, _02130_);
  or (_05890_, _05878_, _02131_);
  nor (_05892_, _05890_, _05788_);
  or (_05894_, _05892_, _02016_);
  nor (_05896_, _05894_, _05888_);
  nor (_05898_, _05659_, _05800_);
  nor (_05900_, _05898_, _05778_);
  and (_05902_, _05900_, _02016_);
  nor (_05904_, _05902_, _05896_);
  and (_05906_, _05904_, _05474_);
  nor (_05908_, _05673_, _05800_);
  nor (_05910_, _05908_, _05778_);
  nor (_05912_, _05910_, _05474_);
  or (_05914_, _05912_, _05906_);
  and (_05916_, _05914_, _02168_);
  nor (_05918_, _05804_, _02168_);
  or (_05920_, _05918_, _01594_);
  nor (_05922_, _05920_, _05916_);
  and (_05924_, _05759_, _04147_);
  nor (_05926_, _05924_, _05778_);
  and (_05928_, _05926_, _01594_);
  nor (_05930_, _05928_, _05922_);
  or (_05932_, _05930_, _26506_);
  or (_05934_, _26505_, \oc8051_golden_model_1.TL1 [7]);
  and (_05936_, _05934_, _25964_);
  and (_25312_, _05936_, _05932_);
  not (_05939_, \oc8051_golden_model_1.TL0 [7]);
  nor (_05941_, _04143_, _05939_);
  and (_05943_, _04143_, _02962_);
  nor (_05945_, _05943_, _05941_);
  and (_05947_, _05945_, _02019_);
  and (_05949_, _04143_, \oc8051_golden_model_1.ACC [7]);
  nor (_05951_, _05949_, _05941_);
  nor (_05953_, _05951_, _01964_);
  nor (_05955_, _05951_, _05488_);
  nor (_05957_, _04571_, _05939_);
  or (_05959_, _05957_, _05955_);
  and (_05961_, _05959_, _02438_);
  not (_05963_, _04143_);
  nor (_05965_, _05499_, _05963_);
  nor (_05967_, _05965_, _05941_);
  nor (_05969_, _05967_, _02438_);
  or (_05971_, _05969_, _05961_);
  and (_05973_, _05971_, _05487_);
  nor (_05975_, _05963_, _02786_);
  nor (_05977_, _05975_, _05941_);
  nor (_05979_, _05977_, _05487_);
  nor (_05981_, _05979_, _05973_);
  nor (_05982_, _05981_, _01963_);
  or (_05983_, _05982_, _04950_);
  nor (_05984_, _05983_, _05953_);
  and (_05985_, _05977_, _04950_);
  nor (_05986_, _05985_, _05984_);
  nor (_05987_, _05986_, _04951_);
  and (_05988_, _04143_, _03796_);
  nor (_05989_, _05941_, _05513_);
  not (_05990_, _05989_);
  nor (_05991_, _05990_, _05988_);
  or (_05992_, _05991_, _01602_);
  nor (_05993_, _05992_, _05987_);
  nor (_05994_, _05647_, _05963_);
  nor (_05995_, _05994_, _05941_);
  nor (_05996_, _05995_, _01923_);
  or (_05997_, _05996_, _02019_);
  nor (_05998_, _05997_, _05993_);
  nor (_05999_, _05998_, _05947_);
  or (_06000_, _05999_, _02018_);
  and (_06001_, _05662_, _04143_);
  or (_06002_, _06001_, _05941_);
  or (_06003_, _06002_, _05049_);
  and (_06004_, _06003_, _02136_);
  and (_06005_, _06004_, _06000_);
  and (_06006_, _05676_, _04143_);
  nor (_06007_, _06006_, _05941_);
  nor (_06008_, _06007_, _02136_);
  nor (_06009_, _06008_, _06005_);
  nor (_06010_, _06009_, _02039_);
  nor (_06011_, _05941_, _05687_);
  not (_06012_, _06011_);
  nor (_06013_, _05945_, _05076_);
  and (_06014_, _06013_, _06012_);
  nor (_06015_, _06014_, _06010_);
  nor (_06016_, _06015_, _02130_);
  or (_06017_, _06011_, _02131_);
  nor (_06018_, _06017_, _05951_);
  or (_06019_, _06018_, _02016_);
  nor (_06020_, _06019_, _06016_);
  nor (_06021_, _05659_, _05963_);
  nor (_06022_, _06021_, _05941_);
  and (_06023_, _06022_, _02016_);
  nor (_06024_, _06023_, _06020_);
  and (_06025_, _06024_, _05474_);
  nor (_06026_, _05673_, _05963_);
  nor (_06027_, _06026_, _05941_);
  nor (_06028_, _06027_, _05474_);
  or (_06029_, _06028_, _06025_);
  and (_06030_, _06029_, _02168_);
  nor (_06031_, _05967_, _02168_);
  or (_06032_, _06031_, _01594_);
  nor (_06033_, _06032_, _06030_);
  and (_06034_, _05759_, _04143_);
  nor (_06035_, _06034_, _05941_);
  and (_06036_, _06035_, _01594_);
  nor (_06037_, _06036_, _06033_);
  or (_06038_, _06037_, _26506_);
  or (_06039_, _26505_, \oc8051_golden_model_1.TL0 [7]);
  and (_06040_, _06039_, _25964_);
  and (_25313_, _06040_, _06038_);
  not (_06041_, \oc8051_golden_model_1.TH1 [7]);
  nor (_06042_, _04138_, _06041_);
  and (_06043_, _04138_, _02962_);
  nor (_06044_, _06043_, _06042_);
  and (_06045_, _06044_, _02019_);
  not (_06046_, _04138_);
  nor (_06047_, _06046_, _02786_);
  nor (_06048_, _06047_, _06042_);
  and (_06049_, _06048_, _04950_);
  and (_06050_, _04138_, \oc8051_golden_model_1.ACC [7]);
  nor (_06051_, _06050_, _06042_);
  nor (_06052_, _06051_, _05488_);
  nor (_06053_, _04571_, _06041_);
  or (_06054_, _06053_, _06052_);
  and (_06055_, _06054_, _02438_);
  nor (_06056_, _05499_, _06046_);
  nor (_06057_, _06056_, _06042_);
  nor (_06058_, _06057_, _02438_);
  or (_06059_, _06058_, _06055_);
  and (_06060_, _06059_, _05487_);
  nor (_06061_, _06048_, _05487_);
  nor (_06062_, _06061_, _06060_);
  nor (_06063_, _06062_, _01963_);
  nor (_06064_, _06051_, _01964_);
  nor (_06065_, _06064_, _04950_);
  not (_06066_, _06065_);
  nor (_06067_, _06066_, _06063_);
  nor (_06068_, _06067_, _06049_);
  nor (_06069_, _06068_, _04951_);
  and (_06070_, _04138_, _03796_);
  nor (_06071_, _06042_, _05513_);
  not (_06072_, _06071_);
  nor (_06073_, _06072_, _06070_);
  or (_06074_, _06073_, _01602_);
  nor (_06075_, _06074_, _06069_);
  nor (_06076_, _05647_, _06046_);
  nor (_06077_, _06076_, _06042_);
  nor (_06078_, _06077_, _01923_);
  or (_06079_, _06078_, _02019_);
  nor (_06080_, _06079_, _06075_);
  nor (_06081_, _06080_, _06045_);
  or (_06082_, _06081_, _02018_);
  and (_06083_, _05662_, _04138_);
  or (_06084_, _06083_, _06042_);
  or (_06085_, _06084_, _05049_);
  and (_06086_, _06085_, _02136_);
  and (_06087_, _06086_, _06082_);
  and (_06088_, _05676_, _04138_);
  nor (_06089_, _06088_, _06042_);
  nor (_06090_, _06089_, _02136_);
  nor (_06091_, _06090_, _06087_);
  nor (_06092_, _06091_, _02039_);
  nor (_06093_, _06042_, _05687_);
  not (_06094_, _06093_);
  nor (_06095_, _06044_, _05076_);
  and (_06096_, _06095_, _06094_);
  nor (_06097_, _06096_, _06092_);
  nor (_06098_, _06097_, _02130_);
  or (_06099_, _06093_, _02131_);
  nor (_06100_, _06099_, _06051_);
  or (_06101_, _06100_, _02016_);
  nor (_06102_, _06101_, _06098_);
  nor (_06103_, _05659_, _06046_);
  nor (_06104_, _06103_, _06042_);
  and (_06105_, _06104_, _02016_);
  nor (_06106_, _06105_, _06102_);
  and (_06107_, _06106_, _05474_);
  nor (_06108_, _05673_, _06046_);
  nor (_06109_, _06108_, _06042_);
  nor (_06110_, _06109_, _05474_);
  or (_06111_, _06110_, _06107_);
  and (_06112_, _06111_, _02168_);
  nor (_06113_, _06057_, _02168_);
  or (_06114_, _06113_, _01594_);
  nor (_06115_, _06114_, _06112_);
  and (_06116_, _05759_, _04138_);
  nor (_06117_, _06116_, _06042_);
  and (_06118_, _06117_, _01594_);
  nor (_06119_, _06118_, _06115_);
  or (_06120_, _06119_, _26506_);
  or (_06121_, _26505_, \oc8051_golden_model_1.TH1 [7]);
  and (_06122_, _06121_, _25964_);
  and (_25314_, _06122_, _06120_);
  not (_06123_, \oc8051_golden_model_1.TH0 [7]);
  nor (_06124_, _04125_, _06123_);
  and (_06125_, _04125_, _02962_);
  nor (_06126_, _06125_, _06124_);
  and (_06127_, _06126_, _02019_);
  not (_06128_, _04125_);
  nor (_06129_, _06128_, _02786_);
  nor (_06130_, _06129_, _06124_);
  and (_06131_, _06130_, _04950_);
  and (_06132_, _04125_, \oc8051_golden_model_1.ACC [7]);
  nor (_06133_, _06132_, _06124_);
  nor (_06134_, _06133_, _01964_);
  nor (_06135_, _06133_, _05488_);
  nor (_06136_, _04571_, _06123_);
  or (_06137_, _06136_, _06135_);
  and (_06138_, _06137_, _02438_);
  nor (_06139_, _05499_, _06128_);
  nor (_06140_, _06139_, _06124_);
  nor (_06141_, _06140_, _02438_);
  or (_06142_, _06141_, _06138_);
  and (_06143_, _06142_, _05487_);
  nor (_06144_, _06130_, _05487_);
  nor (_06145_, _06144_, _06143_);
  nor (_06146_, _06145_, _01963_);
  or (_06147_, _06146_, _04950_);
  nor (_06148_, _06147_, _06134_);
  nor (_06149_, _06148_, _06131_);
  nor (_06150_, _06149_, _04951_);
  and (_06151_, _04125_, _03796_);
  nor (_06152_, _06124_, _05513_);
  not (_06153_, _06152_);
  nor (_06154_, _06153_, _06151_);
  or (_06155_, _06154_, _01602_);
  nor (_06156_, _06155_, _06150_);
  nor (_06157_, _05647_, _06128_);
  nor (_06158_, _06157_, _06124_);
  nor (_06159_, _06158_, _01923_);
  or (_06160_, _06159_, _02019_);
  nor (_06161_, _06160_, _06156_);
  nor (_06162_, _06161_, _06127_);
  or (_06163_, _06162_, _02018_);
  and (_06164_, _05662_, _04125_);
  or (_06165_, _06164_, _06124_);
  or (_06166_, _06165_, _05049_);
  and (_06167_, _06166_, _02136_);
  and (_06168_, _06167_, _06163_);
  and (_06169_, _05676_, _04125_);
  nor (_06170_, _06169_, _06124_);
  nor (_06171_, _06170_, _02136_);
  nor (_06172_, _06171_, _06168_);
  nor (_06173_, _06172_, _02039_);
  nor (_06174_, _06124_, _05687_);
  not (_06175_, _06174_);
  nor (_06176_, _06126_, _05076_);
  and (_06177_, _06176_, _06175_);
  nor (_06178_, _06177_, _06173_);
  nor (_06179_, _06178_, _02130_);
  or (_06180_, _06174_, _02131_);
  nor (_06181_, _06180_, _06133_);
  or (_06182_, _06181_, _02016_);
  nor (_06183_, _06182_, _06179_);
  nor (_06184_, _05659_, _06128_);
  nor (_06185_, _06184_, _06124_);
  and (_06186_, _06185_, _02016_);
  nor (_06187_, _06186_, _06183_);
  and (_06188_, _06187_, _05474_);
  nor (_06189_, _05673_, _06128_);
  nor (_06190_, _06189_, _06124_);
  nor (_06191_, _06190_, _05474_);
  or (_06192_, _06191_, _06188_);
  and (_06193_, _06192_, _02168_);
  nor (_06194_, _06140_, _02168_);
  or (_06195_, _06194_, _01594_);
  nor (_06196_, _06195_, _06193_);
  and (_06197_, _05759_, _04125_);
  nor (_06198_, _06197_, _06124_);
  and (_06199_, _06198_, _01594_);
  nor (_06200_, _06199_, _06196_);
  or (_06201_, _06200_, _26506_);
  or (_06202_, _26505_, \oc8051_golden_model_1.TH0 [7]);
  and (_06203_, _06202_, _25964_);
  and (_25315_, _06203_, _06201_);
  not (_06204_, \oc8051_golden_model_1.TCON [7]);
  nor (_06205_, _04119_, _06204_);
  not (_06206_, _04119_);
  nor (_06207_, _06206_, _02786_);
  nor (_06208_, _06207_, _06205_);
  and (_06209_, _06208_, _04950_);
  nor (_06210_, _05167_, _06204_);
  not (_06211_, _06210_);
  and (_06212_, _04099_, \oc8051_golden_model_1.P0 [7]);
  and (_06213_, _05189_, \oc8051_golden_model_1.P2 [7]);
  nor (_06214_, _06213_, _06212_);
  and (_06215_, _05195_, \oc8051_golden_model_1.P1 [7]);
  and (_06216_, _05191_, \oc8051_golden_model_1.P3 [7]);
  nor (_06217_, _06216_, _06215_);
  and (_06218_, _06217_, _06214_);
  and (_06219_, _06218_, _05268_);
  and (_06220_, _06219_, _05265_);
  and (_06221_, _06220_, _04079_);
  nor (_06222_, _06221_, _05255_);
  and (_06223_, _06222_, _06211_);
  nand (_06224_, _06221_, _05255_);
  and (_06225_, _06224_, _05167_);
  nor (_06226_, _06225_, _06210_);
  or (_06227_, _06226_, _04885_);
  nor (_06228_, _06227_, _06223_);
  not (_06229_, _01957_);
  nor (_06230_, _05499_, _06206_);
  nor (_06231_, _06230_, _06205_);
  and (_06232_, _06231_, _01969_);
  not (_06233_, _01968_);
  and (_06234_, _04119_, \oc8051_golden_model_1.ACC [7]);
  nor (_06235_, _06234_, _06205_);
  nor (_06236_, _06235_, _05488_);
  nor (_06237_, _04571_, _06204_);
  or (_06238_, _06237_, _01969_);
  nor (_06239_, _06238_, _06236_);
  or (_06240_, _06239_, _06233_);
  nor (_06241_, _06240_, _06232_);
  nor (_06242_, _06208_, _05487_);
  nor (_06243_, _06226_, _02223_);
  nor (_06244_, _06243_, _06242_);
  nand (_06245_, _06244_, _01964_);
  or (_06246_, _06245_, _06241_);
  nand (_06247_, _06235_, _01963_);
  and (_06248_, _06247_, _06246_);
  and (_06249_, _06248_, _06229_);
  nor (_06250_, _06221_, _04176_);
  and (_06251_, _06250_, _05167_);
  nor (_06252_, _06251_, _06210_);
  nor (_06253_, _06252_, _06229_);
  or (_06254_, _06253_, _06249_);
  and (_06255_, _06254_, _04885_);
  nor (_06256_, _06255_, _06228_);
  nor (_06257_, _06256_, _01924_);
  not (_06258_, _05167_);
  nor (_06259_, _05278_, _04176_);
  and (_06260_, _04100_, \oc8051_golden_model_1.PSW [7]);
  and (_06261_, _06260_, _02264_);
  nor (_06262_, _06261_, _06259_);
  nor (_06263_, _06262_, _06258_);
  nor (_06264_, _06263_, _06210_);
  nor (_06265_, _06264_, _01925_);
  nor (_06266_, _06265_, _04950_);
  not (_06267_, _06266_);
  nor (_06268_, _06267_, _06257_);
  nor (_06269_, _06268_, _06209_);
  nor (_06270_, _06269_, _04951_);
  and (_06271_, _04119_, _03796_);
  nor (_06272_, _06205_, _05513_);
  not (_06273_, _06272_);
  nor (_06274_, _06273_, _06271_);
  nor (_06275_, _06274_, _01602_);
  not (_06276_, _06275_);
  nor (_06277_, _06276_, _06270_);
  not (_06278_, _02020_);
  nor (_06279_, _05647_, _06206_);
  nor (_06280_, _06279_, _06205_);
  nor (_06281_, _06280_, _01923_);
  or (_06282_, _06281_, _06278_);
  or (_06283_, _06282_, _06277_);
  and (_06284_, _05662_, _04119_);
  or (_06285_, _06205_, _05049_);
  or (_06286_, _06285_, _06284_);
  and (_06287_, _04119_, _02962_);
  nor (_06288_, _06287_, _06205_);
  and (_06289_, _06288_, _02019_);
  nor (_06290_, _06289_, _02135_);
  and (_06291_, _06290_, _06286_);
  and (_06292_, _06291_, _06283_);
  and (_06293_, _05676_, _04119_);
  nor (_06294_, _06293_, _06205_);
  nor (_06295_, _06294_, _02136_);
  nor (_06296_, _06295_, _06292_);
  nor (_06297_, _06296_, _02039_);
  nor (_06298_, _06205_, _05687_);
  not (_06299_, _06298_);
  nor (_06300_, _06288_, _05076_);
  and (_06301_, _06300_, _06299_);
  nor (_06302_, _06301_, _06297_);
  nor (_06303_, _06302_, _02130_);
  or (_06304_, _06298_, _02131_);
  nor (_06305_, _06304_, _06235_);
  or (_06306_, _06305_, _02016_);
  nor (_06307_, _06306_, _06303_);
  nor (_06308_, _05659_, _06206_);
  nor (_06309_, _06308_, _06205_);
  and (_06310_, _06309_, _02016_);
  nor (_06311_, _06310_, _06307_);
  and (_06312_, _06311_, _05474_);
  nor (_06313_, _05673_, _06206_);
  nor (_06314_, _06313_, _06205_);
  nor (_06315_, _06314_, _05474_);
  or (_06316_, _06315_, _06312_);
  and (_06317_, _06316_, _02168_);
  nor (_06318_, _06231_, _02168_);
  or (_06319_, _06318_, _02025_);
  or (_06320_, _06319_, _06317_);
  nand (_06321_, _06252_, _02025_);
  and (_06322_, _06321_, _06320_);
  nor (_06323_, _06322_, _01594_);
  and (_06324_, _05759_, _04119_);
  nor (_06325_, _06324_, _06205_);
  and (_06326_, _06325_, _01594_);
  nor (_06327_, _06326_, _06323_);
  or (_06328_, _06327_, _26506_);
  or (_06329_, _26505_, \oc8051_golden_model_1.TCON [7]);
  and (_06330_, _06329_, _25964_);
  and (_25317_, _06330_, _06328_);
  not (_06331_, \oc8051_golden_model_1.SP [7]);
  nor (_06332_, _04111_, _06331_);
  and (_06333_, _05676_, _04111_);
  or (_06334_, _06333_, _06332_);
  and (_06335_, _06334_, _02135_);
  not (_06336_, _04111_);
  nor (_06337_, _06336_, _02786_);
  or (_06338_, _06332_, _04951_);
  or (_06339_, _06338_, _06337_);
  and (_06340_, _06339_, _04953_);
  nor (_06341_, _05499_, _06336_);
  or (_06342_, _06341_, _06332_);
  or (_06343_, _06342_, _02438_);
  and (_06344_, _04396_, \oc8051_golden_model_1.ACC [7]);
  or (_06345_, _06344_, _06332_);
  or (_06346_, _06345_, _05488_);
  or (_06347_, _04571_, \oc8051_golden_model_1.SP [7]);
  and (_06348_, _06347_, _01625_);
  and (_06349_, _06348_, _06346_);
  and (_06350_, \oc8051_golden_model_1.SP [3], \oc8051_golden_model_1.SP [2]);
  and (_06351_, _06350_, \oc8051_golden_model_1.SP [1]);
  and (_06352_, _06351_, \oc8051_golden_model_1.SP [4]);
  and (_06353_, _06352_, \oc8051_golden_model_1.SP [5]);
  and (_06354_, _06353_, \oc8051_golden_model_1.SP [6]);
  or (_06355_, _06354_, \oc8051_golden_model_1.SP [7]);
  nand (_06356_, _06354_, \oc8051_golden_model_1.SP [7]);
  and (_06357_, _06356_, _06355_);
  and (_06358_, _06357_, _04568_);
  or (_06359_, _06358_, _01969_);
  or (_06360_, _06359_, _06349_);
  and (_06361_, _06360_, _01621_);
  and (_06362_, _06361_, _06343_);
  not (_06363_, _01621_);
  and (_06364_, _06357_, _06363_);
  or (_06365_, _06364_, _01967_);
  or (_06366_, _06365_, _06362_);
  not (_06367_, \oc8051_golden_model_1.SP [6]);
  not (_06368_, \oc8051_golden_model_1.SP [5]);
  not (_06369_, \oc8051_golden_model_1.SP [4]);
  and (_06370_, _03418_, _06369_);
  and (_06371_, _06370_, _06368_);
  and (_06372_, _06371_, _06367_);
  and (_06373_, _06372_, _02441_);
  nor (_06374_, _06373_, _06331_);
  and (_06375_, _06373_, _06331_);
  nor (_06376_, _06375_, _06374_);
  nand (_06377_, _06376_, _01967_);
  and (_06378_, _06377_, _06366_);
  or (_06379_, _06378_, _01963_);
  or (_06380_, _06345_, _01964_);
  and (_06382_, _06380_, _02457_);
  and (_06383_, _06382_, _06379_);
  and (_06384_, _06350_, _03399_);
  and (_06385_, _06384_, \oc8051_golden_model_1.SP [4]);
  and (_06386_, _06385_, \oc8051_golden_model_1.SP [5]);
  and (_06387_, _06386_, \oc8051_golden_model_1.SP [6]);
  nor (_06388_, _06387_, _06331_);
  and (_06389_, _06387_, _06331_);
  or (_06390_, _06389_, _06388_);
  nand (_06391_, _06390_, _01953_);
  not (_06393_, _01632_);
  nor (_06394_, _01606_, _06393_);
  nand (_06395_, _06394_, _06391_);
  or (_06396_, _06395_, _06383_);
  not (_06397_, _04950_);
  or (_06398_, _06394_, _06357_);
  and (_06399_, _06398_, _06397_);
  and (_06400_, _06399_, _06396_);
  or (_06401_, _06400_, _06340_);
  or (_06402_, _06332_, _05513_);
  and (_06404_, _04396_, _03796_);
  or (_06405_, _06404_, _06402_);
  and (_06406_, _06405_, _01923_);
  and (_06407_, _06406_, _06401_);
  nor (_06408_, _05647_, _06336_);
  or (_06409_, _06408_, _06332_);
  and (_06410_, _06409_, _01602_);
  or (_06411_, _06410_, _02019_);
  or (_06412_, _06411_, _06407_);
  and (_06413_, _04396_, _02962_);
  or (_06415_, _06413_, _06332_);
  or (_06416_, _06415_, _04979_);
  and (_06417_, _06416_, _06412_);
  or (_06418_, _06417_, _01650_);
  or (_06419_, _06357_, _01651_);
  and (_06420_, _06419_, _06418_);
  or (_06421_, _06420_, _02018_);
  and (_06422_, _05662_, _04111_);
  or (_06423_, _06332_, _05049_);
  or (_06424_, _06423_, _06422_);
  and (_06426_, _06424_, _02136_);
  and (_06427_, _06426_, _06421_);
  or (_06428_, _06427_, _06335_);
  and (_06429_, _06428_, _05076_);
  or (_06430_, _06332_, _05687_);
  and (_06431_, _06415_, _02039_);
  and (_06432_, _06431_, _06430_);
  or (_06433_, _06432_, _06429_);
  and (_06434_, _06433_, _05082_);
  and (_06435_, _06357_, _01666_);
  or (_06437_, _06435_, _02016_);
  and (_06438_, _06345_, _02130_);
  and (_06439_, _06438_, _06430_);
  or (_06440_, _06439_, _06437_);
  or (_06441_, _06440_, _06434_);
  not (_06442_, _04396_);
  nor (_06443_, _05659_, _06442_);
  or (_06444_, _06443_, _06332_);
  or (_06445_, _06444_, _05104_);
  and (_06446_, _06445_, _06441_);
  or (_06447_, _06446_, _02126_);
  nor (_06448_, _05673_, _06336_);
  or (_06449_, _06332_, _05474_);
  or (_06450_, _06449_, _06448_);
  and (_06451_, _06450_, _02718_);
  and (_06452_, _06451_, _06447_);
  or (_06453_, _06372_, \oc8051_golden_model_1.SP [7]);
  nand (_06454_, _06372_, \oc8051_golden_model_1.SP [7]);
  and (_06455_, _06454_, _06453_);
  and (_06456_, _06455_, _02146_);
  or (_06457_, _06456_, _01660_);
  or (_06458_, _06457_, _06452_);
  or (_06459_, _06357_, _05157_);
  and (_06460_, _06459_, _06458_);
  or (_06461_, _06460_, _01585_);
  or (_06462_, _06455_, _01596_);
  and (_06463_, _06462_, _02168_);
  and (_06464_, _06463_, _06461_);
  and (_06465_, _06342_, _02164_);
  nor (_06466_, _02023_, _01670_);
  not (_06467_, _06466_);
  or (_06468_, _06467_, _06465_);
  or (_06469_, _06468_, _06464_);
  or (_06470_, _06466_, _06357_);
  and (_06471_, _06470_, _01595_);
  and (_06472_, _06471_, _06469_);
  and (_06473_, _05759_, _04111_);
  or (_06474_, _06473_, _06332_);
  and (_06475_, _06474_, _01594_);
  or (_06476_, _06475_, _26506_);
  or (_06477_, _06476_, _06472_);
  or (_06478_, _26505_, \oc8051_golden_model_1.SP [7]);
  and (_06479_, _06478_, _25964_);
  and (_25318_, _06479_, _06477_);
  not (_06480_, \oc8051_golden_model_1.SCON [7]);
  nor (_06481_, _04129_, _06480_);
  not (_06482_, _04129_);
  nor (_06483_, _06482_, _02786_);
  nor (_06484_, _06483_, _06481_);
  and (_06485_, _06484_, _04950_);
  nor (_06486_, _05184_, _06480_);
  not (_06487_, _06486_);
  and (_06488_, _06487_, _06222_);
  and (_06489_, _06224_, _05184_);
  nor (_06490_, _06489_, _06486_);
  or (_06491_, _06490_, _04885_);
  nor (_06492_, _06491_, _06488_);
  nor (_06493_, _05499_, _06482_);
  nor (_06494_, _06493_, _06481_);
  and (_06495_, _06494_, _01969_);
  and (_06496_, _04129_, \oc8051_golden_model_1.ACC [7]);
  nor (_06497_, _06496_, _06481_);
  nor (_06498_, _06497_, _05488_);
  nor (_06499_, _04571_, _06480_);
  or (_06500_, _06499_, _01969_);
  nor (_06501_, _06500_, _06498_);
  or (_06502_, _06501_, _06233_);
  nor (_06503_, _06502_, _06495_);
  nor (_06504_, _06484_, _05487_);
  nor (_06505_, _06490_, _02223_);
  nor (_06506_, _06505_, _06504_);
  nand (_06507_, _06506_, _01964_);
  or (_06508_, _06507_, _06503_);
  nand (_06509_, _06497_, _01963_);
  and (_06510_, _06509_, _06508_);
  and (_06511_, _06510_, _06229_);
  and (_06512_, _06250_, _05184_);
  nor (_06513_, _06512_, _06486_);
  nor (_06514_, _06513_, _06229_);
  or (_06515_, _06514_, _06511_);
  and (_06516_, _06515_, _04885_);
  nor (_06517_, _06516_, _06492_);
  nor (_06518_, _06517_, _01924_);
  not (_06519_, _05184_);
  nor (_06520_, _06262_, _06519_);
  nor (_06521_, _06520_, _06486_);
  nor (_06522_, _06521_, _01925_);
  nor (_06523_, _06522_, _04950_);
  not (_06524_, _06523_);
  nor (_06525_, _06524_, _06518_);
  nor (_06526_, _06525_, _06485_);
  nor (_06527_, _06526_, _04951_);
  and (_06528_, _04129_, _03796_);
  nor (_06529_, _06481_, _05513_);
  not (_06530_, _06529_);
  nor (_06531_, _06530_, _06528_);
  nor (_06532_, _06531_, _01602_);
  not (_06533_, _06532_);
  nor (_06534_, _06533_, _06527_);
  nor (_06535_, _05647_, _06482_);
  nor (_06536_, _06535_, _06481_);
  nor (_06537_, _06536_, _01923_);
  or (_06538_, _06537_, _06278_);
  or (_06539_, _06538_, _06534_);
  and (_06540_, _05662_, _04129_);
  or (_06541_, _06481_, _05049_);
  or (_06542_, _06541_, _06540_);
  and (_06543_, _04129_, _02962_);
  nor (_06544_, _06543_, _06481_);
  and (_06545_, _06544_, _02019_);
  nor (_06546_, _06545_, _02135_);
  and (_06547_, _06546_, _06542_);
  and (_06548_, _06547_, _06539_);
  and (_06549_, _05676_, _04129_);
  nor (_06550_, _06549_, _06481_);
  nor (_06551_, _06550_, _02136_);
  nor (_06552_, _06551_, _06548_);
  nor (_06553_, _06552_, _02039_);
  nor (_06554_, _06481_, _05687_);
  not (_06555_, _06554_);
  nor (_06556_, _06544_, _05076_);
  and (_06557_, _06556_, _06555_);
  nor (_06558_, _06557_, _06553_);
  nor (_06559_, _06558_, _02130_);
  or (_06560_, _06554_, _02131_);
  nor (_06561_, _06560_, _06497_);
  or (_06562_, _06561_, _02016_);
  nor (_06563_, _06562_, _06559_);
  nor (_06564_, _05659_, _06482_);
  nor (_06565_, _06564_, _06481_);
  and (_06566_, _06565_, _02016_);
  nor (_06567_, _06566_, _06563_);
  and (_06568_, _06567_, _05474_);
  nor (_06569_, _05673_, _06482_);
  nor (_06570_, _06569_, _06481_);
  nor (_06571_, _06570_, _05474_);
  or (_06572_, _06571_, _06568_);
  and (_06573_, _06572_, _02168_);
  nor (_06574_, _06494_, _02168_);
  or (_06575_, _06574_, _02025_);
  or (_06576_, _06575_, _06573_);
  nand (_06577_, _06513_, _02025_);
  and (_06578_, _06577_, _06576_);
  nor (_06579_, _06578_, _01594_);
  and (_06580_, _05759_, _04129_);
  nor (_06581_, _06580_, _06481_);
  and (_06582_, _06581_, _01594_);
  nor (_06583_, _06582_, _06579_);
  or (_06584_, _06583_, _26506_);
  or (_06585_, _26505_, \oc8051_golden_model_1.SCON [7]);
  and (_06586_, _06585_, _25964_);
  and (_25320_, _06586_, _06584_);
  not (_06587_, \oc8051_golden_model_1.SBUF [7]);
  nor (_06588_, _04180_, _06587_);
  and (_06589_, _04180_, _02962_);
  nor (_06590_, _06589_, _06588_);
  and (_06591_, _06590_, _02019_);
  and (_06592_, _04180_, \oc8051_golden_model_1.ACC [7]);
  nor (_06593_, _06592_, _06588_);
  nor (_06594_, _06593_, _01964_);
  nor (_06595_, _06593_, _05488_);
  nor (_06596_, _04571_, _06587_);
  or (_06597_, _06596_, _06595_);
  and (_06598_, _06597_, _02438_);
  not (_06599_, _04180_);
  nor (_06600_, _05499_, _06599_);
  nor (_06601_, _06600_, _06588_);
  nor (_06602_, _06601_, _02438_);
  or (_06603_, _06602_, _06598_);
  and (_06604_, _06603_, _05487_);
  nor (_06605_, _06599_, _02786_);
  nor (_06606_, _06605_, _06588_);
  nor (_06607_, _06606_, _05487_);
  nor (_06608_, _06607_, _06604_);
  nor (_06609_, _06608_, _01963_);
  or (_06610_, _06609_, _04950_);
  nor (_06611_, _06610_, _06594_);
  and (_06612_, _06606_, _04950_);
  nor (_06613_, _06612_, _06611_);
  nor (_06614_, _06613_, _04951_);
  and (_06615_, _04180_, _03796_);
  nor (_06616_, _06588_, _05513_);
  not (_06617_, _06616_);
  nor (_06618_, _06617_, _06615_);
  or (_06619_, _06618_, _01602_);
  nor (_06620_, _06619_, _06614_);
  nor (_06621_, _05647_, _06599_);
  nor (_06622_, _06621_, _06588_);
  nor (_06623_, _06622_, _01923_);
  or (_06624_, _06623_, _02019_);
  nor (_06625_, _06624_, _06620_);
  nor (_06626_, _06625_, _06591_);
  or (_06627_, _06626_, _02018_);
  and (_06628_, _05662_, _04180_);
  or (_06629_, _06628_, _06588_);
  or (_06630_, _06629_, _05049_);
  and (_06631_, _06630_, _02136_);
  and (_06632_, _06631_, _06627_);
  and (_06633_, _05676_, _04180_);
  nor (_06634_, _06633_, _06588_);
  nor (_06635_, _06634_, _02136_);
  nor (_06636_, _06635_, _06632_);
  nor (_06637_, _06636_, _02039_);
  nor (_06638_, _06588_, _05687_);
  not (_06639_, _06638_);
  nor (_06640_, _06590_, _05076_);
  and (_06641_, _06640_, _06639_);
  nor (_06642_, _06641_, _06637_);
  nor (_06643_, _06642_, _02130_);
  or (_06644_, _06638_, _02131_);
  nor (_06645_, _06644_, _06593_);
  or (_06646_, _06645_, _02016_);
  nor (_06647_, _06646_, _06643_);
  nor (_06648_, _05659_, _06599_);
  nor (_06649_, _06648_, _06588_);
  and (_06650_, _06649_, _02016_);
  nor (_06651_, _06650_, _06647_);
  and (_06652_, _06651_, _05474_);
  nor (_06653_, _05673_, _06599_);
  nor (_06654_, _06653_, _06588_);
  nor (_06655_, _06654_, _05474_);
  or (_06656_, _06655_, _06652_);
  and (_06657_, _06656_, _02168_);
  nor (_06658_, _06601_, _02168_);
  or (_06659_, _06658_, _01594_);
  nor (_06660_, _06659_, _06657_);
  and (_06661_, _05759_, _04180_);
  nor (_06662_, _06661_, _06588_);
  and (_06663_, _06662_, _01594_);
  nor (_06664_, _06663_, _06660_);
  or (_06665_, _06664_, _26506_);
  or (_06666_, _26505_, \oc8051_golden_model_1.SBUF [7]);
  and (_06667_, _06666_, _25964_);
  and (_25322_, _06667_, _06665_);
  not (_06668_, \oc8051_golden_model_1.PCON [7]);
  nor (_06669_, _04177_, _06668_);
  and (_06670_, _04177_, _02962_);
  nor (_06671_, _06670_, _06669_);
  and (_06672_, _06671_, _02019_);
  and (_06673_, _04177_, \oc8051_golden_model_1.ACC [7]);
  nor (_06674_, _06673_, _06669_);
  nor (_06675_, _06674_, _01964_);
  nor (_06676_, _06674_, _05488_);
  nor (_06677_, _04571_, _06668_);
  or (_06678_, _06677_, _06676_);
  and (_06679_, _06678_, _02438_);
  not (_06680_, _04177_);
  nor (_06681_, _05499_, _06680_);
  nor (_06682_, _06681_, _06669_);
  nor (_06683_, _06682_, _02438_);
  or (_06684_, _06683_, _06679_);
  and (_06685_, _06684_, _05487_);
  nor (_06686_, _06680_, _02786_);
  nor (_06687_, _06686_, _06669_);
  nor (_06688_, _06687_, _05487_);
  nor (_06689_, _06688_, _06685_);
  nor (_06690_, _06689_, _01963_);
  or (_06691_, _06690_, _04950_);
  nor (_06692_, _06691_, _06675_);
  and (_06693_, _06687_, _04950_);
  nor (_06694_, _06693_, _06692_);
  nor (_06695_, _06694_, _04951_);
  and (_06696_, _04177_, _03796_);
  nor (_06697_, _06669_, _05513_);
  not (_06698_, _06697_);
  nor (_06699_, _06698_, _06696_);
  or (_06700_, _06699_, _01602_);
  nor (_06701_, _06700_, _06695_);
  nor (_06702_, _05647_, _06680_);
  nor (_06703_, _06702_, _06669_);
  nor (_06704_, _06703_, _01923_);
  or (_06705_, _06704_, _02019_);
  nor (_06706_, _06705_, _06701_);
  nor (_06707_, _06706_, _06672_);
  or (_06708_, _06707_, _02018_);
  and (_06709_, _05662_, _04177_);
  or (_06710_, _06709_, _06669_);
  or (_06711_, _06710_, _05049_);
  and (_06712_, _06711_, _02136_);
  and (_06713_, _06712_, _06708_);
  and (_06714_, _05676_, _04177_);
  nor (_06715_, _06714_, _06669_);
  nor (_06716_, _06715_, _02136_);
  nor (_06717_, _06716_, _06713_);
  nor (_06718_, _06717_, _02039_);
  nor (_06719_, _06669_, _05687_);
  not (_06720_, _06719_);
  nor (_06721_, _06671_, _05076_);
  and (_06722_, _06721_, _06720_);
  nor (_06723_, _06722_, _06718_);
  nor (_06724_, _06723_, _02130_);
  or (_06725_, _06719_, _02131_);
  nor (_06726_, _06725_, _06674_);
  or (_06727_, _06726_, _02016_);
  nor (_06728_, _06727_, _06724_);
  nor (_06729_, _05659_, _06680_);
  nor (_06730_, _06729_, _06669_);
  and (_06731_, _06730_, _02016_);
  nor (_06732_, _06731_, _06728_);
  and (_06733_, _06732_, _05474_);
  nor (_06734_, _05673_, _06680_);
  nor (_06735_, _06734_, _06669_);
  nor (_06736_, _06735_, _05474_);
  or (_06737_, _06736_, _06733_);
  and (_06738_, _06737_, _02168_);
  nor (_06739_, _06682_, _02168_);
  or (_06740_, _06739_, _01594_);
  nor (_06741_, _06740_, _06738_);
  and (_06742_, _05759_, _04177_);
  nor (_06743_, _06742_, _06669_);
  and (_06744_, _06743_, _01594_);
  nor (_06745_, _06744_, _06741_);
  or (_06746_, _06745_, _26506_);
  or (_06747_, _26505_, \oc8051_golden_model_1.PCON [7]);
  and (_06748_, _06747_, _25964_);
  and (_25323_, _06748_, _06746_);
  or (_06749_, _05092_, rst);
  nor (_25324_, _06749_, _26505_);
  and (_06750_, _26505_, _25964_);
  nor (_06751_, \oc8051_golden_model_1.P3 [7], rst);
  nor (_25325_, _06751_, _06750_);
  nor (_06752_, \oc8051_golden_model_1.P2 [7], rst);
  nor (_25326_, _06752_, _06750_);
  nor (_06753_, \oc8051_golden_model_1.P1 [7], rst);
  nor (_25328_, _06753_, _06750_);
  nor (_06754_, \oc8051_golden_model_1.P0 [7], rst);
  nor (_25330_, _06754_, _06750_);
  not (_06755_, \oc8051_golden_model_1.IP [7]);
  nor (_06756_, _04155_, _06755_);
  not (_06757_, _04155_);
  nor (_06758_, _06757_, _02786_);
  nor (_06759_, _06758_, _06756_);
  and (_06760_, _06759_, _04950_);
  nor (_06761_, _05174_, _06755_);
  not (_06762_, _06761_);
  and (_06763_, _06762_, _06222_);
  and (_06764_, _06224_, _05174_);
  nor (_06765_, _06764_, _06761_);
  or (_06766_, _06765_, _04885_);
  nor (_06767_, _06766_, _06763_);
  nor (_06768_, _05499_, _06757_);
  nor (_06769_, _06768_, _06756_);
  and (_06770_, _06769_, _01969_);
  and (_06771_, _04155_, \oc8051_golden_model_1.ACC [7]);
  nor (_06772_, _06771_, _06756_);
  nor (_06773_, _06772_, _05488_);
  nor (_06774_, _04571_, _06755_);
  or (_06775_, _06774_, _01969_);
  nor (_06776_, _06775_, _06773_);
  or (_06777_, _06776_, _06233_);
  nor (_06778_, _06777_, _06770_);
  nor (_06779_, _06759_, _05487_);
  nor (_06780_, _06765_, _02223_);
  nor (_06781_, _06780_, _06779_);
  nand (_06782_, _06781_, _01964_);
  or (_06783_, _06782_, _06778_);
  nand (_06784_, _06772_, _01963_);
  and (_06785_, _06784_, _06783_);
  and (_06786_, _06785_, _06229_);
  and (_06787_, _06250_, _05174_);
  nor (_06788_, _06787_, _06761_);
  nor (_06789_, _06788_, _06229_);
  or (_06790_, _06789_, _06786_);
  and (_06791_, _06790_, _04885_);
  nor (_06792_, _06791_, _06767_);
  nor (_06793_, _06792_, _01924_);
  not (_06794_, _05174_);
  nor (_06795_, _06262_, _06794_);
  nor (_06796_, _06795_, _06761_);
  nor (_06797_, _06796_, _01925_);
  nor (_06798_, _06797_, _04950_);
  not (_06799_, _06798_);
  nor (_06800_, _06799_, _06793_);
  nor (_06801_, _06800_, _06760_);
  nor (_06802_, _06801_, _04951_);
  and (_06803_, _04155_, _03796_);
  nor (_06804_, _06756_, _05513_);
  not (_06805_, _06804_);
  nor (_06806_, _06805_, _06803_);
  nor (_06807_, _06806_, _01602_);
  not (_06808_, _06807_);
  nor (_06809_, _06808_, _06802_);
  nor (_06810_, _05647_, _06757_);
  nor (_06811_, _06810_, _06756_);
  nor (_06812_, _06811_, _01923_);
  or (_06813_, _06812_, _06278_);
  or (_06814_, _06813_, _06809_);
  and (_06815_, _05662_, _04155_);
  or (_06816_, _06756_, _05049_);
  or (_06817_, _06816_, _06815_);
  and (_06818_, _04155_, _02962_);
  nor (_06819_, _06818_, _06756_);
  and (_06820_, _06819_, _02019_);
  nor (_06821_, _06820_, _02135_);
  and (_06822_, _06821_, _06817_);
  and (_06823_, _06822_, _06814_);
  and (_06824_, _05676_, _04155_);
  nor (_06825_, _06824_, _06756_);
  nor (_06826_, _06825_, _02136_);
  nor (_06827_, _06826_, _06823_);
  nor (_06828_, _06827_, _02039_);
  nor (_06829_, _06756_, _05687_);
  not (_06830_, _06829_);
  nor (_06831_, _06819_, _05076_);
  and (_06832_, _06831_, _06830_);
  nor (_06833_, _06832_, _06828_);
  nor (_06834_, _06833_, _02130_);
  or (_06835_, _06829_, _02131_);
  nor (_06836_, _06835_, _06772_);
  or (_06837_, _06836_, _02016_);
  nor (_06838_, _06837_, _06834_);
  nor (_06839_, _05659_, _06757_);
  nor (_06840_, _06839_, _06756_);
  and (_06841_, _06840_, _02016_);
  nor (_06842_, _06841_, _06838_);
  and (_06843_, _06842_, _05474_);
  nor (_06844_, _05673_, _06757_);
  nor (_06845_, _06844_, _06756_);
  nor (_06846_, _06845_, _05474_);
  or (_06847_, _06846_, _06843_);
  and (_06848_, _06847_, _02168_);
  nor (_06849_, _06769_, _02168_);
  or (_06850_, _06849_, _02025_);
  or (_06851_, _06850_, _06848_);
  nand (_06852_, _06788_, _02025_);
  and (_06853_, _06852_, _06851_);
  nor (_06854_, _06853_, _01594_);
  and (_06855_, _05759_, _04155_);
  nor (_06856_, _06855_, _06756_);
  and (_06857_, _06856_, _01594_);
  nor (_06858_, _06857_, _06854_);
  or (_06859_, _06858_, _26506_);
  or (_06860_, _26505_, \oc8051_golden_model_1.IP [7]);
  and (_06861_, _06860_, _25964_);
  and (_25331_, _06861_, _06859_);
  not (_06862_, \oc8051_golden_model_1.IE [7]);
  nor (_06863_, _04183_, _06862_);
  not (_06864_, _04183_);
  nor (_06865_, _06864_, _02786_);
  nor (_06866_, _06865_, _06863_);
  and (_06867_, _06866_, _04950_);
  nor (_06868_, _05186_, _06862_);
  not (_06869_, _06868_);
  and (_06870_, _06869_, _06222_);
  and (_06871_, _06224_, _05186_);
  nor (_06872_, _06871_, _06868_);
  or (_06873_, _06872_, _04885_);
  nor (_06874_, _06873_, _06870_);
  nor (_06875_, _05499_, _06864_);
  nor (_06876_, _06875_, _06863_);
  and (_06877_, _06876_, _01969_);
  and (_06878_, _04183_, \oc8051_golden_model_1.ACC [7]);
  nor (_06879_, _06878_, _06863_);
  nor (_06880_, _06879_, _05488_);
  nor (_06881_, _04571_, _06862_);
  or (_06882_, _06881_, _01969_);
  nor (_06883_, _06882_, _06880_);
  or (_06884_, _06883_, _06233_);
  nor (_06885_, _06884_, _06877_);
  nor (_06886_, _06866_, _05487_);
  nor (_06887_, _06872_, _02223_);
  nor (_06888_, _06887_, _06886_);
  nand (_06889_, _06888_, _01964_);
  or (_06890_, _06889_, _06885_);
  nand (_06891_, _06879_, _01963_);
  and (_06892_, _06891_, _06890_);
  and (_06893_, _06892_, _06229_);
  and (_06894_, _06250_, _05186_);
  nor (_06895_, _06894_, _06868_);
  nor (_06896_, _06895_, _06229_);
  or (_06897_, _06896_, _06893_);
  and (_06898_, _06897_, _04885_);
  nor (_06899_, _06898_, _06874_);
  nor (_06900_, _06899_, _01924_);
  not (_06901_, _05186_);
  nor (_06902_, _06262_, _06901_);
  nor (_06903_, _06902_, _06868_);
  nor (_06904_, _06903_, _01925_);
  nor (_06905_, _06904_, _04950_);
  not (_06906_, _06905_);
  nor (_06907_, _06906_, _06900_);
  nor (_06908_, _06907_, _06867_);
  nor (_06909_, _06908_, _04951_);
  and (_06910_, _04183_, _03796_);
  nor (_06911_, _06863_, _05513_);
  not (_06912_, _06911_);
  nor (_06913_, _06912_, _06910_);
  nor (_06914_, _06913_, _01602_);
  not (_06915_, _06914_);
  nor (_06916_, _06915_, _06909_);
  nor (_06917_, _05647_, _06864_);
  nor (_06918_, _06917_, _06863_);
  nor (_06919_, _06918_, _01923_);
  or (_06920_, _06919_, _06278_);
  or (_06921_, _06920_, _06916_);
  and (_06922_, _05662_, _04183_);
  or (_06923_, _06863_, _05049_);
  or (_06924_, _06923_, _06922_);
  and (_06925_, _04183_, _02962_);
  nor (_06926_, _06925_, _06863_);
  and (_06927_, _06926_, _02019_);
  nor (_06928_, _06927_, _02135_);
  and (_06929_, _06928_, _06924_);
  and (_06930_, _06929_, _06921_);
  and (_06931_, _05676_, _04183_);
  nor (_06932_, _06931_, _06863_);
  nor (_06933_, _06932_, _02136_);
  nor (_06934_, _06933_, _06930_);
  nor (_06935_, _06934_, _02039_);
  nor (_06936_, _06863_, _05687_);
  not (_06937_, _06936_);
  nor (_06938_, _06926_, _05076_);
  and (_06939_, _06938_, _06937_);
  nor (_06940_, _06939_, _06935_);
  nor (_06941_, _06940_, _02130_);
  or (_06942_, _06936_, _02131_);
  nor (_06943_, _06942_, _06879_);
  or (_06944_, _06943_, _02016_);
  nor (_06945_, _06944_, _06941_);
  nor (_06946_, _05659_, _06864_);
  nor (_06947_, _06946_, _06863_);
  and (_06948_, _06947_, _02016_);
  nor (_06949_, _06948_, _06945_);
  and (_06950_, _06949_, _05474_);
  nor (_06951_, _05673_, _06864_);
  nor (_06952_, _06951_, _06863_);
  nor (_06953_, _06952_, _05474_);
  or (_06954_, _06953_, _06950_);
  and (_06955_, _06954_, _02168_);
  nor (_06956_, _06876_, _02168_);
  or (_06957_, _06956_, _02025_);
  or (_06958_, _06957_, _06955_);
  nand (_06959_, _06895_, _02025_);
  and (_06960_, _06959_, _06958_);
  nor (_06961_, _06960_, _01594_);
  and (_06962_, _05759_, _04183_);
  nor (_06963_, _06962_, _06863_);
  and (_06964_, _06963_, _01594_);
  nor (_06965_, _06964_, _06961_);
  or (_06966_, _06965_, _26506_);
  or (_06967_, _26505_, \oc8051_golden_model_1.IE [7]);
  and (_06968_, _06967_, _25964_);
  and (_25333_, _06968_, _06966_);
  or (_06969_, _04987_, rst);
  nor (_25334_, _06969_, _26505_);
  nand (_06970_, \oc8051_golden_model_1.DPL [7], _25964_);
  nor (_25335_, _06970_, _26505_);
  or (_06971_, _05671_, rst);
  nor (_25336_, _06971_, _26505_);
  nand (_06972_, \oc8051_golden_model_1.B [7], _25964_);
  nor (_25338_, _06972_, _26505_);
  and (_06973_, _02025_, _01853_);
  not (_06974_, _06973_);
  and (_06975_, _01660_, _02441_);
  and (_06976_, _02019_, _01853_);
  and (_06977_, _06976_, _02478_);
  and (_06978_, _01953_, _02441_);
  and (_06979_, _01957_, _01853_);
  not (_06980_, _06979_);
  and (_06981_, _02450_, _01959_);
  and (_06982_, _01959_, _01853_);
  and (_06983_, _02857_, _02412_);
  nor (_06984_, _04715_, _06983_);
  or (_06985_, _06984_, _03334_);
  and (_06986_, _01969_, _01853_);
  not (_06987_, _06986_);
  and (_06988_, _04571_, _01853_);
  nor (_06989_, _02857_, _01624_);
  not (_06990_, _06989_);
  nor (_06991_, _06990_, _02446_);
  nor (_06992_, _06991_, _06988_);
  and (_06993_, _06988_, _02478_);
  or (_06994_, _06993_, _04568_);
  or (_06995_, _06994_, _06992_);
  nor (_06996_, _01625_, _02441_);
  and (_06997_, _04557_, _01414_);
  nor (_06998_, _06997_, _06996_);
  and (_06999_, _06998_, _06995_);
  and (_07000_, _06999_, _06987_);
  and (_07001_, _07000_, _06985_);
  and (_07002_, _06986_, _02478_);
  nor (_07003_, _07002_, _07001_);
  nor (_07004_, _07003_, _06982_);
  nor (_07005_, _07004_, _06981_);
  nor (_07006_, _01621_, _02441_);
  nor (_07007_, _07006_, _07005_);
  and (_07008_, _01967_, _01853_);
  and (_07009_, _07008_, _02409_);
  nor (_07010_, _07009_, _02447_);
  and (_07011_, _07010_, _07007_);
  and (_07012_, _02857_, _01952_);
  and (_07013_, _07012_, _03917_);
  not (_07014_, _07013_);
  nand (_07015_, _07014_, _07011_);
  and (_07016_, _01963_, _01853_);
  and (_07017_, _07016_, _02409_);
  nor (_07018_, _07017_, _07015_);
  and (_07019_, _07018_, _06980_);
  or (_07020_, _07019_, _02459_);
  and (_07021_, _07020_, _02457_);
  nor (_07022_, _07021_, _06978_);
  and (_07023_, _01946_, _01853_);
  and (_07024_, _07023_, _03188_);
  nor (_07025_, _07024_, _07022_);
  nor (_07026_, _02446_, _01617_);
  nor (_07027_, _01632_, _02441_);
  nor (_07028_, _07027_, _07026_);
  and (_07029_, _07028_, _07025_);
  and (_07030_, _03917_, _03273_);
  nor (_07031_, _07030_, _02217_);
  and (_07032_, _07031_, _07029_);
  nor (_07033_, _07032_, _02482_);
  nor (_07034_, _07033_, _01606_);
  and (_07035_, _01606_, _02441_);
  nor (_07036_, _07035_, _07034_);
  and (_07037_, _04951_, _01853_);
  and (_07038_, _01853_, _01601_);
  and (_07039_, _07038_, _01382_);
  nor (_07040_, _07039_, _07037_);
  and (_07041_, _01853_, _01602_);
  not (_07042_, _07041_);
  and (_07043_, _07042_, _07040_);
  nor (_07044_, _07043_, _02478_);
  nor (_07045_, _02446_, _02856_);
  nor (_07046_, _07045_, _07044_);
  not (_07047_, _07046_);
  nor (_07048_, _07047_, _07036_);
  and (_07049_, _02857_, _01649_);
  and (_07050_, _07049_, _03917_);
  nor (_07051_, _07050_, _06976_);
  and (_07052_, _07051_, _07048_);
  nor (_07053_, _07052_, _06977_);
  nor (_07054_, _07053_, _01650_);
  and (_07055_, _01650_, _02441_);
  nor (_07056_, _07055_, _07054_);
  and (_07057_, _02130_, _01853_);
  not (_07058_, _07057_);
  and (_07059_, _02039_, _01853_);
  not (_07060_, _07059_);
  and (_07061_, _02018_, _01853_);
  and (_07062_, _02135_, _01853_);
  nor (_07063_, _07062_, _07061_);
  and (_07064_, _07063_, _07060_);
  and (_07065_, _07064_, _07058_);
  nor (_07066_, _07065_, _02478_);
  nor (_07067_, _07066_, _01666_);
  not (_07068_, _07067_);
  nor (_07069_, _07068_, _07056_);
  and (_07070_, _01666_, _02441_);
  nor (_07071_, _07070_, _07069_);
  nand (_07072_, _02128_, _01853_);
  nor (_07073_, _07072_, _02478_);
  nor (_07074_, _07073_, _01660_);
  not (_07075_, _07074_);
  nor (_07076_, _07075_, _07071_);
  nor (_07077_, _07076_, _06975_);
  nor (_07078_, _02446_, _02560_);
  nor (_07079_, _07078_, _07077_);
  and (_07080_, _02164_, _01853_);
  and (_07081_, _05417_, _03917_);
  nor (_07082_, _07081_, _07080_);
  and (_07083_, _07082_, _07079_);
  and (_07084_, _07080_, _02478_);
  nor (_07085_, _07084_, _07083_);
  nor (_07086_, _06466_, _02441_);
  nor (_07087_, _07086_, _07085_);
  and (_07088_, _07087_, _06974_);
  nor (_07089_, _07088_, _02567_);
  nor (_07090_, _02446_, _02569_);
  nor (_07091_, _07090_, _07089_);
  and (_07092_, _05441_, _03917_);
  not (_07093_, _07092_);
  and (_07094_, _07093_, _07091_);
  and (_07095_, _01853_, _01594_);
  and (_07096_, _07095_, _02409_);
  not (_07097_, _07096_);
  and (_07098_, _07097_, _07094_);
  not (_07099_, _06750_);
  nor (_07100_, _07008_, _06988_);
  nor (_07101_, _07095_, _07016_);
  and (_07102_, _07101_, _07100_);
  and (_07103_, _07102_, _07040_);
  and (_07104_, _07103_, _07064_);
  and (_07105_, _07038_, _01593_);
  not (_07106_, _07105_);
  not (_07107_, _07072_);
  nor (_07108_, _01666_, _01650_);
  and (_07109_, _07108_, _01621_);
  and (_07110_, _07109_, _06394_);
  nor (_07111_, _02703_, _02569_);
  and (_07112_, _01938_, _01958_);
  and (_07113_, _07112_, _01608_);
  or (_07114_, _07113_, _07111_);
  and (_07115_, _01938_, _01669_);
  and (_07116_, _07115_, _01609_);
  and (_07117_, _04886_, _01589_);
  or (_07118_, _07117_, _07116_);
  or (_07119_, _07118_, _07114_);
  nand (_07120_, _04919_, _01669_);
  nor (_07121_, _01660_, _04568_);
  and (_07122_, _07121_, _06466_);
  nand (_07123_, _07122_, _07120_);
  nor (_07124_, _07123_, _07119_);
  nand (_07125_, _07124_, _07110_);
  nand (_07126_, _02434_, _01940_);
  and (_07127_, _01938_, _02412_);
  and (_07128_, _02703_, _01935_);
  nor (_07129_, _01935_, _01629_);
  nor (_07130_, _07129_, _01649_);
  nor (_07131_, _07130_, _07128_);
  or (_07132_, _07131_, _07127_);
  or (_07133_, _07132_, _07126_);
  or (_07134_, _01953_, _01936_);
  or (_07135_, _03273_, _02353_);
  or (_07136_, _07135_, _07134_);
  or (_07137_, _05441_, _02359_);
  or (_07138_, _05417_, _02347_);
  or (_07139_, _07138_, _07137_);
  or (_07140_, _07139_, _07136_);
  and (_07141_, _02321_, _02412_);
  or (_07143_, _06983_, _07141_);
  nor (_07144_, _01935_, _01927_);
  and (_07145_, _07144_, _02412_);
  and (_07146_, _04886_, _01649_);
  or (_07147_, _07146_, _07145_);
  or (_07148_, _07147_, _07143_);
  or (_07149_, _07049_, _04715_);
  and (_07150_, _01938_, _01952_);
  or (_07151_, _07150_, _07012_);
  or (_07152_, _07151_, _07149_);
  or (_07153_, _07152_, _07148_);
  or (_07154_, _07153_, _07140_);
  or (_07155_, _07154_, _07133_);
  or (_07156_, _07155_, _07125_);
  or (_07157_, _07156_, _02217_);
  nor (_07158_, _07157_, _07107_);
  and (_07159_, _07158_, _07106_);
  nor (_07160_, _07080_, _07057_);
  nor (_07161_, _07023_, _06986_);
  and (_07162_, _07161_, _07160_);
  nor (_07163_, _06976_, _06973_);
  nor (_07164_, _06979_, _06982_);
  and (_07165_, _07164_, _07163_);
  and (_07166_, _07165_, _07162_);
  and (_07167_, _07166_, _07159_);
  and (_07168_, _07167_, _07104_);
  nor (_07169_, _07168_, _07099_);
  not (_07170_, _07169_);
  and (_07171_, _07095_, _02644_);
  and (_07172_, _02610_, _02025_);
  and (_07173_, _03400_, _01660_);
  and (_07174_, _06976_, _02644_);
  and (_07175_, _02610_, _01957_);
  and (_07176_, _02610_, _01959_);
  and (_07177_, _06986_, _02644_);
  not (_07178_, _03393_);
  or (_07179_, _06984_, _07178_);
  and (_07180_, _02003_, _02412_);
  nor (_07181_, _07180_, _06988_);
  and (_07182_, _06988_, _02644_);
  or (_07183_, _07182_, _04568_);
  or (_07184_, _07183_, _07181_);
  nand (_07185_, _04557_, _01590_);
  nor (_07186_, _03400_, _01625_);
  and (_07187_, _06997_, _01926_);
  nor (_07188_, _07187_, _07186_);
  and (_07189_, _07188_, _07185_);
  and (_07190_, _07189_, _07184_);
  and (_07191_, _07190_, _06987_);
  and (_07192_, _07191_, _07179_);
  nor (_07193_, _07192_, _07177_);
  nor (_07194_, _07193_, _06982_);
  nor (_07195_, _07194_, _07176_);
  nor (_07196_, _03400_, _01621_);
  nor (_07197_, _07196_, _07195_);
  and (_07198_, _07008_, _02643_);
  and (_07199_, _02003_, _01952_);
  nor (_07200_, _07199_, _07198_);
  and (_07201_, _07200_, _07197_);
  and (_07202_, _07012_, _03393_);
  not (_07203_, _07202_);
  nand (_07204_, _07203_, _07201_);
  and (_07205_, _07016_, _02643_);
  nor (_07206_, _07205_, _07204_);
  and (_07207_, _07206_, _06980_);
  nor (_07208_, _07207_, _07175_);
  nor (_07209_, _07208_, _01953_);
  and (_07210_, _03400_, _01953_);
  nor (_07211_, _07210_, _07209_);
  and (_07212_, _07023_, _02606_);
  nor (_07213_, _07212_, _07211_);
  nor (_07214_, _03400_, _01632_);
  and (_07215_, _02003_, _01929_);
  nor (_07216_, _07215_, _07214_);
  and (_07217_, _07216_, _07213_);
  and (_07218_, _03393_, _03273_);
  nor (_07219_, _07218_, _02217_);
  and (_07220_, _07219_, _07217_);
  nor (_07221_, _07220_, _02608_);
  nor (_07222_, _07221_, _01606_);
  and (_07223_, _03400_, _01606_);
  nor (_07224_, _07223_, _07222_);
  nor (_07225_, _07043_, _02644_);
  and (_07226_, _02003_, _01649_);
  nor (_07227_, _07226_, _07225_);
  not (_07228_, _07227_);
  nor (_07229_, _07228_, _07224_);
  and (_07230_, _07049_, _03393_);
  nor (_07231_, _07230_, _06976_);
  and (_07232_, _07231_, _07229_);
  nor (_07233_, _07232_, _07174_);
  nor (_07234_, _07233_, _01650_);
  and (_07235_, _03400_, _01650_);
  nor (_07236_, _07235_, _07234_);
  nor (_07237_, _07065_, _02644_);
  nor (_07238_, _07237_, _01666_);
  not (_07239_, _07238_);
  nor (_07240_, _07239_, _07236_);
  and (_07241_, _03400_, _01666_);
  nor (_07242_, _07241_, _07240_);
  nor (_07243_, _07072_, _02644_);
  nor (_07244_, _07243_, _01660_);
  not (_07245_, _07244_);
  nor (_07246_, _07245_, _07242_);
  nor (_07247_, _07246_, _07173_);
  and (_07248_, _02003_, _01669_);
  nor (_07249_, _07248_, _07247_);
  and (_07250_, _05417_, _03393_);
  nor (_07251_, _07250_, _07080_);
  and (_07252_, _07251_, _07249_);
  and (_07253_, _07080_, _02644_);
  nor (_07254_, _07253_, _07252_);
  nor (_07255_, _06466_, _03400_);
  nor (_07256_, _07255_, _06973_);
  not (_07257_, _07256_);
  nor (_07258_, _07257_, _07254_);
  nor (_07259_, _07258_, _07172_);
  and (_07260_, _02003_, _01589_);
  nor (_07261_, _07260_, _07259_);
  and (_07262_, _05441_, _03393_);
  nor (_07263_, _07262_, _07095_);
  and (_07264_, _07263_, _07261_);
  nor (_07265_, _07264_, _07171_);
  nor (_07266_, _07265_, _07170_);
  and (_07267_, _07266_, _07098_);
  and (_07268_, _05441_, _03473_);
  and (_07269_, _05417_, _03473_);
  not (_07270_, _01606_);
  not (_07271_, _02217_);
  and (_07272_, _03473_, _03273_);
  and (_07273_, _03399_, \oc8051_golden_model_1.SP [2]);
  nor (_07274_, _07273_, \oc8051_golden_model_1.SP [3]);
  nor (_07275_, _07274_, _06384_);
  not (_07276_, _07275_);
  nor (_07277_, _07276_, _01632_);
  and (_07278_, _07012_, _03473_);
  nor (_07279_, _07276_, _01625_);
  nor (_07280_, _06983_, \oc8051_golden_model_1.PSW [3]);
  and (_07281_, _06983_, _03473_);
  or (_07282_, _07281_, _06988_);
  nor (_07283_, _07282_, _07280_);
  and (_07284_, _04571_, _02450_);
  nor (_07285_, _07284_, _07283_);
  nor (_07286_, _07285_, _04568_);
  or (_07287_, _07286_, _04715_);
  nor (_07288_, _07287_, _07279_);
  and (_07289_, _04715_, _03473_);
  nor (_07290_, _07289_, _06986_);
  not (_07291_, _07290_);
  nor (_07292_, _07291_, _07288_);
  and (_07293_, _02450_, _01969_);
  or (_07294_, _07293_, _06982_);
  nor (_07295_, _07294_, _07292_);
  and (_07296_, _06982_, _01885_);
  nor (_07297_, _07296_, _07295_);
  nor (_07298_, _07297_, _06363_);
  nor (_07299_, _07275_, _01621_);
  nor (_07300_, _07299_, _07008_);
  not (_07301_, _07300_);
  nor (_07302_, _07301_, _07298_);
  and (_07303_, _07008_, _01916_);
  or (_07304_, _07303_, _07012_);
  nor (_07305_, _07304_, _07302_);
  or (_07306_, _07305_, _07016_);
  nor (_07307_, _07306_, _07278_);
  and (_07308_, _07016_, _01916_);
  or (_07309_, _07308_, _06979_);
  nor (_07310_, _07309_, _07307_);
  nor (_07311_, _01953_, _01885_);
  nor (_07312_, _07311_, _02455_);
  nor (_07313_, _07312_, _07310_);
  and (_07314_, _07275_, _01953_);
  nor (_07315_, _07314_, _07313_);
  nor (_07316_, _07315_, _07023_);
  and (_07317_, _07023_, _01918_);
  or (_07318_, _07317_, _07316_);
  and (_07319_, _07318_, _01632_);
  or (_07320_, _07319_, _03273_);
  nor (_07321_, _07320_, _07277_);
  nor (_07322_, _07321_, _07272_);
  and (_07323_, _07322_, _07271_);
  and (_07324_, _02217_, _03683_);
  or (_07325_, _07324_, _07323_);
  and (_07326_, _07325_, _07270_);
  and (_07327_, _07275_, _01606_);
  not (_07328_, _07327_);
  and (_07329_, _07328_, _07043_);
  not (_07330_, _07329_);
  nor (_07331_, _07330_, _07326_);
  nor (_07332_, _07043_, _01916_);
  nor (_07333_, _07332_, _07331_);
  nor (_07334_, _07333_, _07049_);
  and (_07335_, _07049_, _03473_);
  nor (_07336_, _07335_, _06976_);
  not (_07337_, _07336_);
  nor (_07338_, _07337_, _07334_);
  and (_07339_, _02450_, _02019_);
  nor (_07340_, _07339_, _07338_);
  nor (_07341_, _07340_, _01650_);
  and (_07342_, _07275_, _01650_);
  not (_07343_, _07342_);
  and (_07344_, _07343_, _07065_);
  not (_07345_, _07344_);
  nor (_07346_, _07345_, _07341_);
  nor (_07347_, _07065_, _01916_);
  nor (_07348_, _07347_, _01666_);
  not (_07349_, _07348_);
  nor (_07350_, _07349_, _07346_);
  and (_07351_, _07275_, _01666_);
  nor (_07352_, _07351_, _07107_);
  not (_07353_, _07352_);
  nor (_07354_, _07353_, _07350_);
  nor (_07355_, _07072_, _01916_);
  nor (_07356_, _07355_, _01660_);
  not (_07357_, _07356_);
  nor (_07358_, _07357_, _07354_);
  and (_07359_, _07275_, _01660_);
  nor (_07360_, _07359_, _05417_);
  not (_07361_, _07360_);
  nor (_07362_, _07361_, _07358_);
  or (_07363_, _07362_, _07080_);
  nor (_07364_, _07363_, _07269_);
  and (_07365_, _07080_, _01916_);
  nor (_07366_, _07365_, _06467_);
  not (_07367_, _07366_);
  nor (_07368_, _07367_, _07364_);
  nor (_07369_, _07275_, _06466_);
  nor (_07370_, _07369_, _06973_);
  not (_07371_, _07370_);
  nor (_07372_, _07371_, _07368_);
  and (_07373_, _06973_, _03683_);
  or (_07374_, _07373_, _05441_);
  nor (_07375_, _07374_, _07372_);
  or (_07376_, _07375_, _07095_);
  nor (_07377_, _07376_, _07268_);
  and (_07378_, _07095_, _01916_);
  nor (_07379_, _07378_, _07377_);
  and (_07380_, _02221_, _02025_);
  nor (_07381_, _03399_, \oc8051_golden_model_1.SP [2]);
  nor (_07382_, _07381_, _07273_);
  and (_07383_, _07382_, _01660_);
  and (_07384_, _06976_, _02264_);
  and (_07385_, _02221_, _01957_);
  and (_07386_, _02221_, _01959_);
  and (_07387_, _06986_, _02264_);
  not (_07388_, _03272_);
  or (_07389_, _06984_, _07388_);
  nor (_07390_, _06988_, _07127_);
  and (_07391_, _06988_, _02264_);
  or (_07392_, _07391_, _04568_);
  or (_07393_, _07392_, _07390_);
  nor (_07394_, _07382_, _01625_);
  nor (_07395_, _07394_, _07112_);
  and (_07396_, _07395_, _07393_);
  and (_07397_, _07396_, _06987_);
  and (_07398_, _07397_, _07389_);
  nor (_07399_, _07398_, _07387_);
  nor (_07400_, _07399_, _06982_);
  nor (_07401_, _07400_, _07386_);
  nor (_07402_, _07382_, _01621_);
  nor (_07403_, _07402_, _07401_);
  and (_07404_, _07008_, _02263_);
  nor (_07405_, _07404_, _07150_);
  and (_07406_, _07405_, _07403_);
  and (_07407_, _07012_, _03272_);
  not (_07408_, _07407_);
  and (_07409_, _07408_, _07406_);
  and (_07410_, _07016_, _02263_);
  nor (_07411_, _07410_, _06979_);
  and (_07412_, _07411_, _07409_);
  nor (_07413_, _07412_, _07385_);
  nor (_07414_, _07413_, _01953_);
  and (_07415_, _07382_, _01953_);
  nor (_07416_, _07415_, _07414_);
  and (_07417_, _07023_, _02214_);
  nor (_07418_, _07417_, _07416_);
  nor (_07419_, _07382_, _01632_);
  nor (_07420_, _07419_, _01941_);
  and (_07421_, _07420_, _07418_);
  and (_07422_, _03273_, _03272_);
  nor (_07423_, _07422_, _02217_);
  and (_07424_, _07423_, _07421_);
  nor (_07425_, _07424_, _02218_);
  nor (_07426_, _07425_, _01606_);
  and (_07427_, _07382_, _01606_);
  nor (_07428_, _07427_, _07426_);
  nor (_07429_, _07043_, _02264_);
  and (_07430_, _01938_, _01649_);
  nor (_07431_, _07430_, _07429_);
  not (_07432_, _07431_);
  nor (_07433_, _07432_, _07428_);
  and (_07434_, _07049_, _03272_);
  nor (_07435_, _07434_, _06976_);
  and (_07436_, _07435_, _07433_);
  nor (_07437_, _07436_, _07384_);
  nor (_07438_, _07437_, _01650_);
  and (_07439_, _07382_, _01650_);
  nor (_07440_, _07439_, _07438_);
  nor (_07441_, _07065_, _02264_);
  nor (_07442_, _07441_, _01666_);
  not (_07443_, _07442_);
  nor (_07444_, _07443_, _07440_);
  and (_07445_, _07382_, _01666_);
  nor (_07446_, _07445_, _07444_);
  nor (_07447_, _07072_, _02264_);
  nor (_07448_, _07447_, _01660_);
  not (_07449_, _07448_);
  nor (_07450_, _07449_, _07446_);
  nor (_07451_, _07450_, _07383_);
  nor (_07452_, _07451_, _07115_);
  and (_07453_, _05417_, _03272_);
  nor (_07454_, _07453_, _07080_);
  and (_07455_, _07454_, _07452_);
  and (_07456_, _07080_, _02264_);
  nor (_07457_, _07456_, _07455_);
  nor (_07458_, _07382_, _06466_);
  nor (_07459_, _07458_, _06973_);
  not (_07460_, _07459_);
  nor (_07461_, _07460_, _07457_);
  nor (_07462_, _07461_, _07380_);
  nor (_07463_, _07462_, _05443_);
  and (_07464_, _05441_, _03272_);
  nor (_07465_, _07464_, _07095_);
  and (_07466_, _07465_, _07463_);
  and (_07467_, _07095_, _02264_);
  nor (_07468_, _07467_, _07466_);
  nor (_07469_, _07468_, _07170_);
  not (_07470_, _07469_);
  nor (_07471_, _07470_, _07379_);
  and (_07472_, _07471_, _07267_);
  or (_07473_, _07472_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_07474_, _07122_, _07110_);
  nor (_07475_, _07474_, _07099_);
  and (_07476_, _07475_, \oc8051_golden_model_1.SP [0]);
  and (_07477_, _07476_, _02717_);
  and (_07478_, \oc8051_golden_model_1.SP [1], _02441_);
  and (_07479_, _07478_, \oc8051_golden_model_1.SP [2]);
  nor (_07480_, _07478_, _07382_);
  nor (_07481_, _07480_, _07479_);
  and (_07482_, _06351_, _02441_);
  nor (_07483_, _07479_, _07275_);
  nor (_07484_, _07483_, _07482_);
  and (_07485_, _07484_, _07475_);
  and (_07486_, _07485_, _07481_);
  and (_07487_, _07486_, _07477_);
  not (_07488_, _07487_);
  and (_07489_, _07488_, _07473_);
  not (_07490_, _07472_);
  and (_07491_, _07095_, _05759_);
  not (_07492_, _02786_);
  not (_07493_, _04074_);
  not (_07494_, _03976_);
  not (_07495_, _04024_);
  not (_07496_, _03473_);
  nor (_07497_, _03393_, _03917_);
  and (_07498_, _07497_, _07388_);
  and (_07499_, _07498_, _07496_);
  and (_07500_, _07499_, _07495_);
  and (_07501_, _07500_, _07494_);
  and (_07502_, _07501_, _07493_);
  nor (_07503_, _07502_, _07492_);
  and (_07504_, _07502_, _07492_);
  nor (_07505_, _07504_, _07503_);
  nor (_07506_, _07505_, _05444_);
  nand (_07507_, _04623_, _01650_);
  nor (_07508_, _02859_, _02019_);
  or (_07509_, _07508_, _02220_);
  nor (_07510_, _06262_, _07271_);
  nand (_07511_, _04779_, _01950_);
  or (_07512_, _06250_, _06980_);
  not (_07513_, _06982_);
  or (_07514_, _06224_, _07513_);
  not (_07515_, _04715_);
  or (_07516_, _07515_, _03796_);
  and (_07517_, _03393_, _03917_);
  and (_07518_, _07517_, _04701_);
  and (_07519_, _07518_, _04702_);
  and (_07520_, _07519_, _04074_);
  and (_07521_, _07520_, _02786_);
  nor (_07522_, _07520_, _02786_);
  or (_07523_, _07522_, _07521_);
  and (_07524_, _07523_, _04557_);
  and (_07525_, _01625_, \oc8051_golden_model_1.ACC [7]);
  nor (_07526_, _04623_, _01625_);
  or (_07527_, _07526_, _07525_);
  and (_07528_, _07527_, _04709_);
  or (_07529_, _07528_, _04715_);
  or (_07530_, _07529_, _07524_);
  and (_07531_, _07530_, _07516_);
  or (_07532_, _07531_, _06986_);
  nand (_07533_, _06986_, _05499_);
  and (_07534_, _07533_, _07532_);
  or (_07535_, _07534_, _06982_);
  and (_07536_, _07535_, _07514_);
  or (_07537_, _07536_, _06363_);
  nor (_07538_, _04622_, _01621_);
  nor (_07539_, _07538_, _07008_);
  and (_07540_, _07539_, _07537_);
  and (_07541_, _07008_, _07492_);
  or (_07542_, _07541_, _06979_);
  or (_07543_, _07542_, _07540_);
  and (_07544_, _07543_, _07512_);
  or (_07545_, _07544_, _01953_);
  not (_07546_, _07023_);
  nand (_07547_, _04779_, _01953_);
  and (_07548_, _07547_, _07546_);
  and (_07549_, _07548_, _07545_);
  nand (_07550_, _07023_, _06224_);
  nor (_07551_, _07550_, _06222_);
  or (_07552_, _07551_, _07549_);
  and (_07553_, _07552_, _01632_);
  or (_07554_, _04623_, _01632_);
  nand (_07555_, _07554_, _01942_);
  or (_07556_, _07555_, _07553_);
  and (_07557_, _07556_, _07511_);
  or (_07558_, _07557_, _03273_);
  and (_07559_, _04778_, _03273_);
  nand (_07560_, _07559_, _03798_);
  and (_07561_, _07560_, _07271_);
  and (_07562_, _07561_, _07558_);
  or (_07563_, _07562_, _07510_);
  and (_07564_, _07563_, _07270_);
  and (_07565_, _04622_, _01606_);
  or (_07566_, _07565_, _07039_);
  or (_07567_, _07566_, _07564_);
  nand (_07568_, _07039_, _02786_);
  and (_07569_, _07568_, _07567_);
  or (_07570_, _07569_, _07037_);
  not (_07571_, _07037_);
  or (_07572_, _07571_, _03796_);
  and (_07573_, _07572_, _07106_);
  and (_07574_, _07573_, _07570_);
  nor (_07575_, _07042_, _05647_);
  or (_07576_, _07575_, _02859_);
  or (_07577_, _07576_, _07574_);
  and (_07578_, _07577_, _07509_);
  and (_07579_, _06976_, _02962_);
  or (_07580_, _07579_, _01650_);
  or (_07581_, _07580_, _07578_);
  and (_07582_, _07581_, _07507_);
  or (_07583_, _07582_, _07061_);
  not (_07584_, _07062_);
  not (_07585_, _07061_);
  or (_07586_, _07585_, _05662_);
  and (_07587_, _07586_, _07584_);
  and (_07588_, _07587_, _07583_);
  and (_07589_, _07062_, _05676_);
  or (_07590_, _07589_, _07059_);
  or (_07591_, _07590_, _07588_);
  or (_07592_, _07060_, _05661_);
  and (_07593_, _07592_, _07058_);
  and (_07594_, _07593_, _07591_);
  and (_07595_, _07057_, _05674_);
  or (_07596_, _07595_, _01666_);
  or (_07597_, _07596_, _07594_);
  and (_07598_, _02016_, _01853_);
  and (_07599_, _04623_, _01666_);
  nor (_07600_, _07599_, _07598_);
  and (_07601_, _07600_, _07597_);
  and (_07602_, _02126_, _01853_);
  not (_07603_, _07602_);
  nand (_07604_, _07603_, _05659_);
  and (_07605_, _07604_, _07107_);
  or (_07606_, _07605_, _07601_);
  nand (_07607_, _07602_, _05673_);
  and (_07608_, _07607_, _05157_);
  and (_07609_, _07608_, _07606_);
  or (_07610_, _07128_, _02560_);
  nand (_07611_, _04622_, _01660_);
  nand (_07612_, _07611_, _07610_);
  or (_07613_, _07612_, _07609_);
  and (_07614_, _04886_, _01669_);
  not (_07615_, _07614_);
  or (_07616_, _07523_, _07610_);
  and (_07617_, _07616_, _07615_);
  and (_07618_, _07617_, _07613_);
  and (_07619_, _07523_, _07614_);
  or (_07620_, _07619_, _05417_);
  or (_07621_, _07620_, _07618_);
  not (_07622_, _07080_);
  not (_07623_, _05417_);
  not (_07624_, _03796_);
  not (_07625_, _03748_);
  not (_07626_, _03850_);
  not (_07627_, _03903_);
  not (_07628_, _03516_);
  not (_07629_, _03564_);
  nor (_07630_, _03677_, _03613_);
  and (_07631_, _07630_, _07629_);
  and (_07632_, _07631_, _07628_);
  and (_07633_, _07632_, _07627_);
  and (_07634_, _07633_, _07626_);
  and (_07635_, _07634_, _07625_);
  nor (_07636_, _07635_, _07624_);
  and (_07637_, _07635_, _07624_);
  or (_07638_, _07637_, _07636_);
  or (_07639_, _07638_, _07623_);
  and (_07640_, _07639_, _07622_);
  and (_07641_, _07640_, _07621_);
  nor (_07642_, _07622_, _05499_);
  or (_07643_, _07642_, _02023_);
  or (_07644_, _07643_, _07641_);
  nand (_07645_, _02992_, _02023_);
  and (_07646_, _07645_, _07644_);
  or (_07647_, _07646_, _01670_);
  and (_07648_, _04623_, _01670_);
  nor (_07649_, _07648_, _06973_);
  and (_07650_, _07649_, _07647_);
  not (_07651_, _05444_);
  and (_07652_, _06259_, _06973_);
  nor (_07653_, _07652_, _07651_);
  not (_07654_, _07653_);
  nor (_07655_, _07654_, _07650_);
  nor (_07656_, _07655_, _07506_);
  nor (_07657_, _07656_, _05441_);
  and (_07658_, _03677_, _03613_);
  and (_07659_, _07658_, _03564_);
  and (_07660_, _07659_, _03516_);
  and (_07661_, _07660_, _03903_);
  and (_07662_, _07661_, _03850_);
  and (_07663_, _07662_, _03748_);
  nor (_07664_, _07663_, _03796_);
  and (_07665_, _07663_, _03796_);
  nor (_07666_, _07665_, _07664_);
  nor (_07667_, _07666_, _05442_);
  nor (_07668_, _07667_, _07095_);
  not (_07669_, _07668_);
  nor (_07670_, _07669_, _07657_);
  nor (_07671_, _07670_, _07491_);
  nor (_07672_, _07671_, _07170_);
  or (_07673_, _07672_, _07490_);
  and (_07674_, _07673_, _07489_);
  and (_07675_, _02851_, _05429_);
  and (_07676_, _02878_, _02023_);
  or (_07677_, _07676_, _07675_);
  and (_07678_, _07677_, _07475_);
  and (_07679_, _07678_, _07487_);
  or (_29689_, _07679_, _07674_);
  and (_07680_, _07481_, _07475_);
  nor (_07681_, _07485_, _07680_);
  and (_07682_, _07681_, _07475_);
  and (_07683_, _07682_, _07478_);
  not (_07684_, _07683_);
  nor (_07685_, _07379_, _07170_);
  nor (_07686_, _07685_, _07469_);
  and (_07687_, _07169_, _07098_);
  nor (_07688_, _07687_, _07266_);
  and (_07689_, _07688_, _07686_);
  and (_07690_, _07689_, _07169_);
  or (_07691_, _07690_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_07692_, _07691_, _07684_);
  not (_07693_, _07690_);
  and (_07694_, _07651_, _03917_);
  nand (_07695_, _01670_, _01325_);
  nor (_07696_, _04405_, \oc8051_golden_model_1.ACC [0]);
  nand (_07697_, _07696_, _07602_);
  and (_07698_, _04405_, _05531_);
  and (_07699_, _07698_, _07059_);
  not (_07700_, _07039_);
  or (_07701_, _07700_, _03334_);
  nand (_07702_, _04828_, _01950_);
  and (_07703_, _07008_, _03334_);
  or (_07704_, _03917_, _04709_);
  nor (_07705_, _01625_, _01325_);
  and (_07706_, _01625_, \oc8051_golden_model_1.ACC [0]);
  or (_07707_, _07706_, _07705_);
  nor (_07708_, _07707_, _04557_);
  nor (_07709_, _07708_, _06986_);
  and (_07710_, _07709_, _07704_);
  nor (_07711_, _06987_, _04405_);
  or (_07712_, _07711_, _07710_);
  and (_07713_, _07712_, _07513_);
  and (_07714_, _05191_, \oc8051_golden_model_1.P3 [0]);
  nor (_07715_, _07714_, _05296_);
  and (_07716_, _07715_, _05288_);
  and (_07717_, _05195_, \oc8051_golden_model_1.P1 [0]);
  and (_07718_, _05189_, \oc8051_golden_model_1.P2 [0]);
  and (_07719_, _04099_, \oc8051_golden_model_1.P0 [0]);
  or (_07720_, _07719_, _07718_);
  nor (_07721_, _07720_, _07717_);
  and (_07722_, _07721_, _05295_);
  and (_07723_, _07722_, _07716_);
  and (_07724_, _07723_, _04350_);
  nand (_07725_, _07724_, _05282_);
  and (_07726_, _07725_, _06982_);
  or (_07727_, _07726_, _06363_);
  or (_07728_, _07727_, _07713_);
  nor (_07729_, _01621_, \oc8051_golden_model_1.PC [0]);
  nor (_07730_, _07729_, _07008_);
  and (_07731_, _07730_, _07728_);
  or (_07732_, _07731_, _07703_);
  and (_07733_, _07732_, _06980_);
  or (_07734_, _04157_, _06980_);
  nor (_07735_, _07734_, _07724_);
  or (_07736_, _07735_, _01953_);
  or (_07737_, _07736_, _07733_);
  nand (_07738_, _04828_, _01953_);
  and (_07739_, _07738_, _07546_);
  and (_07740_, _07739_, _07737_);
  or (_07741_, _07724_, _05282_);
  and (_07742_, _07725_, _07023_);
  and (_07743_, _07742_, _07741_);
  or (_07744_, _07743_, _07740_);
  and (_07745_, _07744_, _01632_);
  or (_07746_, _01632_, _01325_);
  nand (_07747_, _01942_, _07746_);
  or (_07748_, _07747_, _07745_);
  and (_07749_, _07748_, _07702_);
  or (_07750_, _07749_, _03273_);
  and (_07751_, _03677_, _01853_);
  nand (_07752_, _04827_, _03273_);
  or (_07753_, _07752_, _07751_);
  and (_07754_, _07753_, _07750_);
  or (_07755_, _07754_, _02217_);
  nor (_07756_, _05304_, _04157_);
  and (_07757_, _04115_, \oc8051_golden_model_1.PSW [7]);
  and (_07758_, _07757_, _02263_);
  nor (_07759_, _07758_, _07756_);
  nand (_07760_, _07759_, _02217_);
  and (_07761_, _07760_, _07270_);
  and (_07762_, _07761_, _07755_);
  and (_07763_, _01606_, \oc8051_golden_model_1.PC [0]);
  or (_07764_, _07039_, _07763_);
  or (_07765_, _07764_, _07762_);
  and (_07766_, _07765_, _07701_);
  or (_07767_, _07766_, _07037_);
  or (_07768_, _07571_, _03677_);
  and (_07769_, _07768_, _07106_);
  and (_07770_, _07769_, _07767_);
  and (_07771_, _03334_, _02943_);
  and (_07772_, _05527_, \oc8051_golden_model_1.P1INREG [0]);
  and (_07773_, _05550_, \oc8051_golden_model_1.ACC [0]);
  nor (_07774_, _07773_, _07772_);
  and (_07775_, _05556_, \oc8051_golden_model_1.P0INREG [0]);
  and (_07776_, _05558_, \oc8051_golden_model_1.SCON [0]);
  nor (_07777_, _07776_, _07775_);
  and (_07778_, _07777_, _07774_);
  and (_07779_, _05534_, \oc8051_golden_model_1.SBUF [0]);
  and (_07780_, _05544_, \oc8051_golden_model_1.PSW [0]);
  nor (_07781_, _07780_, _07779_);
  and (_07782_, _05540_, \oc8051_golden_model_1.TCON [0]);
  and (_07783_, _05553_, \oc8051_golden_model_1.B [0]);
  nor (_07784_, _07783_, _07782_);
  and (_07785_, _07784_, _07781_);
  and (_07786_, _07785_, _07778_);
  and (_07787_, _05567_, \oc8051_golden_model_1.PCON [0]);
  and (_07788_, _05569_, \oc8051_golden_model_1.DPH [0]);
  nor (_07789_, _07788_, _07787_);
  and (_07790_, _07789_, _07786_);
  and (_07791_, _05578_, \oc8051_golden_model_1.TL1 [0]);
  and (_07792_, _05633_, \oc8051_golden_model_1.SP [0]);
  nor (_07793_, _07792_, _07791_);
  and (_07794_, _05576_, \oc8051_golden_model_1.DPL [0]);
  and (_07795_, _05629_, \oc8051_golden_model_1.TMOD [0]);
  nor (_07796_, _07795_, _07794_);
  and (_07797_, _07796_, _07793_);
  and (_07798_, _05582_, \oc8051_golden_model_1.TL0 [0]);
  not (_07799_, _07798_);
  and (_07800_, _05603_, \oc8051_golden_model_1.IE [0]);
  and (_07801_, _05619_, \oc8051_golden_model_1.IP [0]);
  nor (_07802_, _07801_, _07800_);
  and (_07803_, _05615_, \oc8051_golden_model_1.P2INREG [0]);
  and (_07804_, _05609_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_07805_, _07804_, _07803_);
  and (_07806_, _07805_, _07802_);
  and (_07807_, _07806_, _07799_);
  and (_07808_, _05595_, \oc8051_golden_model_1.TH1 [0]);
  and (_07809_, _05587_, \oc8051_golden_model_1.TH0 [0]);
  nor (_07810_, _07809_, _07808_);
  and (_07811_, _07810_, _07807_);
  and (_07812_, _07811_, _07797_);
  and (_07813_, _07812_, _07790_);
  not (_07814_, _07813_);
  nor (_07815_, _07814_, _07771_);
  nor (_07816_, _07815_, _07042_);
  or (_07817_, _07816_, _02859_);
  or (_07818_, _07817_, _07770_);
  and (_07819_, _02859_, _02409_);
  nor (_07820_, _07819_, _06976_);
  and (_07821_, _07820_, _07818_);
  and (_07822_, _06976_, _05531_);
  or (_07823_, _07822_, _01650_);
  or (_07824_, _07823_, _07821_);
  and (_07825_, _01650_, _01325_);
  nor (_07826_, _07825_, _07061_);
  and (_07827_, _07826_, _07824_);
  nor (_07828_, _04405_, _05531_);
  nor (_07829_, _07828_, _07698_);
  nor (_07830_, _07829_, _07062_);
  nor (_07831_, _07830_, _07063_);
  or (_07832_, _07831_, _07827_);
  and (_07833_, _04405_, \oc8051_golden_model_1.ACC [0]);
  nor (_07834_, _07833_, _07696_);
  or (_07835_, _07834_, _07584_);
  and (_07836_, _07835_, _07060_);
  and (_07837_, _07836_, _07832_);
  or (_07838_, _07837_, _07699_);
  and (_07839_, _07838_, _07058_);
  and (_07840_, _07833_, _07057_);
  or (_07841_, _07840_, _01666_);
  or (_07842_, _07841_, _07839_);
  and (_07843_, _01666_, _01325_);
  nor (_07844_, _07843_, _07598_);
  and (_07845_, _07844_, _07842_);
  nand (_07846_, _07828_, _07603_);
  and (_07847_, _07846_, _07107_);
  or (_07848_, _07847_, _07845_);
  and (_07849_, _07848_, _07697_);
  or (_07850_, _07849_, _01660_);
  nand (_07851_, _01660_, _01325_);
  and (_07852_, _07851_, _05415_);
  and (_07853_, _07852_, _07850_);
  and (_07854_, _05416_, _03917_);
  or (_07855_, _07854_, _07853_);
  and (_07856_, _07855_, _07623_);
  nor (_07857_, _07623_, _03677_);
  or (_07858_, _07857_, _07080_);
  or (_07859_, _07858_, _07856_);
  nand (_07860_, _07080_, _04405_);
  and (_07861_, _07860_, _05429_);
  and (_07862_, _07861_, _07859_);
  and (_07863_, _02023_, _01325_);
  or (_07864_, _07863_, _01670_);
  or (_07865_, _07864_, _07862_);
  and (_07866_, _07865_, _07695_);
  or (_07867_, _07866_, _06973_);
  or (_07868_, _07756_, _06974_);
  and (_07869_, _07868_, _05444_);
  and (_07870_, _07869_, _07867_);
  or (_07871_, _07870_, _07694_);
  and (_07872_, _07871_, _05442_);
  nor (_07873_, _05442_, _03677_);
  or (_07874_, _07873_, _07095_);
  or (_07875_, _07874_, _07872_);
  nand (_07876_, _07095_, _04405_);
  and (_07877_, _07876_, _07169_);
  and (_07878_, _07877_, _07875_);
  or (_07879_, _07878_, _07693_);
  and (_07880_, _07879_, _07692_);
  nor (_07881_, _04673_, _02023_);
  and (_07882_, _03141_, _02023_);
  or (_07883_, _07882_, _07881_);
  and (_07884_, _07883_, _07683_);
  or (_29636_, _07884_, _07880_);
  or (_07885_, _07690_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_07886_, _07885_, _07684_);
  nor (_07887_, _07658_, _07630_);
  or (_07888_, _07887_, _05442_);
  nor (_07889_, _07887_, _07623_);
  or (_07890_, _07116_, _02347_);
  nor (_07891_, _07517_, _07497_);
  nand (_07892_, _07891_, _07890_);
  nor (_07893_, _04452_, _02676_);
  and (_07894_, _07893_, _07059_);
  nand (_07895_, _07039_, _03393_);
  nand (_07896_, _04759_, _01950_);
  and (_07897_, _04099_, \oc8051_golden_model_1.P0 [1]);
  and (_07898_, _05189_, \oc8051_golden_model_1.P2 [1]);
  nor (_07899_, _07898_, _07897_);
  and (_07900_, _05195_, \oc8051_golden_model_1.P1 [1]);
  and (_07901_, _05191_, \oc8051_golden_model_1.P3 [1]);
  nor (_07902_, _07901_, _07900_);
  and (_07903_, _07902_, _07899_);
  and (_07904_, _07903_, _05216_);
  and (_07905_, _07904_, _05213_);
  and (_07906_, _07905_, _04406_);
  nor (_07907_, _07906_, _04110_);
  or (_07908_, _07907_, _06980_);
  nor (_07909_, _05743_, _05494_);
  nor (_07910_, _07909_, _06987_);
  nand (_07911_, _07891_, _04557_);
  nor (_07912_, _01625_, \oc8051_golden_model_1.PC [1]);
  and (_07913_, _01625_, \oc8051_golden_model_1.ACC [1]);
  or (_07914_, _07913_, _04557_);
  nor (_07915_, _07914_, _07912_);
  nor (_07916_, _07915_, _06986_);
  and (_07917_, _07916_, _07911_);
  or (_07918_, _07917_, _06982_);
  or (_07919_, _07918_, _07910_);
  nand (_07920_, _07906_, _05203_);
  or (_07921_, _07920_, _07513_);
  and (_07922_, _07921_, _07919_);
  or (_07923_, _07922_, _06363_);
  nor (_07924_, _01621_, _01298_);
  nor (_07925_, _07924_, _07008_);
  and (_07926_, _07925_, _07923_);
  and (_07927_, _07008_, _07178_);
  or (_07928_, _07927_, _06979_);
  or (_07929_, _07928_, _07926_);
  and (_07930_, _07929_, _07908_);
  or (_07931_, _07930_, _01953_);
  nand (_07932_, _04759_, _01953_);
  and (_07933_, _07932_, _07546_);
  and (_07934_, _07933_, _07931_);
  or (_07935_, _07906_, _05203_);
  and (_07936_, _07920_, _07935_);
  and (_07937_, _07936_, _07023_);
  or (_07938_, _07937_, _07934_);
  and (_07939_, _07938_, _01632_);
  or (_07940_, _01632_, \oc8051_golden_model_1.PC [1]);
  nand (_07941_, _01942_, _07940_);
  or (_07942_, _07941_, _07939_);
  and (_07943_, _07942_, _07896_);
  or (_07944_, _07943_, _03273_);
  and (_07945_, _03613_, _01853_);
  nand (_07946_, _04758_, _03273_);
  or (_07947_, _07946_, _07945_);
  and (_07948_, _07947_, _07944_);
  or (_07949_, _07948_, _02217_);
  nor (_07950_, _05226_, _04110_);
  and (_07951_, _04109_, \oc8051_golden_model_1.PSW [7]);
  and (_07952_, _07951_, _02263_);
  nor (_07953_, _07952_, _07950_);
  nand (_07954_, _07953_, _02217_);
  and (_07955_, _07954_, _07270_);
  and (_07956_, _07955_, _07949_);
  and (_07957_, _01606_, _01298_);
  or (_07958_, _07039_, _07957_);
  or (_07959_, _07958_, _07956_);
  and (_07960_, _07959_, _07895_);
  or (_07961_, _07960_, _07037_);
  or (_07962_, _07571_, _03613_);
  and (_07963_, _07962_, _07106_);
  and (_07964_, _07963_, _07961_);
  nor (_07965_, _03393_, _02962_);
  and (_07966_, _05544_, \oc8051_golden_model_1.PSW [1]);
  and (_07967_, _05553_, \oc8051_golden_model_1.B [1]);
  nor (_07968_, _07967_, _07966_);
  and (_07969_, _05540_, \oc8051_golden_model_1.TCON [1]);
  and (_07970_, _05550_, \oc8051_golden_model_1.ACC [1]);
  nor (_07971_, _07970_, _07969_);
  and (_07972_, _07971_, _07968_);
  and (_07973_, _05556_, \oc8051_golden_model_1.P0INREG [1]);
  and (_07974_, _05527_, \oc8051_golden_model_1.P1INREG [1]);
  nor (_07975_, _07974_, _07973_);
  and (_07976_, _05558_, \oc8051_golden_model_1.SCON [1]);
  and (_07977_, _05534_, \oc8051_golden_model_1.SBUF [1]);
  nor (_07978_, _07977_, _07976_);
  and (_07979_, _07978_, _07975_);
  and (_07980_, _07979_, _07972_);
  and (_07981_, _05567_, \oc8051_golden_model_1.PCON [1]);
  and (_07982_, _05569_, \oc8051_golden_model_1.DPH [1]);
  nor (_07983_, _07982_, _07981_);
  and (_07984_, _07983_, _07980_);
  and (_07985_, _05582_, \oc8051_golden_model_1.TL0 [1]);
  and (_07986_, _05587_, \oc8051_golden_model_1.TH0 [1]);
  nor (_07987_, _07986_, _07985_);
  and (_07988_, _05576_, \oc8051_golden_model_1.DPL [1]);
  and (_07989_, _05629_, \oc8051_golden_model_1.TMOD [1]);
  nor (_07990_, _07989_, _07988_);
  and (_07991_, _07990_, _07987_);
  and (_07992_, _05595_, \oc8051_golden_model_1.TH1 [1]);
  and (_07993_, _05578_, \oc8051_golden_model_1.TL1 [1]);
  nor (_07994_, _07993_, _07992_);
  and (_07995_, _05633_, \oc8051_golden_model_1.SP [1]);
  not (_07996_, _07995_);
  and (_07997_, _05615_, \oc8051_golden_model_1.P2INREG [1]);
  and (_07998_, _05609_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_07999_, _07998_, _07997_);
  and (_08000_, _05603_, \oc8051_golden_model_1.IE [1]);
  and (_08001_, _05619_, \oc8051_golden_model_1.IP [1]);
  nor (_08002_, _08001_, _08000_);
  and (_08003_, _08002_, _07999_);
  and (_08004_, _08003_, _07996_);
  and (_08005_, _08004_, _07994_);
  and (_08006_, _08005_, _07991_);
  and (_08007_, _08006_, _07984_);
  not (_08008_, _08007_);
  nor (_08009_, _08008_, _07965_);
  nor (_08010_, _08009_, _07042_);
  or (_08011_, _08010_, _02859_);
  or (_08012_, _08011_, _07964_);
  and (_08013_, _02859_, _02643_);
  nor (_08014_, _08013_, _06976_);
  and (_08015_, _08014_, _08012_);
  and (_08016_, _06976_, _05573_);
  or (_08017_, _08016_, _01650_);
  or (_08018_, _08017_, _08015_);
  and (_08019_, _01650_, \oc8051_golden_model_1.PC [1]);
  nor (_08020_, _08019_, _07061_);
  and (_08021_, _08020_, _08018_);
  and (_08022_, _04452_, _02676_);
  nor (_08023_, _08022_, _07893_);
  nor (_08024_, _08023_, _07062_);
  nor (_08025_, _08024_, _07063_);
  or (_08026_, _08025_, _08021_);
  nor (_08027_, _04452_, _01705_);
  and (_08028_, _04452_, _01705_);
  nor (_08029_, _08028_, _08027_);
  or (_08030_, _08029_, _07584_);
  and (_08031_, _08030_, _07060_);
  and (_08032_, _08031_, _08026_);
  or (_08033_, _08032_, _07894_);
  and (_08034_, _08033_, _07058_);
  and (_08035_, _08027_, _07057_);
  or (_08036_, _08035_, _01666_);
  or (_08037_, _08036_, _08034_);
  and (_08038_, _01666_, \oc8051_golden_model_1.PC [1]);
  nor (_08039_, _08038_, _07598_);
  and (_08040_, _08039_, _08037_);
  nand (_08041_, _08022_, _07603_);
  and (_08042_, _08041_, _07107_);
  or (_08043_, _08042_, _08040_);
  nand (_08044_, _08028_, _07602_);
  and (_08045_, _08044_, _05157_);
  and (_08046_, _08045_, _08043_);
  nand (_08047_, _01660_, _01298_);
  nand (_08048_, _02347_, _04918_);
  nand (_08049_, _08048_, _08047_);
  or (_08050_, _07116_, _02348_);
  or (_08051_, _08050_, _08049_);
  or (_08052_, _08051_, _08046_);
  nand (_08053_, _08052_, _07892_);
  nand (_08054_, _08053_, _07120_);
  not (_08055_, _07120_);
  nand (_08056_, _07891_, _08055_);
  and (_08057_, _08056_, _07623_);
  and (_08058_, _08057_, _08054_);
  or (_08059_, _08058_, _07889_);
  and (_08060_, _08059_, _07622_);
  nor (_08061_, _07909_, _07622_);
  or (_08062_, _08061_, _02023_);
  or (_08063_, _08062_, _08060_);
  nand (_08064_, _02023_, _03115_);
  and (_08065_, _08064_, _01671_);
  and (_08066_, _08065_, _08063_);
  and (_08067_, _01670_, _01298_);
  or (_08068_, _06973_, _08067_);
  or (_08069_, _08068_, _08066_);
  or (_08070_, _07950_, _06974_);
  and (_08071_, _08070_, _05444_);
  and (_08072_, _08071_, _08069_);
  and (_08073_, _07891_, _07651_);
  or (_08074_, _08073_, _05441_);
  or (_08075_, _08074_, _08072_);
  and (_08076_, _08075_, _07888_);
  or (_08077_, _08076_, _07095_);
  not (_08078_, _07095_);
  or (_08079_, _07909_, _08078_);
  and (_08080_, _08079_, _07169_);
  and (_08081_, _08080_, _08077_);
  or (_08082_, _08081_, _07693_);
  and (_08083_, _08082_, _07886_);
  nor (_08084_, _04616_, _02023_);
  and (_08085_, _02983_, _02023_);
  or (_08086_, _08085_, _08084_);
  and (_08087_, _08086_, _07683_);
  or (_29637_, _08087_, _08083_);
  or (_08088_, _07690_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_08089_, _08088_, _07684_);
  nor (_08090_, _07497_, _07388_);
  nor (_08091_, _08090_, _07498_);
  and (_08092_, _08091_, _07651_);
  and (_08093_, _05494_, _04252_);
  nor (_08094_, _05494_, _04252_);
  nor (_08095_, _08094_, _08093_);
  nand (_08096_, _08095_, _07080_);
  nor (_08097_, _04252_, _02309_);
  and (_08098_, _08097_, _07059_);
  and (_08099_, _04099_, \oc8051_golden_model_1.P0 [2]);
  and (_08100_, _05189_, \oc8051_golden_model_1.P2 [2]);
  nor (_08101_, _08100_, _08099_);
  and (_08102_, _05195_, \oc8051_golden_model_1.P1 [2]);
  and (_08103_, _05191_, \oc8051_golden_model_1.P3 [2]);
  nor (_08104_, _08103_, _08102_);
  and (_08105_, _08104_, _08101_);
  and (_08106_, _08105_, _05188_);
  and (_08107_, _08106_, _05183_);
  and (_08108_, _08107_, _04205_);
  nor (_08109_, _08108_, _04106_);
  or (_08110_, _08109_, _06980_);
  nand (_08111_, _08108_, _05162_);
  or (_08112_, _08111_, _07513_);
  nor (_08113_, _08095_, _06987_);
  and (_08114_, _07517_, _03272_);
  nor (_08115_, _07517_, _03272_);
  or (_08116_, _08115_, _08114_);
  or (_08117_, _08116_, _04709_);
  nor (_08118_, _01792_, _01625_);
  and (_08119_, _01625_, \oc8051_golden_model_1.ACC [2]);
  or (_08120_, _08119_, _08118_);
  nor (_08121_, _08120_, _04557_);
  nor (_08122_, _08121_, _06986_);
  and (_08123_, _08122_, _08117_);
  or (_08124_, _08123_, _06982_);
  or (_08125_, _08124_, _08113_);
  and (_08126_, _08125_, _08112_);
  or (_08127_, _08126_, _06363_);
  nor (_08128_, _01770_, _01621_);
  nor (_08129_, _08128_, _07008_);
  and (_08130_, _08129_, _08127_);
  and (_08131_, _07008_, _07388_);
  or (_08132_, _08131_, _06979_);
  or (_08133_, _08132_, _08130_);
  and (_08134_, _08133_, _08110_);
  or (_08135_, _08134_, _01953_);
  nand (_08136_, _04793_, _01953_);
  and (_08137_, _08136_, _07546_);
  and (_08138_, _08137_, _08135_);
  or (_08139_, _08108_, _05162_);
  and (_08140_, _08111_, _08139_);
  and (_08141_, _08140_, _07023_);
  or (_08142_, _08141_, _08138_);
  and (_08143_, _08142_, _01632_);
  or (_08144_, _01792_, _01632_);
  nand (_08145_, _01942_, _08144_);
  or (_08146_, _08145_, _08143_);
  nand (_08147_, _04793_, _01950_);
  and (_08148_, _08147_, _08146_);
  or (_08149_, _08148_, _03273_);
  and (_08150_, _03564_, _01853_);
  nand (_08151_, _04792_, _03273_);
  or (_08152_, _08151_, _08150_);
  and (_08153_, _08152_, _08149_);
  or (_08154_, _08153_, _02217_);
  nor (_08155_, _05201_, _04106_);
  and (_08156_, _04105_, \oc8051_golden_model_1.PSW [7]);
  and (_08157_, _08156_, _02263_);
  nor (_08158_, _08157_, _08155_);
  nand (_08159_, _08158_, _02217_);
  and (_08160_, _08159_, _07270_);
  and (_08161_, _08160_, _08154_);
  and (_08162_, _01770_, _01606_);
  or (_08163_, _07039_, _08162_);
  or (_08164_, _08163_, _08161_);
  nand (_08165_, _07039_, _03272_);
  and (_08166_, _08165_, _08164_);
  or (_08167_, _08166_, _07037_);
  or (_08168_, _07571_, _03564_);
  and (_08169_, _08168_, _07106_);
  and (_08170_, _08169_, _08167_);
  nor (_08171_, _03272_, _02962_);
  and (_08172_, _05540_, \oc8051_golden_model_1.TCON [2]);
  and (_08173_, _05550_, \oc8051_golden_model_1.ACC [2]);
  nor (_08174_, _08173_, _08172_);
  and (_08175_, _05556_, \oc8051_golden_model_1.P0INREG [2]);
  and (_08176_, _05558_, \oc8051_golden_model_1.SCON [2]);
  nor (_08177_, _08176_, _08175_);
  and (_08178_, _08177_, _08174_);
  and (_08179_, _05534_, \oc8051_golden_model_1.SBUF [2]);
  and (_08180_, _05553_, \oc8051_golden_model_1.B [2]);
  nor (_08181_, _08180_, _08179_);
  and (_08182_, _05527_, \oc8051_golden_model_1.P1INREG [2]);
  and (_08183_, _05544_, \oc8051_golden_model_1.PSW [2]);
  nor (_08184_, _08183_, _08182_);
  and (_08185_, _08184_, _08181_);
  and (_08186_, _08185_, _08178_);
  and (_08187_, _05567_, \oc8051_golden_model_1.PCON [2]);
  and (_08188_, _05569_, \oc8051_golden_model_1.DPH [2]);
  nor (_08189_, _08188_, _08187_);
  and (_08190_, _08189_, _08186_);
  and (_08191_, _05576_, \oc8051_golden_model_1.DPL [2]);
  and (_08193_, _05578_, \oc8051_golden_model_1.TL1 [2]);
  nor (_08194_, _08193_, _08191_);
  and (_08195_, _05633_, \oc8051_golden_model_1.SP [2]);
  and (_08196_, _05587_, \oc8051_golden_model_1.TH0 [2]);
  nor (_08197_, _08196_, _08195_);
  and (_08198_, _08197_, _08194_);
  and (_08199_, _05582_, \oc8051_golden_model_1.TL0 [2]);
  not (_08200_, _08199_);
  and (_08201_, _05603_, \oc8051_golden_model_1.IE [2]);
  and (_08202_, _05609_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_08203_, _08202_, _08201_);
  and (_08204_, _05615_, \oc8051_golden_model_1.P2INREG [2]);
  and (_08205_, _05619_, \oc8051_golden_model_1.IP [2]);
  nor (_08206_, _08205_, _08204_);
  and (_08207_, _08206_, _08203_);
  and (_08208_, _08207_, _08200_);
  and (_08209_, _05595_, \oc8051_golden_model_1.TH1 [2]);
  and (_08210_, _05629_, \oc8051_golden_model_1.TMOD [2]);
  nor (_08211_, _08210_, _08209_);
  and (_08212_, _08211_, _08208_);
  and (_08213_, _08212_, _08198_);
  and (_08214_, _08213_, _08190_);
  not (_08215_, _08214_);
  nor (_08216_, _08215_, _08171_);
  nor (_08217_, _08216_, _07042_);
  or (_08218_, _08217_, _02859_);
  or (_08219_, _08218_, _08170_);
  and (_08220_, _02859_, _02263_);
  nor (_08221_, _08220_, _06976_);
  and (_08222_, _08221_, _08219_);
  and (_08223_, _06976_, _05563_);
  or (_08224_, _08223_, _01650_);
  or (_08225_, _08224_, _08222_);
  and (_08226_, _01792_, _01650_);
  nor (_08227_, _08226_, _07061_);
  and (_08228_, _08227_, _08225_);
  and (_08229_, _04252_, _02309_);
  nor (_08230_, _08229_, _08097_);
  nor (_08231_, _08230_, _07062_);
  nor (_08232_, _08231_, _07063_);
  or (_08233_, _08232_, _08228_);
  not (_08234_, \oc8051_golden_model_1.ACC [2]);
  nor (_08235_, _04252_, _08234_);
  and (_08236_, _04252_, _08234_);
  nor (_08237_, _08236_, _08235_);
  or (_08238_, _08237_, _07584_);
  and (_08239_, _08238_, _07060_);
  and (_08240_, _08239_, _08233_);
  or (_08241_, _08240_, _08098_);
  and (_08242_, _08241_, _07058_);
  and (_08243_, _08235_, _07057_);
  or (_08244_, _08243_, _01666_);
  or (_08245_, _08244_, _08242_);
  and (_08246_, _01792_, _01666_);
  nor (_08247_, _08246_, _07598_);
  and (_08248_, _08247_, _08245_);
  nand (_08249_, _08229_, _07603_);
  and (_08250_, _08249_, _07107_);
  or (_08251_, _08250_, _08248_);
  nand (_08252_, _08236_, _07602_);
  and (_08253_, _08252_, _05157_);
  and (_08254_, _08253_, _08251_);
  and (_08255_, _01770_, _01660_);
  or (_08256_, _05416_, _08255_);
  or (_08257_, _08256_, _08254_);
  or (_08258_, _08116_, _05415_);
  and (_08259_, _08258_, _07623_);
  and (_08260_, _08259_, _08257_);
  nor (_08261_, _07630_, _07629_);
  or (_08262_, _08261_, _07631_);
  and (_08263_, _08262_, _05417_);
  or (_08264_, _08263_, _07080_);
  or (_08265_, _08264_, _08260_);
  and (_08266_, _08265_, _08096_);
  or (_08267_, _08266_, _02023_);
  nand (_08268_, _03113_, _02023_);
  and (_08269_, _08268_, _01671_);
  and (_08270_, _08269_, _08267_);
  and (_08271_, _01770_, _01670_);
  or (_08272_, _06973_, _08271_);
  or (_08273_, _08272_, _08270_);
  or (_08274_, _08155_, _06974_);
  and (_08275_, _08274_, _05444_);
  and (_08276_, _08275_, _08273_);
  or (_08277_, _08276_, _08092_);
  and (_08278_, _08277_, _05442_);
  or (_08279_, _07658_, _03564_);
  nor (_08280_, _07659_, _05442_);
  and (_08281_, _08280_, _08279_);
  or (_08282_, _08281_, _07095_);
  or (_08283_, _08282_, _08278_);
  nor (_08284_, _05743_, _05739_);
  nor (_08285_, _08284_, _05745_);
  or (_08286_, _08285_, _08078_);
  and (_08287_, _08286_, _07169_);
  and (_08288_, _08287_, _08283_);
  or (_08289_, _08288_, _07693_);
  and (_08291_, _08289_, _08089_);
  and (_08292_, _02967_, _02023_);
  nor (_08294_, _04601_, _02023_);
  or (_08295_, _08294_, _08292_);
  and (_08297_, _08295_, _07683_);
  or (_29638_, _08297_, _08291_);
  or (_08299_, _07690_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_08300_, _08299_, _07684_);
  and (_08301_, _01720_, _01660_);
  nor (_08302_, _04204_, _01732_);
  and (_08303_, _04204_, _01732_);
  nor (_08304_, _08303_, _08302_);
  and (_08305_, _08304_, _07062_);
  nor (_08306_, _05357_, _04101_);
  and (_08307_, _06260_, _02263_);
  nor (_08308_, _08307_, _08306_);
  nor (_08309_, _08308_, _07271_);
  nand (_08310_, _03516_, _01853_);
  nand (_08311_, _08310_, _04854_);
  and (_08312_, _08311_, _03273_);
  and (_08313_, _05195_, \oc8051_golden_model_1.P1 [3]);
  and (_08314_, _05191_, \oc8051_golden_model_1.P3 [3]);
  nor (_08315_, _08314_, _08313_);
  and (_08316_, _05189_, \oc8051_golden_model_1.P2 [3]);
  and (_08317_, _04099_, \oc8051_golden_model_1.P0 [3]);
  nor (_08318_, _08317_, _08316_);
  and (_08319_, _08318_, _08315_);
  and (_08320_, _08319_, _05341_);
  and (_08321_, _08320_, _05350_);
  and (_08322_, _08321_, _05343_);
  and (_08323_, _08322_, _04095_);
  nor (_08324_, _08323_, _04101_);
  or (_08325_, _08324_, _06980_);
  nor (_08326_, _08114_, _03473_);
  or (_08327_, _08326_, _07518_);
  or (_08328_, _08327_, _04709_);
  and (_08329_, _01625_, \oc8051_golden_model_1.ACC [3]);
  nor (_08330_, _02060_, _01625_);
  or (_08331_, _04557_, _08330_);
  or (_08332_, _08331_, _08329_);
  and (_08333_, _08332_, _08328_);
  and (_08334_, _08333_, _06987_);
  and (_08335_, _05494_, _04253_);
  nor (_08336_, _08093_, _04204_);
  nor (_08337_, _08336_, _08335_);
  nor (_08338_, _08337_, _06987_);
  or (_08339_, _08338_, _08334_);
  or (_08340_, _08339_, _06982_);
  nand (_08341_, _08323_, _05334_);
  or (_08342_, _08341_, _07513_);
  and (_08343_, _08342_, _08340_);
  or (_08344_, _08343_, _06363_);
  nor (_08345_, _01720_, _01621_);
  nor (_08346_, _08345_, _07008_);
  and (_08347_, _08346_, _08344_);
  and (_08348_, _07008_, _07496_);
  or (_08349_, _08348_, _06979_);
  or (_08350_, _08349_, _08347_);
  and (_08351_, _08350_, _08325_);
  or (_08352_, _08351_, _01953_);
  nand (_08353_, _04855_, _01953_);
  and (_08354_, _08353_, _07546_);
  and (_08355_, _08354_, _08352_);
  nor (_08356_, _08323_, _05334_);
  not (_08357_, _08356_);
  and (_08358_, _08341_, _08357_);
  and (_08359_, _08358_, _07023_);
  or (_08360_, _08359_, _08355_);
  and (_08361_, _08360_, _01632_);
  or (_08362_, _02060_, _01632_);
  nand (_08363_, _01942_, _08362_);
  or (_08364_, _08363_, _08361_);
  nand (_08365_, _04855_, _01950_);
  and (_08366_, _08365_, _03274_);
  and (_08367_, _08366_, _08364_);
  or (_08368_, _08367_, _08312_);
  and (_08369_, _08368_, _07271_);
  or (_08370_, _08369_, _08309_);
  and (_08371_, _08370_, _07270_);
  and (_08372_, _01720_, _01606_);
  or (_08373_, _07039_, _08372_);
  or (_08374_, _08373_, _08371_);
  nand (_08375_, _07039_, _03473_);
  and (_08376_, _08375_, _08374_);
  or (_08377_, _08376_, _07037_);
  or (_08378_, _07571_, _03516_);
  and (_08379_, _08378_, _07106_);
  and (_08380_, _08379_, _08377_);
  nor (_08381_, _03473_, _02962_);
  and (_08382_, _05540_, \oc8051_golden_model_1.TCON [3]);
  and (_08383_, _05550_, \oc8051_golden_model_1.ACC [3]);
  nor (_08384_, _08383_, _08382_);
  and (_08385_, _05556_, \oc8051_golden_model_1.P0INREG [3]);
  and (_08386_, _05527_, \oc8051_golden_model_1.P1INREG [3]);
  nor (_08387_, _08386_, _08385_);
  and (_08388_, _08387_, _08384_);
  and (_08389_, _05544_, \oc8051_golden_model_1.PSW [3]);
  and (_08390_, _05553_, \oc8051_golden_model_1.B [3]);
  nor (_08391_, _08390_, _08389_);
  and (_08392_, _05558_, \oc8051_golden_model_1.SCON [3]);
  and (_08393_, _05534_, \oc8051_golden_model_1.SBUF [3]);
  nor (_08394_, _08393_, _08392_);
  and (_08395_, _08394_, _08391_);
  and (_08396_, _08395_, _08388_);
  and (_08397_, _05567_, \oc8051_golden_model_1.PCON [3]);
  and (_08398_, _05569_, \oc8051_golden_model_1.DPH [3]);
  nor (_08399_, _08398_, _08397_);
  and (_08400_, _08399_, _08396_);
  and (_08401_, _05576_, \oc8051_golden_model_1.DPL [3]);
  and (_08402_, _05629_, \oc8051_golden_model_1.TMOD [3]);
  nor (_08403_, _08402_, _08401_);
  and (_08404_, _05582_, \oc8051_golden_model_1.TL0 [3]);
  and (_08405_, _05595_, \oc8051_golden_model_1.TH1 [3]);
  nor (_08406_, _08405_, _08404_);
  and (_08407_, _08406_, _08403_);
  and (_08408_, _05578_, \oc8051_golden_model_1.TL1 [3]);
  not (_08409_, _08408_);
  and (_08410_, _05615_, \oc8051_golden_model_1.P2INREG [3]);
  and (_08411_, _05609_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_08412_, _08411_, _08410_);
  and (_08413_, _05603_, \oc8051_golden_model_1.IE [3]);
  and (_08414_, _05619_, \oc8051_golden_model_1.IP [3]);
  nor (_08415_, _08414_, _08413_);
  and (_08416_, _08415_, _08412_);
  and (_08417_, _08416_, _08409_);
  and (_08418_, _05633_, \oc8051_golden_model_1.SP [3]);
  and (_08419_, _05587_, \oc8051_golden_model_1.TH0 [3]);
  nor (_08420_, _08419_, _08418_);
  and (_08421_, _08420_, _08417_);
  and (_08422_, _08421_, _08407_);
  and (_08423_, _08422_, _08400_);
  not (_08424_, _08423_);
  nor (_08425_, _08424_, _08381_);
  nor (_08426_, _08425_, _07042_);
  or (_08427_, _08426_, _02859_);
  or (_08428_, _08427_, _08380_);
  not (_08429_, _02859_);
  nor (_08430_, _08429_, _01916_);
  nor (_08431_, _08430_, _06976_);
  and (_08432_, _08431_, _08428_);
  and (_08433_, _06976_, _05529_);
  or (_08434_, _08433_, _01650_);
  or (_08435_, _08434_, _08432_);
  and (_08436_, _02060_, _01650_);
  nor (_08437_, _08436_, _07061_);
  and (_08438_, _08437_, _08435_);
  nor (_08439_, _04204_, _02119_);
  and (_08440_, _04204_, _02119_);
  nor (_08441_, _08440_, _08439_);
  and (_08442_, _08441_, _07061_);
  or (_08443_, _08442_, _08438_);
  and (_08444_, _08443_, _07584_);
  or (_08445_, _08444_, _08305_);
  and (_08446_, _08445_, _07060_);
  and (_08447_, _08439_, _07059_);
  or (_08448_, _08447_, _08446_);
  and (_08449_, _08448_, _07058_);
  and (_08450_, _08302_, _07057_);
  or (_08452_, _08450_, _01666_);
  or (_08454_, _08452_, _08449_);
  and (_08456_, _02060_, _01666_);
  nor (_08458_, _08456_, _07598_);
  and (_08460_, _08458_, _08454_);
  nand (_08462_, _08440_, _07603_);
  and (_08464_, _08462_, _07107_);
  or (_08466_, _08464_, _08460_);
  nand (_08468_, _08303_, _07602_);
  and (_08469_, _08468_, _05157_);
  and (_08470_, _08469_, _08466_);
  or (_08471_, _08470_, _08301_);
  and (_08472_, _08471_, _07610_);
  or (_08473_, _08327_, _07614_);
  and (_08474_, _08473_, _05416_);
  or (_08475_, _08474_, _08472_);
  or (_08476_, _08327_, _07615_);
  and (_08477_, _08476_, _07623_);
  and (_08478_, _08477_, _08475_);
  nor (_08479_, _07631_, _07628_);
  or (_08480_, _08479_, _07632_);
  and (_08481_, _08480_, _05417_);
  or (_08482_, _08481_, _08478_);
  and (_08483_, _08482_, _07622_);
  nor (_08484_, _08337_, _07622_);
  or (_08485_, _08484_, _02023_);
  or (_08486_, _08485_, _08483_);
  nand (_08487_, _03108_, _02023_);
  and (_08488_, _08487_, _01671_);
  and (_08489_, _08488_, _08486_);
  and (_08490_, _01720_, _01670_);
  or (_08491_, _06973_, _08490_);
  or (_08492_, _08491_, _08489_);
  or (_08493_, _08306_, _06974_);
  and (_08494_, _08493_, _05444_);
  and (_08495_, _08494_, _08492_);
  nor (_08496_, _07498_, _07496_);
  nor (_08497_, _08496_, _07499_);
  and (_08498_, _08497_, _07651_);
  or (_08499_, _08498_, _05441_);
  or (_08500_, _08499_, _08495_);
  nor (_08501_, _07659_, _03516_);
  nor (_08502_, _08501_, _07660_);
  or (_08503_, _08502_, _05442_);
  and (_08504_, _08503_, _08078_);
  and (_08505_, _08504_, _08500_);
  nor (_08506_, _05745_, _05737_);
  nor (_08507_, _08506_, _05747_);
  and (_08508_, _08507_, _07095_);
  nor (_08509_, _08508_, _08505_);
  nor (_08510_, _08509_, _07170_);
  or (_08511_, _08510_, _07693_);
  and (_08512_, _08511_, _08300_);
  and (_08513_, _02974_, _02023_);
  nor (_08514_, _04607_, _02023_);
  or (_08515_, _08514_, _08513_);
  and (_08516_, _08515_, _07683_);
  or (_29639_, _08516_, _08512_);
  and (_08517_, _02010_, _01589_);
  nor (_08518_, _07499_, _07495_);
  nor (_08519_, _08518_, _07500_);
  and (_08520_, _08519_, _08517_);
  nor (_08521_, _07632_, _07627_);
  or (_08522_, _08521_, _07633_);
  and (_08523_, _08522_, _05417_);
  not (_08524_, \oc8051_golden_model_1.ACC [4]);
  nor (_08525_, _04299_, _08524_);
  and (_08526_, _04299_, _08524_);
  nor (_08527_, _08526_, _08525_);
  and (_08528_, _08527_, _07062_);
  nor (_08529_, _04299_, _03101_);
  and (_08530_, _04299_, _03101_);
  nor (_08531_, _08530_, _08529_);
  and (_08532_, _08531_, _07061_);
  and (_08533_, _04641_, _01606_);
  and (_08534_, _04099_, \oc8051_golden_model_1.P0 [4]);
  and (_08535_, _05191_, \oc8051_golden_model_1.P3 [4]);
  nor (_08536_, _08535_, _08534_);
  and (_08537_, _05195_, \oc8051_golden_model_1.P1 [4]);
  and (_08538_, _05189_, \oc8051_golden_model_1.P2 [4]);
  nor (_08539_, _08538_, _08537_);
  and (_08540_, _08539_, _08536_);
  and (_08541_, _08540_, _05241_);
  and (_08542_, _08541_, _05238_);
  and (_08543_, _08542_, _04254_);
  nor (_08544_, _08543_, _05252_);
  or (_08545_, _08544_, _06980_);
  nor (_08546_, _08335_, _04299_);
  and (_08547_, _08335_, _04299_);
  nor (_08548_, _08547_, _08546_);
  nor (_08549_, _08548_, _06987_);
  or (_08550_, _07515_, _03903_);
  nor (_08551_, _07518_, _04024_);
  and (_08552_, _07518_, _04024_);
  or (_08553_, _08552_, _08551_);
  and (_08554_, _08553_, _04557_);
  nor (_08555_, _04642_, _01625_);
  and (_08556_, _01625_, \oc8051_golden_model_1.ACC [4]);
  or (_08557_, _08556_, _08555_);
  and (_08558_, _08557_, _04709_);
  or (_08559_, _08558_, _04715_);
  or (_08560_, _08559_, _08554_);
  and (_08561_, _08560_, _06987_);
  and (_08562_, _08561_, _08550_);
  or (_08563_, _08562_, _08549_);
  and (_08564_, _08563_, _07513_);
  nand (_08565_, _08543_, _05253_);
  and (_08566_, _08565_, _06982_);
  or (_08567_, _08566_, _06363_);
  or (_08568_, _08567_, _08564_);
  nor (_08569_, _04641_, _01621_);
  nor (_08570_, _08569_, _07008_);
  and (_08571_, _08570_, _08568_);
  and (_08572_, _07008_, _07495_);
  or (_08573_, _08572_, _06979_);
  or (_08574_, _08573_, _08571_);
  and (_08575_, _08574_, _08545_);
  or (_08576_, _08575_, _01953_);
  nand (_08577_, _04841_, _01953_);
  and (_08578_, _08577_, _07546_);
  and (_08579_, _08578_, _08576_);
  nor (_08580_, _08543_, _05253_);
  not (_08581_, _08580_);
  and (_08582_, _08565_, _08581_);
  and (_08583_, _08582_, _07023_);
  or (_08584_, _08583_, _08579_);
  and (_08585_, _08584_, _01632_);
  nor (_08586_, _04642_, _01632_);
  not (_08587_, _02030_);
  nand (_08588_, _07128_, _08587_);
  and (_08589_, _08588_, _01929_);
  or (_08590_, _08589_, _08586_);
  or (_08591_, _08590_, _08585_);
  and (_08592_, _02010_, _01929_);
  and (_08593_, _08589_, _04841_);
  nor (_08594_, _08593_, _08592_);
  and (_08595_, _08594_, _08591_);
  not (_08596_, _08592_);
  nor (_08597_, _04841_, _08596_);
  or (_08598_, _08597_, _03273_);
  or (_08599_, _08598_, _08595_);
  and (_08600_, _03903_, _01853_);
  nand (_08601_, _04840_, _03273_);
  or (_08602_, _08601_, _08600_);
  and (_08603_, _08602_, _08599_);
  or (_08604_, _08603_, _02217_);
  nor (_08605_, _05252_, _05251_);
  and (_08606_, _07757_, _02264_);
  nor (_08607_, _08606_, _08605_);
  nand (_08608_, _08607_, _02217_);
  and (_08609_, _08608_, _07270_);
  and (_08610_, _08609_, _08604_);
  or (_08611_, _08610_, _08533_);
  and (_08612_, _08611_, _07700_);
  nor (_08613_, _07700_, _04024_);
  or (_08614_, _08613_, _07037_);
  or (_08615_, _08614_, _08612_);
  or (_08616_, _07571_, _03903_);
  and (_08617_, _08616_, _07042_);
  and (_08618_, _08617_, _08615_);
  nor (_08619_, _04024_, _02962_);
  and (_08620_, _05556_, \oc8051_golden_model_1.P0INREG [4]);
  and (_08621_, _05534_, \oc8051_golden_model_1.SBUF [4]);
  nor (_08622_, _08621_, _08620_);
  and (_08623_, _05553_, \oc8051_golden_model_1.B [4]);
  and (_08624_, _05544_, \oc8051_golden_model_1.PSW [4]);
  nor (_08625_, _08624_, _08623_);
  and (_08626_, _08625_, _08622_);
  and (_08627_, _05540_, \oc8051_golden_model_1.TCON [4]);
  and (_08628_, _05527_, \oc8051_golden_model_1.P1INREG [4]);
  nor (_08629_, _08628_, _08627_);
  and (_08630_, _05558_, \oc8051_golden_model_1.SCON [4]);
  and (_08631_, _05550_, \oc8051_golden_model_1.ACC [4]);
  nor (_08632_, _08631_, _08630_);
  and (_08633_, _08632_, _08629_);
  and (_08634_, _08633_, _08626_);
  and (_08635_, _05567_, \oc8051_golden_model_1.PCON [4]);
  and (_08636_, _05569_, \oc8051_golden_model_1.DPH [4]);
  nor (_08637_, _08636_, _08635_);
  and (_08638_, _08637_, _08634_);
  and (_08639_, _05576_, \oc8051_golden_model_1.DPL [4]);
  and (_08640_, _05633_, \oc8051_golden_model_1.SP [4]);
  nor (_08641_, _08640_, _08639_);
  and (_08642_, _05582_, \oc8051_golden_model_1.TL0 [4]);
  and (_08643_, _05595_, \oc8051_golden_model_1.TH1 [4]);
  nor (_08644_, _08643_, _08642_);
  and (_08645_, _08644_, _08641_);
  and (_08646_, _05587_, \oc8051_golden_model_1.TH0 [4]);
  not (_08647_, _08646_);
  and (_08648_, _05615_, \oc8051_golden_model_1.P2INREG [4]);
  and (_08649_, _05603_, \oc8051_golden_model_1.IE [4]);
  nor (_08650_, _08649_, _08648_);
  and (_08651_, _05609_, \oc8051_golden_model_1.P3INREG [4]);
  and (_08652_, _05619_, \oc8051_golden_model_1.IP [4]);
  nor (_08653_, _08652_, _08651_);
  and (_08654_, _08653_, _08650_);
  and (_08655_, _08654_, _08647_);
  and (_08656_, _05629_, \oc8051_golden_model_1.TMOD [4]);
  and (_08657_, _05578_, \oc8051_golden_model_1.TL1 [4]);
  nor (_08658_, _08657_, _08656_);
  and (_08659_, _08658_, _08655_);
  and (_08660_, _08659_, _08645_);
  and (_08661_, _08660_, _08638_);
  not (_08662_, _08661_);
  nor (_08663_, _08662_, _08619_);
  nor (_08664_, _08663_, _07042_);
  or (_08665_, _08664_, _02859_);
  or (_08666_, _08665_, _08618_);
  and (_08667_, _02859_, _02606_);
  nor (_08668_, _08667_, _06976_);
  and (_08669_, _08668_, _08666_);
  and (_08670_, _06976_, _05524_);
  or (_08671_, _08670_, _01650_);
  or (_08672_, _08671_, _08669_);
  and (_08673_, _04642_, _01650_);
  nor (_08674_, _08673_, _07061_);
  and (_08675_, _08674_, _08672_);
  or (_08676_, _08675_, _08532_);
  and (_08677_, _08676_, _07584_);
  or (_08678_, _08677_, _08528_);
  and (_08679_, _08678_, _07060_);
  and (_08680_, _08529_, _07059_);
  or (_08681_, _08680_, _08679_);
  and (_08682_, _08681_, _07058_);
  and (_08683_, _08525_, _07057_);
  or (_08684_, _08683_, _01666_);
  or (_08685_, _08684_, _08682_);
  and (_08686_, _04642_, _01666_);
  nor (_08687_, _08686_, _07598_);
  and (_08688_, _08687_, _08685_);
  nand (_08689_, _08530_, _07603_);
  and (_08690_, _08689_, _07107_);
  or (_08691_, _08690_, _08688_);
  nand (_08692_, _08526_, _07602_);
  and (_08693_, _08692_, _05157_);
  and (_08694_, _08693_, _08691_);
  and (_08695_, _04641_, _01660_);
  or (_08696_, _08695_, _05416_);
  or (_08697_, _08696_, _08694_);
  or (_08698_, _08553_, _05415_);
  and (_08699_, _08698_, _07623_);
  and (_08700_, _08699_, _08697_);
  or (_08701_, _08700_, _08523_);
  and (_08702_, _08701_, _07622_);
  nor (_08703_, _08548_, _07622_);
  or (_08704_, _08703_, _02023_);
  or (_08705_, _08704_, _08702_);
  nand (_08706_, _03104_, _02023_);
  and (_08707_, _08706_, _01671_);
  and (_08708_, _08707_, _08705_);
  and (_08709_, _04641_, _01670_);
  or (_08710_, _08709_, _06973_);
  or (_08711_, _08710_, _08708_);
  and (_08712_, _01938_, _04918_);
  and (_08713_, _08712_, _01589_);
  nor (_08714_, _08713_, _02359_);
  or (_08715_, _08605_, _06974_);
  and (_08716_, _08715_, _08714_);
  and (_08717_, _08716_, _08711_);
  not (_08718_, _08714_);
  and (_08719_, _08519_, _08718_);
  nor (_08720_, _08719_, _08717_);
  nor (_08721_, _08720_, _08517_);
  or (_08722_, _08721_, _08520_);
  and (_08723_, _08722_, _05442_);
  or (_08724_, _07660_, _03903_);
  nor (_08725_, _07661_, _05442_);
  and (_08726_, _08725_, _08724_);
  or (_08727_, _08726_, _07095_);
  or (_08728_, _08727_, _08723_);
  not (_08729_, _04299_);
  and (_08730_, _05747_, _08729_);
  nor (_08731_, _05747_, _08729_);
  nor (_08732_, _08731_, _08730_);
  or (_08733_, _08732_, _08078_);
  and (_08734_, _08733_, _07169_);
  and (_08735_, _08734_, _08728_);
  or (_08736_, _08735_, _07693_);
  or (_08737_, _07690_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_08738_, _08737_, _07684_);
  and (_08739_, _08738_, _08736_);
  and (_08740_, _02964_, _02023_);
  nor (_08741_, _04597_, _02023_);
  or (_08742_, _08741_, _08740_);
  and (_08743_, _08742_, _07683_);
  or (_29640_, _08743_, _08739_);
  nor (_08744_, _08552_, _03976_);
  or (_08745_, _08744_, _07519_);
  or (_08746_, _08745_, _05415_);
  not (_08747_, \oc8051_golden_model_1.ACC [5]);
  nor (_08748_, _04347_, _08747_);
  and (_08749_, _04347_, _08747_);
  nor (_08750_, _08749_, _08748_);
  and (_08751_, _08750_, _07062_);
  nor (_08752_, _05381_, _05380_);
  and (_08753_, _07951_, _02264_);
  nor (_08754_, _08753_, _08752_);
  nor (_08755_, _08754_, _07271_);
  nand (_08756_, _04868_, _01950_);
  and (_08757_, _05191_, \oc8051_golden_model_1.P3 [5]);
  nor (_08758_, _08757_, _05372_);
  and (_08759_, _08758_, _05364_);
  and (_08760_, _05195_, \oc8051_golden_model_1.P1 [5]);
  and (_08761_, _05189_, \oc8051_golden_model_1.P2 [5]);
  and (_08762_, _04099_, \oc8051_golden_model_1.P0 [5]);
  or (_08763_, _08762_, _08761_);
  nor (_08764_, _08763_, _08760_);
  and (_08765_, _08764_, _05371_);
  and (_08766_, _08765_, _08759_);
  and (_08767_, _08766_, _04300_);
  nor (_08768_, _08767_, _05381_);
  or (_08769_, _08768_, _06980_);
  nor (_08770_, _08547_, _04347_);
  nor (_08771_, _08770_, _05495_);
  nor (_08772_, _08771_, _06987_);
  or (_08773_, _07515_, _03850_);
  and (_08774_, _08745_, _04557_);
  and (_08775_, _01625_, \oc8051_golden_model_1.ACC [5]);
  nor (_08776_, _04637_, _01625_);
  or (_08777_, _08776_, _08775_);
  and (_08778_, _08777_, _04709_);
  or (_08779_, _08778_, _04715_);
  or (_08780_, _08779_, _08774_);
  and (_08781_, _08780_, _06987_);
  and (_08782_, _08781_, _08773_);
  or (_08783_, _08782_, _08772_);
  and (_08784_, _08783_, _07513_);
  nand (_08785_, _08767_, _05382_);
  and (_08786_, _08785_, _06982_);
  or (_08787_, _08786_, _06363_);
  or (_08788_, _08787_, _08784_);
  nor (_08789_, _04636_, _01621_);
  nor (_08790_, _08789_, _07008_);
  and (_08791_, _08790_, _08788_);
  and (_08792_, _07008_, _07494_);
  or (_08793_, _08792_, _06979_);
  or (_08794_, _08793_, _08791_);
  and (_08795_, _08794_, _08769_);
  or (_08796_, _08795_, _01953_);
  nand (_08797_, _04868_, _01953_);
  and (_08798_, _08797_, _07546_);
  and (_08799_, _08798_, _08796_);
  nor (_08800_, _08767_, _05382_);
  not (_08801_, _08800_);
  and (_08802_, _08785_, _08801_);
  and (_08803_, _08802_, _07023_);
  or (_08804_, _08803_, _08799_);
  and (_08805_, _08804_, _01632_);
  or (_08806_, _04637_, _01632_);
  nand (_08807_, _08806_, _01942_);
  or (_08808_, _08807_, _08805_);
  and (_08809_, _08808_, _08756_);
  or (_08810_, _08809_, _03273_);
  and (_08811_, _03850_, _01853_);
  nand (_08812_, _04867_, _03273_);
  or (_08813_, _08812_, _08811_);
  and (_08814_, _08813_, _07271_);
  and (_08815_, _08814_, _08810_);
  or (_08816_, _08815_, _08755_);
  and (_08817_, _08816_, _07270_);
  and (_08818_, _04636_, _01606_);
  or (_08819_, _08818_, _07039_);
  or (_08820_, _08819_, _08817_);
  nand (_08821_, _07039_, _03976_);
  and (_08822_, _08821_, _08820_);
  or (_08823_, _08822_, _07037_);
  or (_08824_, _07571_, _03850_);
  and (_08825_, _08824_, _07106_);
  and (_08826_, _08825_, _08823_);
  nor (_08827_, _03976_, _02962_);
  and (_08828_, _05527_, \oc8051_golden_model_1.P1INREG [5]);
  and (_08829_, _05534_, \oc8051_golden_model_1.SBUF [5]);
  nor (_08830_, _08829_, _08828_);
  and (_08831_, _05556_, \oc8051_golden_model_1.P0INREG [5]);
  and (_08832_, _05540_, \oc8051_golden_model_1.TCON [5]);
  nor (_08833_, _08832_, _08831_);
  and (_08834_, _08833_, _08830_);
  and (_08835_, _05544_, \oc8051_golden_model_1.PSW [5]);
  and (_08836_, _05553_, \oc8051_golden_model_1.B [5]);
  nor (_08837_, _08836_, _08835_);
  and (_08838_, _05558_, \oc8051_golden_model_1.SCON [5]);
  and (_08839_, _05550_, \oc8051_golden_model_1.ACC [5]);
  nor (_08840_, _08839_, _08838_);
  and (_08841_, _08840_, _08837_);
  and (_08842_, _08841_, _08834_);
  and (_08843_, _05567_, \oc8051_golden_model_1.PCON [5]);
  and (_08844_, _05569_, \oc8051_golden_model_1.DPH [5]);
  nor (_08845_, _08844_, _08843_);
  and (_08846_, _08845_, _08842_);
  and (_08847_, _05582_, \oc8051_golden_model_1.TL0 [5]);
  and (_08848_, _05629_, \oc8051_golden_model_1.TMOD [5]);
  nor (_08849_, _08848_, _08847_);
  and (_08850_, _05576_, \oc8051_golden_model_1.DPL [5]);
  and (_08852_, _05633_, \oc8051_golden_model_1.SP [5]);
  nor (_08853_, _08852_, _08850_);
  and (_08854_, _08853_, _08849_);
  and (_08855_, _05595_, \oc8051_golden_model_1.TH1 [5]);
  and (_08856_, _05578_, \oc8051_golden_model_1.TL1 [5]);
  nor (_08857_, _08856_, _08855_);
  and (_08858_, _05587_, \oc8051_golden_model_1.TH0 [5]);
  not (_08859_, _08858_);
  and (_08860_, _05615_, \oc8051_golden_model_1.P2INREG [5]);
  and (_08861_, _05603_, \oc8051_golden_model_1.IE [5]);
  nor (_08863_, _08861_, _08860_);
  and (_08864_, _05609_, \oc8051_golden_model_1.P3INREG [5]);
  and (_08865_, _05619_, \oc8051_golden_model_1.IP [5]);
  nor (_08866_, _08865_, _08864_);
  and (_08867_, _08866_, _08863_);
  and (_08868_, _08867_, _08859_);
  and (_08869_, _08868_, _08857_);
  and (_08870_, _08869_, _08854_);
  and (_08871_, _08870_, _08846_);
  not (_08872_, _08871_);
  nor (_08874_, _08872_, _08827_);
  nor (_08875_, _08874_, _07042_);
  or (_08876_, _08875_, _02859_);
  or (_08877_, _08876_, _08826_);
  and (_08878_, _02859_, _02214_);
  nor (_08879_, _08878_, _06976_);
  and (_08880_, _08879_, _08877_);
  and (_08881_, _06976_, _05548_);
  or (_08882_, _08881_, _01650_);
  or (_08883_, _08882_, _08880_);
  and (_08885_, _04637_, _01650_);
  nor (_08886_, _08885_, _07061_);
  and (_08887_, _08886_, _08883_);
  nor (_08888_, _04347_, _03064_);
  and (_08889_, _04347_, _03064_);
  nor (_08890_, _08889_, _08888_);
  and (_08891_, _08890_, _07061_);
  or (_08892_, _08891_, _08887_);
  and (_08893_, _08892_, _07584_);
  or (_08894_, _08893_, _08751_);
  and (_08896_, _08894_, _07060_);
  and (_08897_, _08888_, _07059_);
  or (_08898_, _08897_, _08896_);
  and (_08899_, _08898_, _07058_);
  and (_08900_, _08748_, _07057_);
  or (_08901_, _08900_, _01666_);
  or (_08902_, _08901_, _08899_);
  and (_08903_, _04637_, _01666_);
  nor (_08904_, _08903_, _07598_);
  and (_08905_, _08904_, _08902_);
  nand (_08907_, _08889_, _07603_);
  and (_08908_, _08907_, _07107_);
  or (_08909_, _08908_, _08905_);
  nand (_08910_, _08749_, _07602_);
  and (_08911_, _08910_, _05157_);
  and (_08912_, _08911_, _08909_);
  and (_08913_, _04636_, _01660_);
  or (_08914_, _08913_, _05416_);
  or (_08915_, _08914_, _08912_);
  and (_08916_, _08915_, _08746_);
  or (_08918_, _08916_, _05417_);
  nor (_08919_, _07633_, _07626_);
  or (_08920_, _08919_, _07634_);
  or (_08921_, _08920_, _07623_);
  and (_08922_, _08921_, _07622_);
  and (_08923_, _08922_, _08918_);
  nor (_08924_, _08771_, _07622_);
  or (_08925_, _08924_, _02023_);
  or (_08926_, _08925_, _08923_);
  nand (_08927_, _03068_, _02023_);
  and (_08928_, _08927_, _01671_);
  and (_08929_, _08928_, _08926_);
  and (_08930_, _04636_, _01670_);
  or (_08931_, _08930_, _06973_);
  or (_08932_, _08931_, _08929_);
  or (_08933_, _08752_, _06974_);
  and (_08934_, _08933_, _05444_);
  and (_08935_, _08934_, _08932_);
  or (_08936_, _07500_, _07494_);
  nor (_08937_, _07501_, _05444_);
  and (_08938_, _08937_, _08936_);
  or (_08939_, _08938_, _08935_);
  and (_08940_, _08939_, _05442_);
  or (_08941_, _07661_, _03850_);
  nor (_08942_, _07662_, _05442_);
  and (_08943_, _08942_, _08941_);
  or (_08944_, _08943_, _07095_);
  or (_08945_, _08944_, _08940_);
  not (_08946_, _04347_);
  and (_08947_, _08730_, _08946_);
  nor (_08948_, _08730_, _08946_);
  nor (_08949_, _08948_, _08947_);
  or (_08950_, _08949_, _08078_);
  and (_08951_, _08950_, _07169_);
  and (_08952_, _08951_, _08945_);
  or (_08953_, _08952_, _07693_);
  or (_08954_, _07690_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_08955_, _08954_, _07684_);
  and (_08956_, _08955_, _08953_);
  and (_08957_, _04592_, _05429_);
  and (_08958_, _02958_, _02023_);
  or (_08959_, _08958_, _08957_);
  and (_08960_, _08959_, _07683_);
  or (_29641_, _08960_, _08956_);
  or (_08961_, _07690_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_08962_, _08961_, _07684_);
  and (_08963_, _05751_, _04501_);
  nor (_08964_, _05751_, _04501_);
  or (_08965_, _08964_, _08963_);
  and (_08966_, _08965_, _07095_);
  and (_08967_, _02413_, _01589_);
  nor (_08968_, _07634_, _07625_);
  or (_08969_, _08968_, _07635_);
  and (_08970_, _08969_, _05417_);
  and (_08971_, _04628_, _01660_);
  not (_08972_, \oc8051_golden_model_1.ACC [6]);
  nor (_08973_, _04501_, _08972_);
  and (_08974_, _04501_, _08972_);
  nor (_08975_, _08974_, _08973_);
  and (_08976_, _08975_, _07062_);
  nor (_08977_, _05330_, _05329_);
  and (_08978_, _08156_, _02264_);
  nor (_08979_, _08978_, _08977_);
  nor (_08980_, _08979_, _07271_);
  nand (_08981_, _04806_, _01950_);
  and (_08982_, _04099_, \oc8051_golden_model_1.P0 [6]);
  and (_08983_, _05189_, \oc8051_golden_model_1.P2 [6]);
  nor (_08984_, _08983_, _08982_);
  and (_08985_, _05195_, \oc8051_golden_model_1.P1 [6]);
  and (_08986_, _05191_, \oc8051_golden_model_1.P3 [6]);
  nor (_08987_, _08986_, _08985_);
  and (_08988_, _08987_, _08984_);
  and (_08989_, _08988_, _05318_);
  and (_08990_, _08989_, _05315_);
  and (_08991_, _08990_, _04454_);
  nor (_08992_, _08991_, _05330_);
  or (_08993_, _08992_, _06980_);
  nor (_08994_, _05495_, _04501_);
  nor (_08995_, _08994_, _05496_);
  nor (_08996_, _08995_, _06987_);
  or (_08997_, _07515_, _03748_);
  nor (_08998_, _07519_, _04074_);
  or (_08999_, _08998_, _07520_);
  and (_09000_, _08999_, _04557_);
  nor (_09001_, _04629_, _01625_);
  and (_09002_, _01625_, \oc8051_golden_model_1.ACC [6]);
  or (_09003_, _09002_, _09001_);
  and (_09004_, _09003_, _04709_);
  or (_09005_, _09004_, _04715_);
  or (_09006_, _09005_, _09000_);
  and (_09007_, _09006_, _06987_);
  and (_09008_, _09007_, _08997_);
  or (_09009_, _09008_, _08996_);
  and (_09010_, _09009_, _07513_);
  nand (_09011_, _08991_, _05331_);
  and (_09012_, _09011_, _06982_);
  or (_09013_, _09012_, _06363_);
  or (_09014_, _09013_, _09010_);
  nor (_09015_, _04628_, _01621_);
  nor (_09016_, _09015_, _07008_);
  and (_09017_, _09016_, _09014_);
  and (_09018_, _07008_, _07493_);
  or (_09019_, _09018_, _06979_);
  or (_09020_, _09019_, _09017_);
  and (_09021_, _09020_, _08993_);
  or (_09022_, _09021_, _01953_);
  nand (_09023_, _04806_, _01953_);
  and (_09024_, _09023_, _07546_);
  nand (_09025_, _09024_, _09022_);
  nor (_09026_, _08991_, _05331_);
  nand (_09027_, _09011_, _07023_);
  or (_09028_, _09027_, _09026_);
  nand (_09029_, _09028_, _09025_);
  and (_09030_, _09029_, _01632_);
  or (_09031_, _04629_, _01632_);
  nand (_09032_, _09031_, _01942_);
  or (_09033_, _09032_, _09030_);
  and (_09034_, _09033_, _08981_);
  or (_09035_, _09034_, _03273_);
  and (_09036_, _03748_, _01853_);
  nand (_09037_, _04805_, _03273_);
  or (_09038_, _09037_, _09036_);
  and (_09039_, _09038_, _07271_);
  and (_09040_, _09039_, _09035_);
  or (_09041_, _09040_, _08980_);
  and (_09042_, _09041_, _07270_);
  and (_09043_, _04628_, _01606_);
  or (_09044_, _09043_, _07039_);
  or (_09045_, _09044_, _09042_);
  nand (_09046_, _07039_, _04074_);
  and (_09047_, _09046_, _09045_);
  or (_09048_, _09047_, _07037_);
  or (_09049_, _07571_, _03748_);
  and (_09050_, _09049_, _07106_);
  and (_09051_, _09050_, _09048_);
  nor (_09052_, _04074_, _02962_);
  and (_09053_, _05540_, \oc8051_golden_model_1.TCON [6]);
  and (_09054_, _05544_, \oc8051_golden_model_1.PSW [6]);
  nor (_09055_, _09054_, _09053_);
  and (_09056_, _05556_, \oc8051_golden_model_1.P0INREG [6]);
  and (_09057_, _05558_, \oc8051_golden_model_1.SCON [6]);
  nor (_09058_, _09057_, _09056_);
  and (_09059_, _09058_, _09055_);
  and (_09060_, _05550_, \oc8051_golden_model_1.ACC [6]);
  and (_09061_, _05553_, \oc8051_golden_model_1.B [6]);
  nor (_09062_, _09061_, _09060_);
  and (_09063_, _05527_, \oc8051_golden_model_1.P1INREG [6]);
  and (_09064_, _05534_, \oc8051_golden_model_1.SBUF [6]);
  nor (_09065_, _09064_, _09063_);
  and (_09066_, _09065_, _09062_);
  and (_09067_, _09066_, _09059_);
  and (_09068_, _05567_, \oc8051_golden_model_1.PCON [6]);
  and (_09069_, _05569_, \oc8051_golden_model_1.DPH [6]);
  nor (_09070_, _09069_, _09068_);
  and (_09071_, _09070_, _09067_);
  and (_09072_, _05633_, \oc8051_golden_model_1.SP [6]);
  and (_09073_, _05578_, \oc8051_golden_model_1.TL1 [6]);
  nor (_09074_, _09073_, _09072_);
  and (_09075_, _05595_, \oc8051_golden_model_1.TH1 [6]);
  and (_09076_, _05629_, \oc8051_golden_model_1.TMOD [6]);
  nor (_09077_, _09076_, _09075_);
  and (_09078_, _09077_, _09074_);
  and (_09079_, _05576_, \oc8051_golden_model_1.DPL [6]);
  not (_09080_, _09079_);
  and (_09081_, _05603_, \oc8051_golden_model_1.IE [6]);
  and (_09082_, _05609_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_09083_, _09082_, _09081_);
  and (_09084_, _05615_, \oc8051_golden_model_1.P2INREG [6]);
  and (_09085_, _05619_, \oc8051_golden_model_1.IP [6]);
  nor (_09086_, _09085_, _09084_);
  and (_09087_, _09086_, _09083_);
  and (_09088_, _09087_, _09080_);
  and (_09089_, _05582_, \oc8051_golden_model_1.TL0 [6]);
  and (_09090_, _05587_, \oc8051_golden_model_1.TH0 [6]);
  nor (_09091_, _09090_, _09089_);
  and (_09092_, _09091_, _09088_);
  and (_09093_, _09092_, _09078_);
  and (_09094_, _09093_, _09071_);
  not (_09095_, _09094_);
  nor (_09096_, _09095_, _09052_);
  nor (_09097_, _09096_, _07042_);
  or (_09098_, _09097_, _02859_);
  or (_09099_, _09098_, _09051_);
  and (_09100_, _02859_, _01884_);
  nor (_09101_, _09100_, _06976_);
  and (_09102_, _09101_, _09099_);
  not (_09103_, _03025_);
  and (_09104_, _06976_, _09103_);
  or (_09105_, _09104_, _01650_);
  or (_09106_, _09105_, _09102_);
  and (_09107_, _04629_, _01650_);
  nor (_09108_, _09107_, _07061_);
  and (_09109_, _09108_, _09106_);
  nor (_09110_, _04501_, _03025_);
  and (_09111_, _04501_, _03025_);
  nor (_09112_, _09111_, _09110_);
  and (_09113_, _09112_, _07061_);
  or (_09114_, _09113_, _09109_);
  and (_09115_, _09114_, _07584_);
  or (_09116_, _09115_, _08976_);
  and (_09117_, _09116_, _07060_);
  and (_09118_, _09110_, _07059_);
  or (_09119_, _09118_, _09117_);
  and (_09120_, _09119_, _07058_);
  and (_09121_, _08973_, _07057_);
  or (_09122_, _09121_, _01666_);
  or (_09123_, _09122_, _09120_);
  and (_09124_, _04629_, _01666_);
  nor (_09125_, _09124_, _07598_);
  and (_09126_, _09125_, _09123_);
  nand (_09127_, _09111_, _07603_);
  and (_09128_, _09127_, _07107_);
  or (_09129_, _09128_, _09126_);
  nand (_09130_, _08974_, _07602_);
  and (_09131_, _09130_, _05157_);
  and (_09132_, _09131_, _09129_);
  or (_09133_, _09132_, _08971_);
  and (_09134_, _09133_, _08048_);
  nor (_09135_, _07115_, _02348_);
  not (_09136_, _08048_);
  nand (_09137_, _08999_, _09136_);
  nand (_09138_, _09137_, _09135_);
  or (_09139_, _09138_, _09134_);
  or (_09140_, _08999_, _09135_);
  and (_09141_, _09140_, _07623_);
  and (_09142_, _09141_, _09139_);
  or (_09143_, _09142_, _08970_);
  and (_09144_, _09143_, _07622_);
  nor (_09145_, _08995_, _07622_);
  or (_09146_, _09145_, _02023_);
  or (_09147_, _09146_, _09144_);
  nand (_09148_, _03029_, _02023_);
  and (_09149_, _09148_, _01671_);
  and (_09150_, _09149_, _09147_);
  and (_09151_, _04628_, _01670_);
  or (_09152_, _09151_, _06973_);
  or (_09153_, _09152_, _09150_);
  or (_09154_, _08977_, _06974_);
  and (_09155_, _09154_, _05444_);
  and (_09156_, _09155_, _09153_);
  and (_09157_, _02804_, _01589_);
  nor (_09158_, _07501_, _07493_);
  nor (_09159_, _09158_, _07502_);
  and (_09160_, _09159_, _07651_);
  or (_09161_, _09160_, _09157_);
  or (_09162_, _09161_, _09156_);
  not (_09163_, _09157_);
  nor (_09164_, _07662_, _03748_);
  nor (_09165_, _09164_, _07663_);
  or (_09166_, _09165_, _09163_);
  and (_09167_, _09166_, _09162_);
  or (_09168_, _09167_, _08967_);
  not (_09169_, _08967_);
  or (_09170_, _09165_, _09169_);
  and (_09171_, _09170_, _08078_);
  and (_09172_, _09171_, _09168_);
  nor (_09173_, _09172_, _08966_);
  nand (_09174_, _09173_, _07690_);
  and (_09175_, _09174_, _08962_);
  and (_09176_, _02945_, _02023_);
  nor (_09177_, _04586_, _02023_);
  or (_09178_, _09177_, _09176_);
  and (_09179_, _09178_, _07683_);
  or (_29642_, _09179_, _09175_);
  or (_09180_, _07690_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_09181_, _09180_, _07684_);
  nand (_09182_, _07690_, _07671_);
  and (_09183_, _09182_, _09181_);
  and (_09184_, _07683_, _07677_);
  or (_29643_, _09184_, _09183_);
  and (_09185_, _07687_, _07265_);
  and (_09186_, _09185_, _07686_);
  not (_09187_, _09186_);
  or (_09188_, _09187_, _07878_);
  and (_09189_, _07682_, _03399_);
  not (_09190_, _09189_);
  or (_09191_, _09186_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_09192_, _09191_, _09190_);
  and (_09193_, _09192_, _09188_);
  and (_09194_, _09189_, _07883_);
  or (_29726_[0], _09194_, _09193_);
  or (_09195_, _09190_, _08086_);
  and (_09196_, _09186_, _08081_);
  nor (_09197_, _09186_, _03343_);
  or (_09198_, _09197_, _09189_);
  or (_09199_, _09198_, _09196_);
  and (_29726_[1], _09199_, _09195_);
  or (_09200_, _09190_, _08295_);
  nand (_09201_, _09186_, _08288_);
  or (_09202_, _09186_, _03203_);
  and (_09203_, _09202_, _09190_);
  nand (_09204_, _09203_, _09201_);
  and (_29726_[2], _09204_, _09200_);
  and (_09205_, _09186_, _08510_);
  nor (_09206_, _09186_, _03405_);
  or (_09207_, _09206_, _09189_);
  or (_09208_, _09207_, _09205_);
  or (_09209_, _09190_, _08515_);
  and (_29726_[3], _09209_, _09208_);
  or (_09210_, _09187_, _08735_);
  or (_09211_, _09186_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_09212_, _09211_, _09190_);
  and (_09213_, _09212_, _09210_);
  and (_09214_, _09189_, _08742_);
  or (_29726_[4], _09214_, _09213_);
  or (_09215_, _09187_, _08952_);
  or (_09216_, _09186_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_09217_, _09216_, _09190_);
  and (_09218_, _09217_, _09215_);
  and (_09219_, _09189_, _08959_);
  or (_29726_[5], _09219_, _09218_);
  nor (_09220_, _09173_, _07168_);
  and (_09221_, _09220_, _26505_);
  and (_09222_, _09221_, _25964_);
  or (_09223_, _09187_, _09222_);
  or (_09224_, _09186_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_09225_, _09224_, _09190_);
  and (_09226_, _09225_, _09223_);
  and (_09227_, _09189_, _09178_);
  or (_29726_[6], _09227_, _09226_);
  or (_09228_, _09187_, _07672_);
  or (_09229_, _09186_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_09230_, _09229_, _09190_);
  and (_09231_, _09230_, _09228_);
  and (_09232_, _09189_, _07677_);
  or (_29726_[7], _09232_, _09231_);
  not (_09233_, _07098_);
  and (_09234_, _07266_, _09233_);
  and (_09235_, _09234_, _07686_);
  not (_09236_, _09235_);
  or (_09237_, _09236_, _07878_);
  and (_09238_, _07682_, _03190_);
  not (_09239_, _09238_);
  or (_09240_, _09235_, \oc8051_golden_model_1.IRAM[2] [0]);
  and (_09241_, _09240_, _09239_);
  and (_09242_, _09241_, _09237_);
  and (_09243_, _09238_, _07883_);
  or (_29727_[0], _09243_, _09242_);
  or (_09244_, _09236_, _08081_);
  or (_09245_, _09235_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_09246_, _09245_, _09239_);
  and (_09247_, _09246_, _09244_);
  and (_09248_, _08086_, _07475_);
  and (_09249_, _09248_, _09238_);
  or (_29727_[1], _09249_, _09247_);
  or (_09250_, _09236_, _08288_);
  or (_09251_, _09235_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_09252_, _09251_, _09239_);
  and (_09253_, _09252_, _09250_);
  and (_09254_, _08295_, _07475_);
  and (_09255_, _09254_, _09238_);
  or (_29727_[2], _09255_, _09253_);
  or (_09256_, _09236_, _08510_);
  or (_09257_, _09235_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_09258_, _09257_, _09239_);
  and (_09259_, _09258_, _09256_);
  and (_09260_, _09238_, _08515_);
  or (_29727_[3], _09260_, _09259_);
  or (_09261_, _09236_, _08735_);
  or (_09262_, _09235_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_09263_, _09262_, _09239_);
  and (_09264_, _09263_, _09261_);
  and (_09265_, _08742_, _07475_);
  and (_09266_, _09265_, _09238_);
  or (_29727_[4], _09266_, _09264_);
  or (_09267_, _09236_, _08952_);
  or (_09268_, _09235_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_09269_, _09268_, _09239_);
  and (_09270_, _09269_, _09267_);
  and (_09271_, _08959_, _07475_);
  and (_09272_, _09271_, _09238_);
  or (_29727_[5], _09272_, _09270_);
  or (_09273_, _09236_, _09222_);
  or (_09274_, _09235_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_09275_, _09274_, _09239_);
  and (_09276_, _09275_, _09273_);
  and (_09277_, _09178_, _07475_);
  and (_09278_, _09277_, _09238_);
  or (_29727_[6], _09278_, _09276_);
  or (_09279_, _09236_, _07672_);
  or (_09280_, _09235_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_09281_, _09280_, _09239_);
  and (_09282_, _09281_, _09279_);
  and (_09283_, _09238_, _07678_);
  or (_29727_[7], _09283_, _09282_);
  not (_09284_, _07265_);
  and (_09285_, _07687_, _09284_);
  and (_09286_, _07686_, _09285_);
  not (_09287_, _09286_);
  or (_09288_, _09287_, _07878_);
  and (_09289_, _07681_, _07477_);
  not (_09290_, _09289_);
  or (_09291_, _09286_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_09292_, _09291_, _09290_);
  and (_09293_, _09292_, _09288_);
  and (_09294_, _07883_, _07475_);
  and (_09295_, _09294_, _09289_);
  or (_29728_[0], _09295_, _09293_);
  or (_09296_, _09287_, _08081_);
  or (_09297_, _09286_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_09298_, _09297_, _09290_);
  and (_09299_, _09298_, _09296_);
  and (_09300_, _09289_, _09248_);
  or (_29728_[1], _09300_, _09299_);
  or (_09301_, _09287_, _08288_);
  or (_09302_, _09286_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_09303_, _09302_, _09290_);
  and (_09304_, _09303_, _09301_);
  and (_09305_, _09289_, _09254_);
  or (_29728_[2], _09305_, _09304_);
  and (_09306_, _07686_, _07267_);
  or (_09307_, _09306_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_09308_, _09307_, _09290_);
  not (_09309_, _09306_);
  or (_09310_, _09309_, _08510_);
  and (_09311_, _09310_, _09308_);
  and (_09312_, _08515_, _07475_);
  and (_09313_, _09312_, _09289_);
  or (_29728_[3], _09313_, _09311_);
  or (_09314_, _09306_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_09315_, _09314_, _09290_);
  or (_09316_, _09309_, _08735_);
  and (_09317_, _09316_, _09315_);
  and (_09318_, _09289_, _09265_);
  or (_29728_[4], _09318_, _09317_);
  or (_09319_, _09306_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_09320_, _09319_, _09290_);
  or (_09321_, _09309_, _08952_);
  and (_09322_, _09321_, _09320_);
  and (_09323_, _09289_, _09271_);
  or (_29728_[5], _09323_, _09322_);
  or (_09324_, _09306_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_09325_, _09324_, _09290_);
  or (_09326_, _09309_, _09222_);
  and (_09327_, _09326_, _09325_);
  and (_09328_, _09289_, _09277_);
  or (_29728_[6], _09328_, _09327_);
  or (_09329_, _09306_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_09330_, _09329_, _09290_);
  or (_09331_, _09309_, _07672_);
  and (_09332_, _09331_, _09330_);
  and (_09333_, _09289_, _07678_);
  or (_29728_[7], _09333_, _09332_);
  and (_09334_, _07469_, _07379_);
  and (_09335_, _09334_, _07688_);
  not (_09336_, _09335_);
  or (_09337_, _09336_, _07878_);
  not (_09338_, _07484_);
  and (_09339_, _07680_, _09338_);
  and (_09340_, _09339_, _07478_);
  not (_09341_, _09340_);
  or (_09342_, _09335_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_09343_, _09342_, _09341_);
  and (_09344_, _09343_, _09337_);
  and (_09345_, _09340_, _09294_);
  or (_29729_[0], _09345_, _09344_);
  or (_09346_, _09336_, _08081_);
  or (_09347_, _09335_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_09348_, _09347_, _09341_);
  and (_09349_, _09348_, _09346_);
  and (_09350_, _09340_, _09248_);
  or (_29729_[1], _09350_, _09349_);
  or (_09351_, _09336_, _08288_);
  or (_09352_, _09335_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_09353_, _09352_, _09341_);
  and (_09354_, _09353_, _09351_);
  and (_09355_, _09340_, _09254_);
  or (_29729_[2], _09355_, _09354_);
  or (_09356_, _09336_, _08510_);
  or (_09357_, _09335_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_09358_, _09357_, _09341_);
  and (_09359_, _09358_, _09356_);
  and (_09360_, _09340_, _09312_);
  or (_29729_[3], _09360_, _09359_);
  or (_09361_, _09336_, _08735_);
  or (_09362_, _09335_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_09363_, _09362_, _09341_);
  and (_09364_, _09363_, _09361_);
  and (_09365_, _09340_, _09265_);
  or (_29729_[4], _09365_, _09364_);
  or (_09366_, _09336_, _08952_);
  or (_09367_, _09335_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_09368_, _09367_, _09341_);
  and (_09369_, _09368_, _09366_);
  and (_09370_, _09340_, _09271_);
  or (_29729_[5], _09370_, _09369_);
  or (_09371_, _09336_, _09222_);
  or (_09372_, _09335_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_09373_, _09372_, _09341_);
  and (_09374_, _09373_, _09371_);
  and (_09375_, _09340_, _09277_);
  or (_29729_[6], _09375_, _09374_);
  or (_09376_, _09336_, _07672_);
  or (_09377_, _09335_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_09378_, _09377_, _09341_);
  and (_09379_, _09378_, _09376_);
  and (_09380_, _09340_, _07678_);
  or (_29729_[7], _09380_, _09379_);
  and (_09381_, _09334_, _09185_);
  not (_09382_, _09381_);
  or (_09383_, _09382_, _07878_);
  and (_09384_, _09339_, _03399_);
  not (_09385_, _09384_);
  or (_09386_, _09381_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_09387_, _09386_, _09385_);
  and (_09388_, _09387_, _09383_);
  and (_09389_, _09384_, _09294_);
  or (_29690_, _09389_, _09388_);
  or (_09390_, _09382_, _08081_);
  or (_09391_, _09381_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_09392_, _09391_, _09385_);
  and (_09393_, _09392_, _09390_);
  and (_09394_, _09384_, _09248_);
  or (_29691_, _09394_, _09393_);
  or (_09395_, _09382_, _08288_);
  or (_09396_, _09381_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_09397_, _09396_, _09385_);
  and (_09398_, _09397_, _09395_);
  and (_09399_, _09384_, _09254_);
  or (_29692_, _09399_, _09398_);
  or (_09400_, _09382_, _08510_);
  or (_09401_, _09381_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_09402_, _09401_, _09385_);
  and (_09403_, _09402_, _09400_);
  and (_09404_, _09384_, _09312_);
  or (_29693_, _09404_, _09403_);
  or (_09405_, _09382_, _08735_);
  or (_09406_, _09381_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_09407_, _09406_, _09385_);
  and (_09408_, _09407_, _09405_);
  and (_09409_, _09384_, _09265_);
  or (_29694_, _09409_, _09408_);
  or (_09410_, _09382_, _08952_);
  or (_09411_, _09381_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_09412_, _09411_, _09385_);
  and (_09413_, _09412_, _09410_);
  and (_09414_, _09384_, _09271_);
  or (_29695_, _09414_, _09413_);
  and (_09415_, _09381_, _09222_);
  nor (_09416_, _09381_, _03709_);
  or (_09417_, _09416_, _09384_);
  or (_09418_, _09417_, _09415_);
  or (_09419_, _09385_, _09277_);
  and (_29696_, _09419_, _09418_);
  or (_09420_, _09382_, _07672_);
  or (_09421_, _09381_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_09422_, _09421_, _09385_);
  and (_09423_, _09422_, _09420_);
  and (_09424_, _09384_, _07678_);
  or (_29697_, _09424_, _09423_);
  and (_09425_, _09334_, _09234_);
  not (_09426_, _09425_);
  or (_09427_, _09426_, _07878_);
  and (_09428_, _09339_, _03190_);
  not (_09429_, _09428_);
  or (_09430_, _09425_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_09431_, _09430_, _09429_);
  and (_09432_, _09431_, _09427_);
  and (_09433_, _09428_, _09294_);
  or (_29698_, _09433_, _09432_);
  or (_09434_, _09426_, _08081_);
  or (_09435_, _09425_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_09436_, _09435_, _09429_);
  and (_09437_, _09436_, _09434_);
  and (_09438_, _09428_, _09248_);
  or (_29699_, _09438_, _09437_);
  or (_09439_, _09426_, _08288_);
  or (_09440_, _09425_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_09441_, _09440_, _09429_);
  and (_09442_, _09441_, _09439_);
  and (_09443_, _09428_, _09254_);
  or (_29700_, _09443_, _09442_);
  or (_09444_, _09426_, _08510_);
  or (_09445_, _09425_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_09446_, _09445_, _09429_);
  and (_09447_, _09446_, _09444_);
  and (_09448_, _09428_, _09312_);
  or (_29701_, _09448_, _09447_);
  or (_09449_, _09426_, _08735_);
  or (_09450_, _09425_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_09451_, _09450_, _09429_);
  and (_09452_, _09451_, _09449_);
  and (_09453_, _09428_, _09265_);
  or (_29702_, _09453_, _09452_);
  or (_09454_, _09426_, _08952_);
  or (_09455_, _09425_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_09456_, _09455_, _09429_);
  and (_09457_, _09456_, _09454_);
  and (_09458_, _09428_, _09271_);
  or (_29703_, _09458_, _09457_);
  or (_09459_, _09426_, _09222_);
  or (_09460_, _09425_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_09461_, _09460_, _09429_);
  and (_09462_, _09461_, _09459_);
  and (_09463_, _09428_, _09277_);
  or (_29704_, _09463_, _09462_);
  or (_09464_, _09426_, _07672_);
  or (_09465_, _09425_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_09466_, _09465_, _09429_);
  and (_09467_, _09466_, _09464_);
  and (_09468_, _09428_, _07678_);
  or (_29705_, _09468_, _09467_);
  and (_09469_, _09339_, _07477_);
  not (_09470_, _09469_);
  and (_09471_, _09334_, _07267_);
  or (_09472_, _09471_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_09473_, _09472_, _09470_);
  not (_09474_, _09471_);
  or (_09475_, _09474_, _07878_);
  and (_09476_, _09475_, _09473_);
  and (_09477_, _09469_, _09294_);
  or (_29706_, _09477_, _09476_);
  or (_09478_, _09470_, _09248_);
  and (_09479_, _09471_, _08081_);
  nor (_09480_, _09471_, _03355_);
  or (_09481_, _09480_, _09469_);
  or (_09482_, _09481_, _09479_);
  and (_29707_, _09482_, _09478_);
  or (_09483_, _09471_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_09484_, _09483_, _09470_);
  or (_09485_, _09474_, _08288_);
  and (_09486_, _09485_, _09484_);
  and (_09487_, _09469_, _09254_);
  or (_29708_, _09487_, _09486_);
  or (_09488_, _09471_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_09489_, _09488_, _09470_);
  or (_09490_, _09474_, _08510_);
  and (_09491_, _09490_, _09489_);
  and (_09492_, _09469_, _09312_);
  or (_29709_, _09492_, _09491_);
  or (_09493_, _09471_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_09494_, _09493_, _09470_);
  or (_09495_, _09474_, _08735_);
  and (_09496_, _09495_, _09494_);
  and (_09497_, _09469_, _09265_);
  or (_29710_, _09497_, _09496_);
  or (_09498_, _09471_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_09499_, _09498_, _09470_);
  or (_09500_, _09474_, _08952_);
  and (_09501_, _09500_, _09499_);
  and (_09502_, _09469_, _09271_);
  or (_29711_, _09502_, _09501_);
  or (_09503_, _09474_, _09222_);
  or (_09504_, _09471_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_09505_, _09504_, _09470_);
  and (_09506_, _09505_, _09503_);
  and (_09507_, _09469_, _09277_);
  or (_29712_, _09507_, _09506_);
  or (_09508_, _09471_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_09509_, _09508_, _09470_);
  or (_09510_, _09474_, _07672_);
  and (_09511_, _09510_, _09509_);
  and (_09512_, _09469_, _07678_);
  or (_29713_, _09512_, _09511_);
  and (_09513_, _07685_, _07468_);
  and (_09514_, _09513_, _07688_);
  not (_09515_, _09514_);
  or (_09516_, _09515_, _07878_);
  or (_09517_, _09514_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand (_09518_, _07485_, _07479_);
  and (_09519_, _09518_, _09517_);
  and (_09520_, _09519_, _09516_);
  not (_09521_, _07481_);
  and (_09522_, _07485_, _09521_);
  and (_09523_, _09522_, _07478_);
  and (_09524_, _09523_, _09294_);
  or (_29714_, _09524_, _09520_);
  or (_09525_, _09515_, _08081_);
  nor (_09526_, _09514_, \oc8051_golden_model_1.IRAM[8] [1]);
  nor (_09527_, _09526_, _09523_);
  and (_09528_, _09527_, _09525_);
  and (_09529_, _09523_, _09248_);
  or (_29715_, _09529_, _09528_);
  or (_09530_, _09515_, _08288_);
  nor (_09531_, _09514_, \oc8051_golden_model_1.IRAM[8] [2]);
  nor (_09532_, _09531_, _09523_);
  and (_09533_, _09532_, _09530_);
  and (_09534_, _09523_, _09254_);
  or (_29716_, _09534_, _09533_);
  or (_09535_, _09515_, _08510_);
  or (_09536_, _09514_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_09537_, _09536_, _09518_);
  and (_09538_, _09537_, _09535_);
  and (_09539_, _09523_, _09312_);
  or (_29717_, _09539_, _09538_);
  or (_09540_, _09515_, _08735_);
  or (_09541_, _09514_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_09542_, _09541_, _09518_);
  and (_09543_, _09542_, _09540_);
  and (_09544_, _09523_, _09265_);
  or (_29718_, _09544_, _09543_);
  or (_09545_, _09515_, _08952_);
  or (_09546_, _09514_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_09547_, _09546_, _09518_);
  and (_09548_, _09547_, _09545_);
  and (_09549_, _09523_, _09271_);
  or (_29719_, _09549_, _09548_);
  or (_09550_, _09515_, _09222_);
  or (_09551_, _09514_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_09552_, _09551_, _09518_);
  and (_09553_, _09552_, _09550_);
  and (_09554_, _09523_, _09277_);
  or (_29720_, _09554_, _09553_);
  or (_09555_, _09515_, _07672_);
  or (_09556_, _09514_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_09557_, _09556_, _09518_);
  and (_09558_, _09557_, _09555_);
  and (_09559_, _09523_, _07678_);
  or (_29721_, _09559_, _09558_);
  and (_09560_, _09513_, _09185_);
  not (_09561_, _09560_);
  or (_09562_, _09561_, _07878_);
  and (_09563_, _09522_, _03399_);
  not (_09564_, _09563_);
  or (_09565_, _09560_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_09566_, _09565_, _09564_);
  and (_09567_, _09566_, _09562_);
  and (_09568_, _09563_, _09294_);
  or (_29722_, _09568_, _09567_);
  or (_09569_, _09561_, _08081_);
  or (_09570_, _09560_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_09571_, _09570_, _09564_);
  and (_09572_, _09571_, _09569_);
  and (_09573_, _09563_, _09248_);
  or (_29723_, _09573_, _09572_);
  or (_09574_, _09561_, _08288_);
  or (_09575_, _09560_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_09576_, _09575_, _09564_);
  and (_09577_, _09576_, _09574_);
  and (_09578_, _09563_, _09254_);
  or (_29724_, _09578_, _09577_);
  or (_09579_, _09561_, _08510_);
  nand (_09580_, _07485_, _07273_);
  or (_09581_, _09560_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_09582_, _09581_, _09580_);
  and (_09583_, _09582_, _09579_);
  and (_09584_, _09563_, _09312_);
  or (_29725_, _09584_, _09583_);
  or (_09585_, _09561_, _08735_);
  or (_09586_, _09560_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_09587_, _09586_, _09580_);
  and (_09588_, _09587_, _09585_);
  and (_09589_, _09563_, _09265_);
  or (_29730_[4], _09589_, _09588_);
  or (_09590_, _09561_, _08952_);
  or (_09591_, _09560_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_09592_, _09591_, _09580_);
  and (_09593_, _09592_, _09590_);
  and (_09594_, _09563_, _09271_);
  or (_29730_[5], _09594_, _09593_);
  or (_09595_, _09561_, _09222_);
  or (_09596_, _09560_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_09597_, _09596_, _09580_);
  and (_09598_, _09597_, _09595_);
  and (_09599_, _09563_, _09277_);
  or (_29730_[6], _09599_, _09598_);
  and (_09600_, _09560_, _07672_);
  nand (_09601_, _09561_, \oc8051_golden_model_1.IRAM[9] [7]);
  nand (_09602_, _09601_, _09580_);
  or (_09603_, _09602_, _09600_);
  or (_09604_, _09564_, _07678_);
  and (_29730_[7], _09604_, _09603_);
  and (_09605_, _09513_, _09234_);
  and (_09606_, _09605_, _07878_);
  nor (_09607_, _09605_, _03312_);
  or (_09608_, _09607_, _09606_);
  nor (_09609_, _07474_, _02441_);
  and (_09610_, _09609_, _26505_);
  and (_09611_, _09610_, _25964_);
  nor (_09612_, _07474_, \oc8051_golden_model_1.SP [1]);
  and (_09613_, _09612_, _26505_);
  and (_09614_, _09613_, _25964_);
  not (_09615_, _09614_);
  nor (_09616_, _09615_, _09611_);
  nor (_09617_, _09521_, _07474_);
  and (_09618_, _09617_, _26505_);
  and (_09619_, _09618_, _25964_);
  nor (_09620_, _09338_, _07474_);
  and (_09621_, _09620_, _26505_);
  and (_09622_, _09621_, _25964_);
  not (_09623_, _09622_);
  nor (_09624_, _09623_, _09619_);
  nand (_09625_, _09624_, _09616_);
  and (_09626_, _09625_, _09608_);
  and (_09627_, _09522_, _03190_);
  and (_09628_, _09627_, _09294_);
  or (_25573_, _09628_, _09626_);
  not (_09629_, _09605_);
  or (_09630_, _09629_, _08081_);
  not (_09631_, _09627_);
  or (_09632_, _09605_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_09633_, _09632_, _09631_);
  and (_09634_, _09633_, _09630_);
  and (_09635_, _09627_, _09248_);
  or (_25574_, _09635_, _09634_);
  or (_09636_, _09629_, _08288_);
  or (_09637_, _09605_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_09638_, _09637_, _09631_);
  and (_09639_, _09638_, _09636_);
  and (_09640_, _09627_, _09254_);
  or (_29644_, _09640_, _09639_);
  or (_09641_, _09629_, _08510_);
  or (_09642_, _09605_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_09643_, _09642_, _09631_);
  and (_09644_, _09643_, _09641_);
  and (_09645_, _09627_, _09312_);
  or (_29645_, _09645_, _09644_);
  or (_09646_, _09629_, _08735_);
  or (_09647_, _09605_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_09648_, _09647_, _09631_);
  and (_09649_, _09648_, _09646_);
  and (_09650_, _09627_, _09265_);
  or (_29646_, _09650_, _09649_);
  or (_09651_, _09629_, _08952_);
  or (_09652_, _09605_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_09653_, _09652_, _09631_);
  and (_09654_, _09653_, _09651_);
  and (_09655_, _09627_, _09271_);
  or (_29647_, _09655_, _09654_);
  or (_09656_, _09629_, _09222_);
  or (_09657_, _09605_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_09658_, _09657_, _09631_);
  and (_09659_, _09658_, _09656_);
  and (_09660_, _09627_, _09277_);
  or (_29648_, _09660_, _09659_);
  or (_09661_, _09629_, _07672_);
  or (_09662_, _09605_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_09663_, _09662_, _09631_);
  and (_09664_, _09663_, _09661_);
  and (_09665_, _09627_, _07678_);
  or (_29649_, _09665_, _09664_);
  and (_09666_, _09513_, _09285_);
  not (_09667_, _09666_);
  or (_09668_, _09667_, _07878_);
  and (_09669_, _09522_, _07477_);
  not (_09670_, _09669_);
  or (_09671_, _09666_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_09672_, _09671_, _09670_);
  and (_09673_, _09672_, _09668_);
  and (_09674_, _09669_, _09294_);
  or (_29650_, _09674_, _09673_);
  or (_09675_, _09667_, _08081_);
  or (_09676_, _09666_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_09677_, _09676_, _09670_);
  and (_09678_, _09677_, _09675_);
  and (_09679_, _09669_, _09248_);
  or (_29651_, _09679_, _09678_);
  or (_09680_, _09667_, _08288_);
  or (_09681_, _09666_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_09682_, _09681_, _09670_);
  and (_09683_, _09682_, _09680_);
  and (_09684_, _09669_, _09254_);
  or (_29652_, _09684_, _09683_);
  nor (_09685_, _09666_, \oc8051_golden_model_1.IRAM[11] [3]);
  nor (_09686_, _09667_, _08510_);
  or (_09687_, _09686_, _09685_);
  nand (_09688_, _09687_, _09670_);
  or (_09689_, _09670_, _09312_);
  and (_29653_, _09689_, _09688_);
  and (_09690_, _09513_, _07267_);
  or (_09691_, _09690_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_09692_, _09691_, _09670_);
  not (_09693_, _09690_);
  or (_09694_, _09693_, _08735_);
  and (_09695_, _09694_, _09692_);
  and (_09696_, _09669_, _09265_);
  or (_29654_, _09696_, _09695_);
  or (_09697_, _09690_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_09698_, _09697_, _09670_);
  or (_09699_, _09693_, _08952_);
  and (_09700_, _09699_, _09698_);
  and (_09701_, _09669_, _09271_);
  or (_29655_, _09701_, _09700_);
  or (_09702_, _09690_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_09703_, _09702_, _09670_);
  or (_09704_, _09693_, _09222_);
  and (_09705_, _09704_, _09703_);
  and (_09706_, _09669_, _09277_);
  or (_29656_, _09706_, _09705_);
  nor (_09707_, _09666_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor (_09708_, _09667_, _07672_);
  or (_09709_, _09708_, _09707_);
  nand (_09710_, _09709_, _09670_);
  or (_09711_, _09670_, _07678_);
  and (_29657_, _09711_, _09710_);
  not (_09712_, _07468_);
  and (_09713_, _07685_, _09712_);
  and (_09714_, _07688_, _09713_);
  not (_09715_, _09714_);
  or (_09716_, _09715_, _07878_);
  and (_09717_, _07486_, _07478_);
  not (_09718_, _09717_);
  or (_09719_, _09714_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_09720_, _09719_, _09718_);
  and (_09721_, _09720_, _09716_);
  and (_09722_, _09717_, _09294_);
  or (_29658_, _09722_, _09721_);
  or (_09723_, _09715_, _08081_);
  or (_09724_, _09714_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_09725_, _09724_, _09718_);
  and (_09726_, _09725_, _09723_);
  and (_09727_, _09717_, _09248_);
  or (_29659_, _09727_, _09726_);
  or (_09728_, _09715_, _08288_);
  or (_09729_, _09714_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_09730_, _09729_, _09718_);
  and (_09731_, _09730_, _09728_);
  and (_09732_, _09717_, _09254_);
  or (_29660_, _09732_, _09731_);
  and (_09733_, _07688_, _07471_);
  or (_09734_, _09733_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_09735_, _09734_, _09718_);
  or (_09736_, _09715_, _08510_);
  and (_09737_, _09736_, _09735_);
  and (_09738_, _09717_, _09312_);
  or (_29661_, _09738_, _09737_);
  or (_09739_, _09733_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_09740_, _09739_, _09718_);
  or (_09741_, _09715_, _08735_);
  and (_09742_, _09741_, _09740_);
  and (_09743_, _09717_, _09265_);
  or (_29662_, _09743_, _09742_);
  or (_09744_, _09733_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_09745_, _09744_, _09718_);
  or (_09746_, _09715_, _08952_);
  and (_09747_, _09746_, _09745_);
  and (_09748_, _09717_, _09271_);
  or (_29663_, _09748_, _09747_);
  or (_09749_, _09733_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_09750_, _09749_, _09718_);
  or (_09751_, _09715_, _09222_);
  and (_09752_, _09751_, _09750_);
  and (_09753_, _09717_, _09277_);
  or (_29664_, _09753_, _09752_);
  or (_09754_, _09733_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_09755_, _09754_, _09718_);
  or (_09756_, _09715_, _07672_);
  and (_09757_, _09756_, _09755_);
  and (_09758_, _09717_, _07678_);
  or (_29665_, _09758_, _09757_);
  and (_09759_, _09185_, _09713_);
  not (_09760_, _09759_);
  or (_09761_, _09760_, _07878_);
  and (_09762_, _07486_, _03399_);
  not (_09763_, _09762_);
  or (_09764_, _09759_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_09765_, _09764_, _09763_);
  and (_09766_, _09765_, _09761_);
  and (_09767_, _09762_, _09294_);
  or (_29666_, _09767_, _09766_);
  or (_09768_, _09760_, _08081_);
  or (_09769_, _09759_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_09770_, _09769_, _09763_);
  and (_09771_, _09770_, _09768_);
  and (_09772_, _09762_, _09248_);
  or (_29667_, _09772_, _09771_);
  or (_09773_, _09760_, _08288_);
  or (_09774_, _09759_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_09775_, _09774_, _09763_);
  and (_09776_, _09775_, _09773_);
  and (_09777_, _09762_, _09254_);
  or (_29668_, _09777_, _09776_);
  or (_09778_, _09759_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_09779_, _09778_, _09763_);
  or (_09780_, _09760_, _08510_);
  and (_09781_, _09780_, _09779_);
  and (_09782_, _09762_, _09312_);
  or (_29669_, _09782_, _09781_);
  or (_09783_, _09759_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_09784_, _09783_, _09763_);
  or (_09785_, _09760_, _08735_);
  and (_09786_, _09785_, _09784_);
  and (_09787_, _09762_, _09265_);
  or (_29670_, _09787_, _09786_);
  or (_09788_, _09759_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_09789_, _09788_, _09763_);
  or (_09790_, _09760_, _08952_);
  and (_09791_, _09790_, _09789_);
  and (_09792_, _09762_, _09271_);
  or (_29671_, _09792_, _09791_);
  nor (_09793_, _09760_, _09222_);
  nor (_09794_, _09759_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_09795_, _09794_, _09793_);
  nor (_09796_, _09795_, _09762_);
  and (_09797_, _09762_, _09277_);
  or (_29672_, _09797_, _09796_);
  or (_09798_, _09759_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_09799_, _09798_, _09763_);
  or (_09800_, _09760_, _07672_);
  and (_09801_, _09800_, _09799_);
  and (_09802_, _09762_, _07678_);
  or (_29673_, _09802_, _09801_);
  and (_09803_, _09234_, _09713_);
  not (_09804_, _09803_);
  or (_09805_, _09804_, _07878_);
  and (_09806_, _07486_, _03190_);
  not (_09807_, _09806_);
  or (_09808_, _09803_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_09809_, _09808_, _09807_);
  and (_09810_, _09809_, _09805_);
  and (_09811_, _09806_, _09294_);
  or (_29674_, _09811_, _09810_);
  or (_09812_, _09804_, _08081_);
  or (_09813_, _09803_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_09814_, _09813_, _09807_);
  and (_09815_, _09814_, _09812_);
  and (_09816_, _09806_, _09248_);
  or (_29675_, _09816_, _09815_);
  or (_09817_, _09804_, _08288_);
  or (_09818_, _09803_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_09819_, _09818_, _09807_);
  and (_09820_, _09819_, _09817_);
  and (_09821_, _09806_, _09254_);
  or (_29676_, _09821_, _09820_);
  and (_09822_, _09234_, _07471_);
  or (_09823_, _09822_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_09824_, _09823_, _09807_);
  or (_09825_, _09804_, _08510_);
  and (_09826_, _09825_, _09824_);
  and (_09827_, _09806_, _09312_);
  or (_29677_, _09827_, _09826_);
  or (_09828_, _09822_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_09829_, _09828_, _09807_);
  or (_09830_, _09804_, _08735_);
  and (_09831_, _09830_, _09829_);
  and (_09832_, _09806_, _09265_);
  or (_29678_, _09832_, _09831_);
  or (_09833_, _09822_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_09834_, _09833_, _09807_);
  or (_09835_, _09804_, _08952_);
  and (_09836_, _09835_, _09834_);
  and (_09837_, _09806_, _09271_);
  or (_29679_, _09837_, _09836_);
  or (_09838_, _09822_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_09839_, _09838_, _09807_);
  or (_09840_, _09804_, _09222_);
  and (_09841_, _09840_, _09839_);
  and (_09842_, _09806_, _09277_);
  or (_29680_, _09842_, _09841_);
  or (_09843_, _09822_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_09844_, _09843_, _09807_);
  or (_09845_, _09804_, _07672_);
  and (_09846_, _09845_, _09844_);
  and (_09847_, _09806_, _07678_);
  or (_29681_, _09847_, _09846_);
  or (_09848_, _07472_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_09849_, _09848_, _07488_);
  or (_09850_, _07878_, _07490_);
  and (_09851_, _09850_, _09849_);
  and (_09852_, _09294_, _07487_);
  or (_29682_, _09852_, _09851_);
  or (_09853_, _07472_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_09854_, _09853_, _07488_);
  or (_09855_, _08081_, _07490_);
  and (_09856_, _09855_, _09854_);
  and (_09857_, _09248_, _07487_);
  or (_29683_, _09857_, _09856_);
  and (_09858_, _09713_, _09285_);
  not (_09859_, _09858_);
  or (_09860_, _08288_, _09859_);
  or (_09861_, _09858_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_09862_, _09861_, _07488_);
  and (_09863_, _09862_, _09860_);
  and (_09864_, _09254_, _07487_);
  or (_29684_, _09864_, _09863_);
  or (_09865_, _08510_, _07490_);
  or (_09866_, _07472_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_09867_, _09866_, _07488_);
  and (_09868_, _09867_, _09865_);
  and (_09869_, _09312_, _07487_);
  or (_29685_, _09869_, _09868_);
  or (_09870_, _07472_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_09871_, _09870_, _07488_);
  or (_09872_, _08735_, _07490_);
  and (_09873_, _09872_, _09871_);
  and (_09874_, _09265_, _07487_);
  or (_29686_, _09874_, _09873_);
  or (_09875_, _07472_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_09876_, _09875_, _07488_);
  or (_09877_, _08952_, _07490_);
  and (_09878_, _09877_, _09876_);
  and (_09879_, _09271_, _07487_);
  or (_29687_, _09879_, _09878_);
  or (_09880_, _07472_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_09881_, _09880_, _07488_);
  or (_09882_, _09222_, _07490_);
  and (_09883_, _09882_, _09881_);
  and (_09884_, _09277_, _07487_);
  or (_29688_, _09884_, _09883_);
  nand (_09885_, \oc8051_golden_model_1.B [0], _25964_);
  nor (_27719_, _09885_, _26505_);
  nand (_09886_, \oc8051_golden_model_1.B [1], _25964_);
  nor (_27720_, _09886_, _26505_);
  nand (_09887_, \oc8051_golden_model_1.B [2], _25964_);
  nor (_27723_, _09887_, _26505_);
  nand (_09888_, \oc8051_golden_model_1.B [3], _25964_);
  nor (_27724_, _09888_, _26505_);
  nand (_09889_, \oc8051_golden_model_1.B [4], _25964_);
  nor (_27725_, _09889_, _26505_);
  nand (_09890_, \oc8051_golden_model_1.B [5], _25964_);
  nor (_27726_, _09890_, _26505_);
  nand (_09891_, \oc8051_golden_model_1.B [6], _25964_);
  nor (_27727_, _09891_, _26505_);
  or (_09892_, _01679_, rst);
  nor (_27729_, _09892_, _26505_);
  or (_09893_, _01705_, rst);
  nor (_27732_, _09893_, _26505_);
  or (_09894_, _08234_, rst);
  nor (_27733_, _09894_, _26505_);
  or (_09895_, _01732_, rst);
  nor (_27734_, _09895_, _26505_);
  or (_09896_, _08524_, rst);
  nor (_27735_, _09896_, _26505_);
  or (_09897_, _08747_, rst);
  nor (_27736_, _09897_, _26505_);
  or (_09898_, _08972_, rst);
  nor (_27737_, _09898_, _26505_);
  nand (_09899_, \oc8051_golden_model_1.DPL [0], _25964_);
  nor (_27739_, _09899_, _26505_);
  nand (_09900_, \oc8051_golden_model_1.DPL [1], _25964_);
  nor (_27740_, _09900_, _26505_);
  nand (_09901_, \oc8051_golden_model_1.DPL [2], _25964_);
  nor (_27741_, _09901_, _26505_);
  nand (_09902_, \oc8051_golden_model_1.DPL [3], _25964_);
  nor (_27742_, _09902_, _26505_);
  nand (_09903_, \oc8051_golden_model_1.DPL [4], _25964_);
  nor (_27743_, _09903_, _26505_);
  nand (_09904_, \oc8051_golden_model_1.DPL [5], _25964_);
  nor (_27744_, _09904_, _26505_);
  nand (_09905_, \oc8051_golden_model_1.DPL [6], _25964_);
  nor (_27745_, _09905_, _26505_);
  nand (_09906_, \oc8051_golden_model_1.DPH [0], _25964_);
  nor (_27750_, _09906_, _26505_);
  nand (_09907_, \oc8051_golden_model_1.DPH [1], _25964_);
  nor (_27751_, _09907_, _26505_);
  nand (_09908_, \oc8051_golden_model_1.DPH [2], _25964_);
  nor (_27752_, _09908_, _26505_);
  nand (_09909_, \oc8051_golden_model_1.DPH [3], _25964_);
  nor (_27753_, _09909_, _26505_);
  nand (_09910_, \oc8051_golden_model_1.DPH [4], _25964_);
  nor (_27754_, _09910_, _26505_);
  nand (_09911_, \oc8051_golden_model_1.DPH [5], _25964_);
  nor (_27755_, _09911_, _26505_);
  nand (_09912_, \oc8051_golden_model_1.DPH [6], _25964_);
  nor (_27756_, _09912_, _26505_);
  not (_09913_, \oc8051_golden_model_1.IE [0]);
  nor (_09914_, _04183_, _09913_);
  nor (_09915_, _04405_, _06864_);
  nor (_09916_, _09915_, _09914_);
  nor (_09917_, _09916_, _01595_);
  and (_09918_, _04183_, _03677_);
  nor (_09919_, _09914_, _05513_);
  not (_09920_, _09919_);
  nor (_09921_, _09920_, _09918_);
  nor (_09922_, _05186_, _09913_);
  and (_09923_, _07725_, _05186_);
  nor (_09924_, _09923_, _09922_);
  nor (_09925_, _09924_, _02223_);
  and (_09926_, _09916_, _01969_);
  and (_09927_, _04183_, \oc8051_golden_model_1.ACC [0]);
  nor (_09928_, _09927_, _09914_);
  nor (_09929_, _09928_, _05488_);
  nor (_09930_, _04571_, _09913_);
  or (_09931_, _09930_, _01969_);
  nor (_09932_, _09931_, _09929_);
  or (_09933_, _09932_, _06233_);
  nor (_09934_, _09933_, _09926_);
  and (_09935_, _04183_, _03334_);
  nor (_09936_, _09935_, _09914_);
  nor (_09937_, _09936_, _05487_);
  or (_09938_, _09937_, _01963_);
  or (_09939_, _09938_, _09934_);
  nor (_09940_, _09939_, _09925_);
  and (_09941_, _09928_, _01963_);
  nor (_09942_, _09941_, _01957_);
  not (_09943_, _09942_);
  nor (_09944_, _09943_, _09940_);
  and (_09945_, _09914_, _01957_);
  or (_09946_, _09945_, _09944_);
  and (_09947_, _09946_, _04885_);
  nor (_09948_, _09916_, _04885_);
  or (_09949_, _09948_, _09947_);
  nor (_09950_, _09949_, _01924_);
  nor (_09951_, _07759_, _06901_);
  or (_09952_, _09922_, _01925_);
  nor (_09953_, _09952_, _09951_);
  or (_09954_, _09953_, _04950_);
  or (_09955_, _09954_, _09950_);
  or (_09956_, _09936_, _06397_);
  and (_09957_, _09956_, _05513_);
  and (_09958_, _09957_, _09955_);
  nor (_09959_, _09958_, _09921_);
  nor (_09960_, _09959_, _01602_);
  nor (_09961_, _07815_, _06864_);
  or (_09962_, _09914_, _01923_);
  nor (_09963_, _09962_, _09961_);
  or (_09964_, _09963_, _02019_);
  nor (_09965_, _09964_, _09960_);
  and (_09966_, _04183_, _05531_);
  nor (_09967_, _09966_, _09914_);
  nand (_09968_, _09967_, _05049_);
  and (_09969_, _09968_, _06278_);
  nor (_09970_, _09969_, _09965_);
  and (_09971_, _07829_, _04183_);
  nor (_09972_, _09971_, _09914_);
  and (_09973_, _09972_, _02018_);
  nor (_09974_, _09973_, _09970_);
  and (_09975_, _09974_, _02136_);
  and (_09976_, _07834_, _04183_);
  nor (_09977_, _09976_, _09914_);
  nor (_09978_, _09977_, _02136_);
  or (_09979_, _09978_, _09975_);
  and (_09980_, _09979_, _05076_);
  or (_09981_, _09967_, _05076_);
  nor (_09982_, _09981_, _09915_);
  nor (_09983_, _09982_, _09980_);
  nor (_09984_, _09983_, _02130_);
  nor (_09985_, _09914_, _04405_);
  or (_09986_, _09985_, _02131_);
  nor (_09987_, _09986_, _09928_);
  or (_09988_, _09987_, _02016_);
  nor (_09989_, _09988_, _09984_);
  nor (_09990_, _07828_, _06864_);
  nor (_09991_, _09990_, _09914_);
  and (_09992_, _09991_, _02016_);
  nor (_09993_, _09992_, _09989_);
  and (_09994_, _09993_, _05474_);
  nor (_09995_, _07696_, _06864_);
  nor (_09996_, _09995_, _09914_);
  nor (_09997_, _09996_, _05474_);
  or (_09998_, _09997_, _09994_);
  and (_09999_, _09998_, _02168_);
  nor (_10000_, _09916_, _02168_);
  nor (_10001_, _10000_, _02025_);
  not (_10002_, _10001_);
  nor (_10003_, _10002_, _09999_);
  nor (_10004_, _09914_, _02377_);
  nor (_10005_, _10004_, _10003_);
  and (_10006_, _10005_, _01595_);
  nor (_10007_, _10006_, _09917_);
  nand (_10008_, _10007_, _26505_);
  or (_10009_, _26505_, \oc8051_golden_model_1.IE [0]);
  and (_10010_, _10009_, _25964_);
  and (_27757_, _10010_, _10008_);
  not (_10011_, \oc8051_golden_model_1.IE [1]);
  nor (_10012_, _04183_, _10011_);
  and (_10013_, _04183_, _03613_);
  or (_10014_, _10013_, _10012_);
  and (_10015_, _10014_, _04951_);
  nor (_10016_, _07953_, _06901_);
  nor (_10017_, _05186_, _10011_);
  or (_10018_, _10017_, _01925_);
  or (_10019_, _10018_, _10016_);
  nor (_10020_, _04183_, \oc8051_golden_model_1.IE [1]);
  and (_10021_, _07909_, _04183_);
  nor (_10022_, _10021_, _10020_);
  nor (_10023_, _10022_, _02438_);
  and (_10024_, _04183_, _01705_);
  nor (_10025_, _10024_, _10020_);
  and (_10026_, _10025_, _04571_);
  nor (_10027_, _04571_, _10011_);
  or (_10028_, _10027_, _01969_);
  nor (_10029_, _10028_, _10026_);
  or (_10030_, _10029_, _06233_);
  nor (_10031_, _10030_, _10023_);
  nor (_10032_, _06864_, _03393_);
  nor (_10033_, _10032_, _10012_);
  nor (_10034_, _10033_, _05487_);
  and (_10035_, _07920_, _05186_);
  nor (_10036_, _10035_, _10017_);
  nor (_10037_, _10036_, _02223_);
  nor (_10038_, _10037_, _10034_);
  nand (_10039_, _10038_, _01964_);
  or (_10040_, _10039_, _10031_);
  or (_10041_, _10025_, _01964_);
  and (_10042_, _10041_, _10040_);
  and (_10043_, _10042_, _06229_);
  and (_10044_, _07907_, _05186_);
  nor (_10045_, _10044_, _10017_);
  nor (_10046_, _10045_, _06229_);
  or (_10047_, _10046_, _10043_);
  and (_10048_, _10047_, _04885_);
  nor (_10049_, _10017_, _07935_);
  or (_10050_, _10049_, _04885_);
  nor (_10051_, _10050_, _10036_);
  or (_10052_, _10051_, _01924_);
  or (_10053_, _10052_, _10048_);
  and (_10054_, _10053_, _10019_);
  nor (_10055_, _10054_, _04950_);
  and (_10056_, _10033_, _04950_);
  or (_10057_, _10056_, _04951_);
  nor (_10058_, _10057_, _10055_);
  or (_10059_, _10058_, _10015_);
  and (_10060_, _10059_, _01923_);
  nor (_10061_, _08009_, _06864_);
  nor (_10062_, _10061_, _10012_);
  nor (_10063_, _10062_, _01923_);
  nor (_10064_, _10063_, _10060_);
  nor (_10065_, _10064_, _06278_);
  and (_10066_, _04183_, _02676_);
  not (_10067_, _10066_);
  nor (_10068_, _10020_, _04979_);
  and (_10069_, _10068_, _10067_);
  nor (_10070_, _10069_, _10065_);
  not (_10071_, _10012_);
  nand (_10072_, _08023_, _04183_);
  and (_10073_, _10072_, _10071_);
  or (_10074_, _10073_, _05049_);
  and (_10075_, _10074_, _10070_);
  nor (_10076_, _10075_, _02135_);
  not (_10077_, _10020_);
  nor (_10078_, _08029_, _06864_);
  nor (_10079_, _10078_, _02136_);
  and (_10080_, _10079_, _10077_);
  nor (_10081_, _10080_, _10076_);
  nor (_10082_, _10081_, _02039_);
  nor (_10083_, _07893_, _06864_);
  nor (_10084_, _10083_, _05076_);
  and (_10085_, _10084_, _10077_);
  nor (_10086_, _10085_, _10082_);
  nor (_10087_, _10086_, _02130_);
  and (_10088_, _10071_, _04452_);
  nor (_10089_, _10088_, _02131_);
  and (_10090_, _10089_, _10025_);
  nor (_10091_, _10090_, _10087_);
  nor (_10092_, _10091_, _02128_);
  and (_10093_, _10066_, _04452_);
  nor (_10094_, _10093_, _05104_);
  nand (_10095_, _10024_, _04452_);
  and (_10096_, _10095_, _02126_);
  or (_10097_, _10096_, _10094_);
  and (_10098_, _10097_, _10077_);
  or (_10099_, _10098_, _02164_);
  nor (_10100_, _10099_, _10092_);
  nor (_10101_, _10022_, _02168_);
  or (_10102_, _10101_, _02025_);
  nor (_10103_, _10102_, _10100_);
  nor (_10104_, _10045_, _02377_);
  or (_10105_, _10104_, _01594_);
  nor (_10106_, _10105_, _10103_);
  nor (_10107_, _10021_, _10012_);
  and (_10108_, _10107_, _01594_);
  nor (_10109_, _10108_, _10106_);
  or (_10110_, _10109_, _26506_);
  or (_10111_, _26505_, \oc8051_golden_model_1.IE [1]);
  and (_10112_, _10111_, _25964_);
  and (_27758_, _10112_, _10110_);
  not (_10113_, \oc8051_golden_model_1.IE [2]);
  nor (_10114_, _04183_, _10113_);
  and (_10115_, _04183_, _05563_);
  nor (_10116_, _10115_, _10114_);
  and (_10117_, _10116_, _02019_);
  nor (_10118_, _06864_, _03272_);
  nor (_10119_, _10118_, _10114_);
  and (_10120_, _10119_, _04950_);
  nor (_10121_, _08095_, _06864_);
  nor (_10122_, _10121_, _10114_);
  and (_10123_, _10122_, _01969_);
  and (_10124_, _04183_, \oc8051_golden_model_1.ACC [2]);
  nor (_10125_, _10124_, _10114_);
  nor (_10126_, _10125_, _05488_);
  nor (_10127_, _04571_, _10113_);
  or (_10128_, _10127_, _01969_);
  nor (_10129_, _10128_, _10126_);
  or (_10130_, _10129_, _06233_);
  nor (_10131_, _10130_, _10123_);
  nor (_10132_, _10119_, _05487_);
  nor (_10133_, _05186_, _10113_);
  and (_10134_, _08111_, _05186_);
  nor (_10135_, _10134_, _10133_);
  nor (_10136_, _10135_, _02223_);
  nor (_10137_, _10136_, _10132_);
  nand (_10138_, _10137_, _01964_);
  or (_10139_, _10138_, _10131_);
  nand (_10140_, _10125_, _01963_);
  and (_10141_, _10140_, _10139_);
  nor (_10142_, _10141_, _01957_);
  and (_10143_, _08109_, _05186_);
  nor (_10144_, _10143_, _10133_);
  and (_10145_, _10144_, _01957_);
  or (_10146_, _10145_, _01946_);
  nor (_10147_, _10146_, _10142_);
  nor (_10148_, _10133_, _08139_);
  or (_10149_, _10148_, _04885_);
  nor (_10150_, _10149_, _10135_);
  or (_10151_, _10150_, _10147_);
  and (_10152_, _10151_, _01925_);
  nor (_10153_, _08158_, _06901_);
  nor (_10154_, _10133_, _10153_);
  nor (_10155_, _10154_, _01925_);
  or (_10156_, _10155_, _04950_);
  nor (_10157_, _10156_, _10152_);
  nor (_10158_, _10157_, _10120_);
  nor (_10159_, _10158_, _04951_);
  and (_10160_, _04183_, _03564_);
  nor (_10161_, _10114_, _05513_);
  not (_10162_, _10161_);
  nor (_10163_, _10162_, _10160_);
  or (_10164_, _10163_, _01602_);
  nor (_10165_, _10164_, _10159_);
  nor (_10166_, _08216_, _06864_);
  nor (_10167_, _10166_, _10114_);
  nor (_10168_, _10167_, _01923_);
  or (_10169_, _10168_, _02019_);
  nor (_10170_, _10169_, _10165_);
  nor (_10171_, _10170_, _10117_);
  or (_10172_, _10171_, _02018_);
  and (_10173_, _08230_, _04183_);
  or (_10174_, _10173_, _10114_);
  or (_10175_, _10174_, _05049_);
  and (_10176_, _10175_, _02136_);
  and (_10177_, _10176_, _10172_);
  and (_10178_, _08237_, _04183_);
  nor (_10179_, _10178_, _10114_);
  nor (_10180_, _10179_, _02136_);
  nor (_10181_, _10180_, _10177_);
  nor (_10182_, _10181_, _02039_);
  nor (_10183_, _10114_, _05739_);
  not (_10184_, _10183_);
  nor (_10185_, _10116_, _05076_);
  and (_10186_, _10185_, _10184_);
  nor (_10187_, _10186_, _10182_);
  nor (_10188_, _10187_, _02130_);
  or (_10189_, _10183_, _02131_);
  nor (_10190_, _10189_, _10125_);
  or (_10191_, _10190_, _02016_);
  nor (_10192_, _10191_, _10188_);
  nor (_10193_, _08229_, _06864_);
  nor (_10194_, _10193_, _10114_);
  and (_10195_, _10194_, _02016_);
  nor (_10196_, _10195_, _10192_);
  and (_10197_, _10196_, _05474_);
  nor (_10198_, _08236_, _06864_);
  nor (_10199_, _10198_, _10114_);
  nor (_10200_, _10199_, _05474_);
  or (_10201_, _10200_, _10197_);
  and (_10202_, _10201_, _02168_);
  nor (_10203_, _10122_, _02168_);
  or (_10204_, _10203_, _02025_);
  or (_10205_, _10204_, _10202_);
  nand (_10206_, _10144_, _02025_);
  and (_10207_, _10206_, _10205_);
  nor (_10208_, _10207_, _01594_);
  and (_10209_, _08285_, _04183_);
  nor (_10210_, _10209_, _10114_);
  and (_10211_, _10210_, _01594_);
  nor (_10212_, _10211_, _10208_);
  or (_10213_, _10212_, _26506_);
  or (_10214_, _26505_, \oc8051_golden_model_1.IE [2]);
  and (_10215_, _10214_, _25964_);
  and (_27759_, _10215_, _10213_);
  not (_10216_, \oc8051_golden_model_1.IE [3]);
  nor (_10217_, _04183_, _10216_);
  and (_10218_, _04183_, _05529_);
  nor (_10219_, _10218_, _10217_);
  and (_10220_, _10219_, _02019_);
  nor (_10221_, _06864_, _03473_);
  nor (_10222_, _10221_, _10217_);
  and (_10223_, _10222_, _04950_);
  nor (_10224_, _08308_, _06901_);
  nor (_10225_, _05186_, _10216_);
  or (_10226_, _10225_, _01925_);
  or (_10227_, _10226_, _10224_);
  nor (_10228_, _08337_, _06864_);
  nor (_10229_, _10228_, _10217_);
  and (_10230_, _10229_, _01969_);
  and (_10231_, _04183_, \oc8051_golden_model_1.ACC [3]);
  nor (_10232_, _10231_, _10217_);
  nor (_10233_, _10232_, _05488_);
  nor (_10234_, _04571_, _10216_);
  or (_10235_, _10234_, _01969_);
  nor (_10236_, _10235_, _10233_);
  or (_10237_, _10236_, _06233_);
  nor (_10238_, _10237_, _10230_);
  nor (_10239_, _10222_, _05487_);
  and (_10240_, _08341_, _05186_);
  nor (_10241_, _10240_, _10225_);
  nor (_10242_, _10241_, _02223_);
  nor (_10243_, _10242_, _10239_);
  nand (_10244_, _10243_, _01964_);
  or (_10245_, _10244_, _10238_);
  nand (_10246_, _10232_, _01963_);
  and (_10247_, _10246_, _10245_);
  and (_10248_, _10247_, _06229_);
  and (_10249_, _08324_, _05186_);
  nor (_10250_, _10249_, _10225_);
  nor (_10251_, _10250_, _06229_);
  or (_10252_, _10251_, _10248_);
  and (_10253_, _10252_, _04885_);
  nor (_10254_, _10225_, _08357_);
  or (_10255_, _10241_, _04885_);
  nor (_10256_, _10255_, _10254_);
  or (_10257_, _10256_, _01924_);
  or (_10258_, _10257_, _10253_);
  and (_10259_, _10258_, _10227_);
  nor (_10260_, _10259_, _04950_);
  nor (_10261_, _10260_, _10223_);
  nor (_10262_, _10261_, _04951_);
  and (_10263_, _04183_, _03516_);
  nor (_10264_, _10217_, _05513_);
  not (_10265_, _10264_);
  nor (_10266_, _10265_, _10263_);
  or (_10267_, _10266_, _01602_);
  nor (_10268_, _10267_, _10262_);
  nor (_10269_, _08425_, _06864_);
  nor (_10270_, _10269_, _10217_);
  nor (_10271_, _10270_, _01923_);
  or (_10272_, _10271_, _02019_);
  nor (_10273_, _10272_, _10268_);
  nor (_10274_, _10273_, _10220_);
  or (_10275_, _10274_, _02018_);
  and (_10276_, _08441_, _04183_);
  or (_10277_, _10276_, _10217_);
  or (_10278_, _10277_, _05049_);
  and (_10279_, _10278_, _02136_);
  and (_10280_, _10279_, _10275_);
  and (_10281_, _08304_, _04183_);
  nor (_10282_, _10281_, _10217_);
  nor (_10283_, _10282_, _02136_);
  nor (_10284_, _10283_, _10280_);
  nor (_10285_, _10284_, _02039_);
  nor (_10286_, _10217_, _05737_);
  not (_10287_, _10286_);
  nor (_10288_, _10219_, _05076_);
  and (_10289_, _10288_, _10287_);
  nor (_10290_, _10289_, _10285_);
  nor (_10291_, _10290_, _02130_);
  or (_10292_, _10286_, _02131_);
  nor (_10293_, _10292_, _10232_);
  or (_10294_, _10293_, _02016_);
  nor (_10295_, _10294_, _10291_);
  nor (_10296_, _08440_, _06864_);
  nor (_10297_, _10296_, _10217_);
  and (_10298_, _10297_, _02016_);
  nor (_10299_, _10298_, _10295_);
  and (_10300_, _10299_, _05474_);
  nor (_10301_, _08303_, _06864_);
  nor (_10302_, _10301_, _10217_);
  nor (_10303_, _10302_, _05474_);
  or (_10304_, _10303_, _10300_);
  and (_10305_, _10304_, _02168_);
  nor (_10306_, _10229_, _02168_);
  or (_10307_, _10306_, _02025_);
  or (_10308_, _10307_, _10305_);
  nand (_10309_, _10250_, _02025_);
  and (_10310_, _10309_, _10308_);
  nor (_10311_, _10310_, _01594_);
  and (_10312_, _08507_, _04183_);
  nor (_10313_, _10312_, _10217_);
  and (_10314_, _10313_, _01594_);
  nor (_10315_, _10314_, _10311_);
  or (_10316_, _10315_, _26506_);
  or (_10317_, _26505_, \oc8051_golden_model_1.IE [3]);
  and (_10318_, _10317_, _25964_);
  and (_27760_, _10318_, _10316_);
  not (_10319_, \oc8051_golden_model_1.IE [4]);
  nor (_10320_, _04183_, _10319_);
  and (_10321_, _04183_, _05524_);
  nor (_10322_, _10321_, _10320_);
  and (_10323_, _10322_, _02019_);
  nor (_10324_, _06864_, _04024_);
  nor (_10325_, _10324_, _10320_);
  and (_10326_, _10325_, _04950_);
  nor (_10327_, _05186_, _10319_);
  nor (_10328_, _10327_, _08581_);
  and (_10329_, _08565_, _05186_);
  nor (_10330_, _10329_, _10327_);
  or (_10331_, _10330_, _04885_);
  nor (_10332_, _10331_, _10328_);
  nor (_10333_, _08548_, _06864_);
  nor (_10334_, _10333_, _10320_);
  and (_10335_, _10334_, _01969_);
  and (_10336_, _04183_, \oc8051_golden_model_1.ACC [4]);
  nor (_10337_, _10336_, _10320_);
  nor (_10338_, _10337_, _05488_);
  nor (_10339_, _04571_, _10319_);
  or (_10340_, _10339_, _01969_);
  nor (_10341_, _10340_, _10338_);
  or (_10342_, _10341_, _06233_);
  nor (_10343_, _10342_, _10335_);
  nor (_10344_, _10325_, _05487_);
  nor (_10345_, _10330_, _02223_);
  nor (_10346_, _10345_, _10344_);
  nand (_10347_, _10346_, _01964_);
  or (_10348_, _10347_, _10343_);
  nand (_10349_, _10337_, _01963_);
  and (_10350_, _10349_, _10348_);
  and (_10351_, _10350_, _06229_);
  and (_10352_, _08544_, _05186_);
  nor (_10353_, _10352_, _10327_);
  nor (_10354_, _10353_, _06229_);
  or (_10355_, _10354_, _10351_);
  and (_10356_, _10355_, _04885_);
  nor (_10357_, _10356_, _10332_);
  nor (_10358_, _10357_, _01924_);
  nor (_10359_, _08607_, _06901_);
  nor (_10360_, _10359_, _10327_);
  nor (_10361_, _10360_, _01925_);
  nor (_10362_, _10361_, _04950_);
  not (_10363_, _10362_);
  nor (_10364_, _10363_, _10358_);
  nor (_10365_, _10364_, _10326_);
  nor (_10366_, _10365_, _04951_);
  and (_10367_, _04183_, _03903_);
  nor (_10368_, _10320_, _05513_);
  not (_10369_, _10368_);
  nor (_10370_, _10369_, _10367_);
  or (_10371_, _10370_, _01602_);
  nor (_10372_, _10371_, _10366_);
  nor (_10373_, _08663_, _06864_);
  nor (_10374_, _10373_, _10320_);
  nor (_10375_, _10374_, _01923_);
  or (_10376_, _10375_, _02019_);
  nor (_10377_, _10376_, _10372_);
  nor (_10378_, _10377_, _10323_);
  or (_10379_, _10378_, _02018_);
  and (_10380_, _08531_, _04183_);
  or (_10381_, _10380_, _10320_);
  or (_10382_, _10381_, _05049_);
  and (_10383_, _10382_, _02136_);
  and (_10384_, _10383_, _10379_);
  and (_10385_, _08527_, _04183_);
  nor (_10386_, _10385_, _10320_);
  nor (_10387_, _10386_, _02136_);
  nor (_10388_, _10387_, _10384_);
  nor (_10389_, _10388_, _02039_);
  nor (_10390_, _10320_, _08729_);
  not (_10391_, _10390_);
  nor (_10392_, _10322_, _05076_);
  and (_10393_, _10392_, _10391_);
  nor (_10394_, _10393_, _10389_);
  nor (_10395_, _10394_, _02130_);
  or (_10396_, _10390_, _02131_);
  nor (_10397_, _10396_, _10337_);
  or (_10398_, _10397_, _02016_);
  nor (_10399_, _10398_, _10395_);
  nor (_10400_, _08530_, _06864_);
  nor (_10401_, _10400_, _10320_);
  and (_10402_, _10401_, _02016_);
  nor (_10403_, _10402_, _10399_);
  and (_10404_, _10403_, _05474_);
  nor (_10405_, _08526_, _06864_);
  nor (_10406_, _10405_, _10320_);
  nor (_10407_, _10406_, _05474_);
  or (_10408_, _10407_, _10404_);
  and (_10409_, _10408_, _02168_);
  nor (_10410_, _10334_, _02168_);
  or (_10411_, _10410_, _02025_);
  or (_10412_, _10411_, _10409_);
  nand (_10413_, _10353_, _02025_);
  and (_10414_, _10413_, _10412_);
  nor (_10415_, _10414_, _01594_);
  and (_10416_, _08732_, _04183_);
  nor (_10417_, _10416_, _10320_);
  and (_10418_, _10417_, _01594_);
  nor (_10419_, _10418_, _10415_);
  or (_10420_, _10419_, _26506_);
  or (_10421_, _26505_, \oc8051_golden_model_1.IE [4]);
  and (_10422_, _10421_, _25964_);
  and (_27761_, _10422_, _10420_);
  not (_10423_, \oc8051_golden_model_1.IE [5]);
  nor (_10424_, _04183_, _10423_);
  and (_10425_, _04183_, _05548_);
  nor (_10426_, _10425_, _10424_);
  and (_10427_, _10426_, _02019_);
  nor (_10428_, _06864_, _03976_);
  nor (_10429_, _10428_, _10424_);
  and (_10430_, _10429_, _04950_);
  nor (_10431_, _08771_, _06864_);
  nor (_10432_, _10431_, _10424_);
  and (_10433_, _10432_, _01969_);
  and (_10434_, _04183_, \oc8051_golden_model_1.ACC [5]);
  nor (_10435_, _10434_, _10424_);
  nor (_10436_, _10435_, _05488_);
  nor (_10437_, _04571_, _10423_);
  or (_10438_, _10437_, _01969_);
  nor (_10439_, _10438_, _10436_);
  or (_10440_, _10439_, _06233_);
  nor (_10441_, _10440_, _10433_);
  nor (_10442_, _10429_, _05487_);
  nor (_10443_, _05186_, _10423_);
  and (_10444_, _08785_, _05186_);
  nor (_10445_, _10444_, _10443_);
  nor (_10446_, _10445_, _02223_);
  nor (_10447_, _10446_, _10442_);
  nand (_10448_, _10447_, _01964_);
  or (_10449_, _10448_, _10441_);
  nand (_10450_, _10435_, _01963_);
  and (_10451_, _10450_, _10449_);
  and (_10452_, _10451_, _06229_);
  and (_10453_, _08768_, _05186_);
  nor (_10454_, _10453_, _10443_);
  nor (_10455_, _10454_, _06229_);
  or (_10456_, _10455_, _10452_);
  and (_10457_, _10456_, _04885_);
  and (_10458_, _08802_, _05186_);
  nor (_10459_, _10458_, _10443_);
  nor (_10460_, _10459_, _04885_);
  nor (_10461_, _10460_, _10457_);
  nor (_10462_, _10461_, _01924_);
  nor (_10463_, _08754_, _06901_);
  nor (_10464_, _10463_, _10443_);
  nor (_10465_, _10464_, _01925_);
  nor (_10466_, _10465_, _04950_);
  not (_10467_, _10466_);
  nor (_10468_, _10467_, _10462_);
  nor (_10469_, _10468_, _10430_);
  nor (_10470_, _10469_, _04951_);
  and (_10471_, _04183_, _03850_);
  nor (_10472_, _10424_, _05513_);
  not (_10473_, _10472_);
  nor (_10474_, _10473_, _10471_);
  or (_10475_, _10474_, _01602_);
  nor (_10476_, _10475_, _10470_);
  nor (_10477_, _08874_, _06864_);
  nor (_10478_, _10477_, _10424_);
  nor (_10479_, _10478_, _01923_);
  or (_10480_, _10479_, _02019_);
  nor (_10481_, _10480_, _10476_);
  nor (_10482_, _10481_, _10427_);
  or (_10483_, _10482_, _02018_);
  and (_10484_, _08890_, _04183_);
  or (_10485_, _10484_, _10424_);
  or (_10486_, _10485_, _05049_);
  and (_10487_, _10486_, _02136_);
  and (_10488_, _10487_, _10483_);
  and (_10489_, _08750_, _04183_);
  nor (_10490_, _10489_, _10424_);
  nor (_10491_, _10490_, _02136_);
  nor (_10492_, _10491_, _10488_);
  nor (_10493_, _10492_, _02039_);
  nor (_10494_, _10424_, _08946_);
  not (_10495_, _10494_);
  nor (_10496_, _10426_, _05076_);
  and (_10497_, _10496_, _10495_);
  nor (_10498_, _10497_, _10493_);
  nor (_10499_, _10498_, _02130_);
  or (_10500_, _10494_, _02131_);
  nor (_10501_, _10500_, _10435_);
  or (_10502_, _10501_, _02016_);
  nor (_10503_, _10502_, _10499_);
  nor (_10504_, _08889_, _06864_);
  nor (_10505_, _10504_, _10424_);
  and (_10506_, _10505_, _02016_);
  nor (_10507_, _10506_, _10503_);
  and (_10508_, _10507_, _05474_);
  nor (_10509_, _08749_, _06864_);
  nor (_10510_, _10509_, _10424_);
  nor (_10511_, _10510_, _05474_);
  or (_10512_, _10511_, _10508_);
  and (_10513_, _10512_, _02168_);
  nor (_10514_, _10432_, _02168_);
  or (_10515_, _10514_, _02025_);
  or (_10516_, _10515_, _10513_);
  nand (_10517_, _10454_, _02025_);
  and (_10518_, _10517_, _10516_);
  nor (_10519_, _10518_, _01594_);
  and (_10520_, _08949_, _04183_);
  nor (_10521_, _10520_, _10424_);
  and (_10522_, _10521_, _01594_);
  nor (_10523_, _10522_, _10519_);
  or (_10524_, _10523_, _26506_);
  or (_10525_, _26505_, \oc8051_golden_model_1.IE [5]);
  and (_10526_, _10525_, _25964_);
  and (_27764_, _10526_, _10524_);
  not (_10527_, \oc8051_golden_model_1.IE [6]);
  nor (_10528_, _04183_, _10527_);
  and (_10529_, _04183_, _03748_);
  or (_10530_, _10529_, _10528_);
  and (_10531_, _10530_, _04951_);
  nor (_10532_, _05186_, _10527_);
  not (_10533_, _10532_);
  and (_10534_, _10533_, _09026_);
  and (_10535_, _09011_, _05186_);
  nor (_10536_, _10535_, _10532_);
  or (_10537_, _10536_, _04885_);
  nor (_10538_, _10537_, _10534_);
  nor (_10539_, _08995_, _06864_);
  nor (_10540_, _10539_, _10528_);
  and (_10541_, _10540_, _01969_);
  and (_10542_, _04183_, \oc8051_golden_model_1.ACC [6]);
  nor (_10543_, _10542_, _10528_);
  nor (_10544_, _10543_, _05488_);
  nor (_10545_, _04571_, _10527_);
  or (_10546_, _10545_, _01969_);
  nor (_10547_, _10546_, _10544_);
  or (_10548_, _10547_, _06233_);
  nor (_10549_, _10548_, _10541_);
  nor (_10550_, _06864_, _04074_);
  nor (_10551_, _10550_, _10528_);
  nor (_10552_, _10551_, _05487_);
  nor (_10553_, _10536_, _02223_);
  nor (_10554_, _10553_, _10552_);
  nand (_10555_, _10554_, _01964_);
  or (_10556_, _10555_, _10549_);
  nand (_10557_, _10543_, _01963_);
  and (_10558_, _10557_, _10556_);
  and (_10559_, _10558_, _06229_);
  and (_10560_, _08992_, _05186_);
  nor (_10561_, _10560_, _10532_);
  nor (_10562_, _10561_, _06229_);
  or (_10563_, _10562_, _10559_);
  and (_10564_, _10563_, _04885_);
  nor (_10565_, _10564_, _10538_);
  nor (_10566_, _10565_, _01924_);
  nor (_10567_, _08979_, _06901_);
  nor (_10568_, _10567_, _10532_);
  nor (_10569_, _10568_, _01925_);
  nor (_10570_, _10569_, _04950_);
  not (_10571_, _10570_);
  nor (_10572_, _10571_, _10566_);
  and (_10573_, _10551_, _04950_);
  or (_10574_, _10573_, _04951_);
  nor (_10575_, _10574_, _10572_);
  or (_10576_, _10575_, _10531_);
  and (_10577_, _10576_, _01923_);
  nor (_10578_, _09096_, _06864_);
  nor (_10579_, _10578_, _10528_);
  nor (_10580_, _10579_, _01923_);
  or (_10581_, _10580_, _06278_);
  or (_10582_, _10581_, _10577_);
  and (_10583_, _09112_, _04183_);
  or (_10584_, _10528_, _05049_);
  or (_10585_, _10584_, _10583_);
  and (_10586_, _04183_, _09103_);
  nor (_10587_, _10586_, _10528_);
  and (_10588_, _10587_, _02019_);
  nor (_10589_, _10588_, _02135_);
  and (_10590_, _10589_, _10585_);
  and (_10591_, _10590_, _10582_);
  and (_10592_, _08975_, _04183_);
  nor (_10593_, _10592_, _10528_);
  nor (_10594_, _10593_, _02136_);
  nor (_10595_, _10594_, _10591_);
  nor (_10596_, _10595_, _02039_);
  nor (_10597_, _10528_, _05735_);
  not (_10598_, _10597_);
  nor (_10599_, _10587_, _05076_);
  and (_10600_, _10599_, _10598_);
  nor (_10601_, _10600_, _10596_);
  nor (_10602_, _10601_, _02130_);
  or (_10603_, _10597_, _02131_);
  nor (_10604_, _10603_, _10543_);
  or (_10605_, _10604_, _02016_);
  nor (_10606_, _10605_, _10602_);
  nor (_10607_, _09111_, _06864_);
  nor (_10608_, _10607_, _10528_);
  and (_10609_, _10608_, _02016_);
  nor (_10610_, _10609_, _10606_);
  and (_10611_, _10610_, _05474_);
  nor (_10612_, _08974_, _06864_);
  nor (_10613_, _10612_, _10528_);
  nor (_10614_, _10613_, _05474_);
  or (_10615_, _10614_, _10611_);
  and (_10616_, _10615_, _02168_);
  nor (_10617_, _10540_, _02168_);
  or (_10618_, _10617_, _02025_);
  or (_10619_, _10618_, _10616_);
  nand (_10620_, _10561_, _02025_);
  and (_10621_, _10620_, _10619_);
  nor (_10622_, _10621_, _01594_);
  and (_10623_, _08965_, _04183_);
  nor (_10624_, _10623_, _10528_);
  and (_10625_, _10624_, _01594_);
  nor (_10626_, _10625_, _10622_);
  or (_10627_, _10626_, _26506_);
  or (_10628_, _26505_, \oc8051_golden_model_1.IE [6]);
  and (_10629_, _10628_, _25964_);
  and (_27765_, _10629_, _10627_);
  not (_10630_, \oc8051_golden_model_1.IP [0]);
  nor (_10631_, _04155_, _10630_);
  nor (_10632_, _04405_, _06757_);
  nor (_10633_, _10632_, _10631_);
  nor (_10634_, _10633_, _01595_);
  and (_10635_, _04155_, _05531_);
  nor (_10636_, _10635_, _10631_);
  nor (_10637_, _10636_, _05076_);
  not (_10638_, _10637_);
  nor (_10639_, _10638_, _10632_);
  and (_10640_, _04155_, _03677_);
  nor (_10641_, _10631_, _05513_);
  not (_10642_, _10641_);
  nor (_10643_, _10642_, _10640_);
  nor (_10644_, _05174_, _10630_);
  and (_10645_, _07725_, _05174_);
  nor (_10646_, _10645_, _10644_);
  nor (_10647_, _10646_, _02223_);
  and (_10648_, _10633_, _01969_);
  and (_10649_, _04155_, \oc8051_golden_model_1.ACC [0]);
  nor (_10650_, _10649_, _10631_);
  nor (_10651_, _10650_, _05488_);
  nor (_10652_, _04571_, _10630_);
  or (_10653_, _10652_, _01969_);
  nor (_10654_, _10653_, _10651_);
  or (_10655_, _10654_, _06233_);
  nor (_10656_, _10655_, _10648_);
  and (_10657_, _04155_, _03334_);
  nor (_10658_, _10657_, _10631_);
  nor (_10659_, _10658_, _05487_);
  or (_10660_, _10659_, _01963_);
  or (_10661_, _10660_, _10656_);
  nor (_10662_, _10661_, _10647_);
  and (_10663_, _10650_, _01963_);
  nor (_10664_, _10663_, _01957_);
  not (_10665_, _10664_);
  nor (_10666_, _10665_, _10662_);
  and (_10667_, _10631_, _01957_);
  or (_10668_, _10667_, _10666_);
  and (_10669_, _10668_, _04885_);
  nor (_10670_, _10633_, _04885_);
  or (_10671_, _10670_, _10669_);
  nor (_10672_, _10671_, _01924_);
  nor (_10673_, _07759_, _06794_);
  or (_10674_, _10644_, _01925_);
  nor (_10675_, _10674_, _10673_);
  or (_10676_, _10675_, _04950_);
  or (_10677_, _10676_, _10672_);
  or (_10678_, _10658_, _06397_);
  and (_10679_, _10678_, _05513_);
  and (_10680_, _10679_, _10677_);
  nor (_10681_, _10680_, _10643_);
  nor (_10682_, _10681_, _01602_);
  nor (_10683_, _07815_, _06757_);
  or (_10684_, _10631_, _01923_);
  nor (_10685_, _10684_, _10683_);
  or (_10686_, _10685_, _02019_);
  nor (_10687_, _10686_, _10682_);
  nand (_10688_, _10636_, _05049_);
  and (_10689_, _10688_, _06278_);
  nor (_10690_, _10689_, _10687_);
  and (_10691_, _07829_, _04155_);
  nor (_10692_, _10691_, _10631_);
  and (_10693_, _10692_, _02018_);
  nor (_10694_, _10693_, _10690_);
  and (_10695_, _10694_, _02136_);
  and (_10696_, _07834_, _04155_);
  nor (_10697_, _10696_, _10631_);
  nor (_10698_, _10697_, _02136_);
  or (_10699_, _10698_, _10695_);
  and (_10700_, _10699_, _05076_);
  nor (_10701_, _10700_, _10639_);
  nor (_10702_, _10701_, _02130_);
  nor (_10703_, _10631_, _04405_);
  or (_10704_, _10703_, _02131_);
  nor (_10705_, _10704_, _10650_);
  or (_10706_, _10705_, _02016_);
  nor (_10707_, _10706_, _10702_);
  nor (_10708_, _07828_, _06757_);
  nor (_10709_, _10708_, _10631_);
  and (_10710_, _10709_, _02016_);
  nor (_10711_, _10710_, _10707_);
  and (_10712_, _10711_, _05474_);
  nor (_10713_, _07696_, _06757_);
  nor (_10714_, _10713_, _10631_);
  nor (_10715_, _10714_, _05474_);
  or (_10716_, _10715_, _10712_);
  and (_10717_, _10716_, _02168_);
  nor (_10718_, _10633_, _02168_);
  nor (_10719_, _10718_, _02025_);
  not (_10720_, _10719_);
  nor (_10721_, _10720_, _10717_);
  nor (_10722_, _10631_, _02377_);
  nor (_10723_, _10722_, _10721_);
  and (_10724_, _10723_, _01595_);
  nor (_10725_, _10724_, _10634_);
  nand (_10726_, _10725_, _26505_);
  or (_10727_, _26505_, \oc8051_golden_model_1.IP [0]);
  and (_10728_, _10727_, _25964_);
  and (_27766_, _10728_, _10726_);
  nor (_10729_, _04155_, \oc8051_golden_model_1.IP [1]);
  not (_10730_, _10729_);
  nor (_10731_, _08029_, _06757_);
  nor (_10732_, _10731_, _02136_);
  and (_10733_, _10732_, _10730_);
  not (_10734_, \oc8051_golden_model_1.IP [1]);
  nor (_10735_, _04155_, _10734_);
  and (_10736_, _04155_, _03613_);
  or (_10737_, _10736_, _10735_);
  and (_10738_, _10737_, _04951_);
  nor (_10739_, _07953_, _06794_);
  nor (_10740_, _05174_, _10734_);
  or (_10741_, _10740_, _01925_);
  or (_10742_, _10741_, _10739_);
  and (_10743_, _07909_, _04155_);
  nor (_10744_, _10743_, _10729_);
  nor (_10745_, _10744_, _02438_);
  and (_10746_, _04155_, _01705_);
  nor (_10747_, _10746_, _10729_);
  and (_10748_, _10747_, _04571_);
  nor (_10749_, _04571_, _10734_);
  or (_10750_, _10749_, _01969_);
  nor (_10751_, _10750_, _10748_);
  or (_10752_, _10751_, _06233_);
  nor (_10753_, _10752_, _10745_);
  nor (_10754_, _06757_, _03393_);
  nor (_10755_, _10754_, _10735_);
  nor (_10756_, _10755_, _05487_);
  and (_10757_, _07920_, _05174_);
  nor (_10758_, _10757_, _10740_);
  nor (_10759_, _10758_, _02223_);
  nor (_10760_, _10759_, _10756_);
  nand (_10761_, _10760_, _01964_);
  or (_10762_, _10761_, _10753_);
  or (_10763_, _10747_, _01964_);
  and (_10764_, _10763_, _10762_);
  and (_10765_, _10764_, _06229_);
  and (_10766_, _07907_, _05174_);
  nor (_10767_, _10766_, _10740_);
  nor (_10768_, _10767_, _06229_);
  or (_10769_, _10768_, _10765_);
  and (_10770_, _10769_, _04885_);
  nor (_10771_, _10740_, _07935_);
  or (_10772_, _10771_, _04885_);
  nor (_10773_, _10772_, _10758_);
  or (_10774_, _10773_, _01924_);
  or (_10775_, _10774_, _10770_);
  and (_10776_, _10775_, _10742_);
  nor (_10777_, _10776_, _04950_);
  and (_10778_, _10755_, _04950_);
  or (_10779_, _10778_, _04951_);
  nor (_10780_, _10779_, _10777_);
  or (_10781_, _10780_, _10738_);
  and (_10782_, _10781_, _01923_);
  nor (_10783_, _08009_, _06757_);
  nor (_10784_, _10783_, _10735_);
  nor (_10785_, _10784_, _01923_);
  nor (_10786_, _10785_, _10782_);
  nor (_10787_, _10786_, _06278_);
  nor (_10788_, _08023_, _06757_);
  nor (_10789_, _10788_, _05049_);
  and (_10790_, _04155_, _02676_);
  nor (_10791_, _10790_, _04979_);
  or (_10792_, _10791_, _10789_);
  and (_10793_, _10792_, _10730_);
  nor (_10794_, _10793_, _10787_);
  nor (_10795_, _10794_, _02135_);
  nor (_10796_, _10795_, _10733_);
  nor (_10797_, _10796_, _02039_);
  nor (_10798_, _07893_, _06757_);
  nor (_10799_, _10798_, _05076_);
  and (_10800_, _10799_, _10730_);
  nor (_10801_, _10800_, _10797_);
  nor (_10802_, _10801_, _02130_);
  nor (_10803_, _10735_, _05741_);
  nor (_10804_, _10803_, _02131_);
  and (_10805_, _10804_, _10747_);
  nor (_10806_, _10805_, _10802_);
  nor (_10807_, _10806_, _02128_);
  and (_10808_, _10790_, _04452_);
  nor (_10809_, _10808_, _05104_);
  nand (_10810_, _10746_, _04452_);
  and (_10811_, _10810_, _02126_);
  or (_10812_, _10811_, _10809_);
  and (_10813_, _10812_, _10730_);
  or (_10814_, _10813_, _02164_);
  nor (_10815_, _10814_, _10807_);
  nor (_10816_, _10744_, _02168_);
  or (_10817_, _10816_, _02025_);
  nor (_10818_, _10817_, _10815_);
  nor (_10819_, _10767_, _02377_);
  or (_10820_, _10819_, _01594_);
  nor (_10821_, _10820_, _10818_);
  nor (_10822_, _10743_, _10735_);
  and (_10823_, _10822_, _01594_);
  nor (_10824_, _10823_, _10821_);
  or (_10825_, _10824_, _26506_);
  or (_10826_, _26505_, \oc8051_golden_model_1.IP [1]);
  and (_10827_, _10826_, _25964_);
  and (_27769_, _10827_, _10825_);
  not (_10828_, \oc8051_golden_model_1.IP [2]);
  nor (_10829_, _04155_, _10828_);
  and (_10830_, _04155_, _05563_);
  nor (_10831_, _10830_, _10829_);
  and (_10832_, _10831_, _02019_);
  nor (_10833_, _06757_, _03272_);
  nor (_10834_, _10833_, _10829_);
  and (_10835_, _10834_, _04950_);
  nor (_10836_, _08095_, _06757_);
  nor (_10837_, _10836_, _10829_);
  and (_10838_, _10837_, _01969_);
  and (_10839_, _04155_, \oc8051_golden_model_1.ACC [2]);
  nor (_10840_, _10839_, _10829_);
  nor (_10841_, _10840_, _05488_);
  nor (_10842_, _04571_, _10828_);
  or (_10843_, _10842_, _01969_);
  nor (_10844_, _10843_, _10841_);
  or (_10845_, _10844_, _06233_);
  nor (_10846_, _10845_, _10838_);
  nor (_10847_, _10834_, _05487_);
  nor (_10848_, _05174_, _10828_);
  and (_10849_, _08111_, _05174_);
  nor (_10850_, _10849_, _10848_);
  nor (_10851_, _10850_, _02223_);
  nor (_10852_, _10851_, _10847_);
  nand (_10853_, _10852_, _01964_);
  or (_10854_, _10853_, _10846_);
  nand (_10855_, _10840_, _01963_);
  and (_10856_, _10855_, _10854_);
  nor (_10857_, _10856_, _01957_);
  and (_10858_, _08109_, _05174_);
  nor (_10859_, _10858_, _10848_);
  and (_10860_, _10859_, _01957_);
  or (_10861_, _10860_, _01946_);
  nor (_10862_, _10861_, _10857_);
  nor (_10863_, _10848_, _08139_);
  or (_10864_, _10863_, _04885_);
  nor (_10865_, _10864_, _10850_);
  or (_10866_, _10865_, _10862_);
  and (_10867_, _10866_, _01925_);
  nor (_10868_, _08158_, _06794_);
  nor (_10869_, _10848_, _10868_);
  nor (_10870_, _10869_, _01925_);
  or (_10871_, _10870_, _04950_);
  nor (_10872_, _10871_, _10867_);
  nor (_10873_, _10872_, _10835_);
  nor (_10874_, _10873_, _04951_);
  and (_10875_, _04155_, _03564_);
  nor (_10876_, _10829_, _05513_);
  not (_10877_, _10876_);
  nor (_10878_, _10877_, _10875_);
  or (_10879_, _10878_, _01602_);
  nor (_10880_, _10879_, _10874_);
  nor (_10881_, _08216_, _06757_);
  nor (_10882_, _10881_, _10829_);
  nor (_10883_, _10882_, _01923_);
  or (_10884_, _10883_, _02019_);
  nor (_10885_, _10884_, _10880_);
  nor (_10886_, _10885_, _10832_);
  or (_10887_, _10886_, _02018_);
  and (_10888_, _08230_, _04155_);
  or (_10889_, _10888_, _10829_);
  or (_10890_, _10889_, _05049_);
  and (_10891_, _10890_, _02136_);
  and (_10892_, _10891_, _10887_);
  and (_10893_, _08237_, _04155_);
  nor (_10894_, _10893_, _10829_);
  nor (_10895_, _10894_, _02136_);
  nor (_10896_, _10895_, _10892_);
  nor (_10897_, _10896_, _02039_);
  nor (_10898_, _10829_, _05739_);
  not (_10899_, _10898_);
  nor (_10900_, _10831_, _05076_);
  and (_10901_, _10900_, _10899_);
  nor (_10902_, _10901_, _10897_);
  nor (_10903_, _10902_, _02130_);
  or (_10904_, _10898_, _02131_);
  nor (_10905_, _10904_, _10840_);
  or (_10906_, _10905_, _02016_);
  nor (_10907_, _10906_, _10903_);
  nor (_10908_, _08229_, _06757_);
  nor (_10909_, _10908_, _10829_);
  and (_10910_, _10909_, _02016_);
  nor (_10911_, _10910_, _10907_);
  and (_10912_, _10911_, _05474_);
  nor (_10913_, _08236_, _06757_);
  nor (_10914_, _10913_, _10829_);
  nor (_10915_, _10914_, _05474_);
  or (_10916_, _10915_, _10912_);
  and (_10917_, _10916_, _02168_);
  nor (_10918_, _10837_, _02168_);
  or (_10919_, _10918_, _02025_);
  or (_10920_, _10919_, _10917_);
  nand (_10921_, _10859_, _02025_);
  and (_10922_, _10921_, _10920_);
  nor (_10923_, _10922_, _01594_);
  and (_10924_, _08285_, _04155_);
  nor (_10925_, _10924_, _10829_);
  and (_10926_, _10925_, _01594_);
  nor (_10927_, _10926_, _10923_);
  or (_10928_, _10927_, _26506_);
  or (_10929_, _26505_, \oc8051_golden_model_1.IP [2]);
  and (_10930_, _10929_, _25964_);
  and (_27770_, _10930_, _10928_);
  not (_10931_, \oc8051_golden_model_1.IP [3]);
  nor (_10932_, _04155_, _10931_);
  and (_10933_, _04155_, _05529_);
  nor (_10934_, _10933_, _10932_);
  and (_10935_, _10934_, _02019_);
  nor (_10936_, _06757_, _03473_);
  nor (_10937_, _10936_, _10932_);
  and (_10938_, _10937_, _04950_);
  nor (_10939_, _08308_, _06794_);
  nor (_10940_, _05174_, _10931_);
  or (_10941_, _10940_, _01925_);
  or (_10942_, _10941_, _10939_);
  nor (_10943_, _08337_, _06757_);
  nor (_10944_, _10943_, _10932_);
  and (_10945_, _10944_, _01969_);
  and (_10946_, _04155_, \oc8051_golden_model_1.ACC [3]);
  nor (_10947_, _10946_, _10932_);
  nor (_10948_, _10947_, _05488_);
  nor (_10949_, _04571_, _10931_);
  or (_10950_, _10949_, _01969_);
  nor (_10951_, _10950_, _10948_);
  or (_10952_, _10951_, _06233_);
  nor (_10953_, _10952_, _10945_);
  nor (_10954_, _10937_, _05487_);
  and (_10955_, _08341_, _05174_);
  nor (_10956_, _10955_, _10940_);
  nor (_10957_, _10956_, _02223_);
  nor (_10958_, _10957_, _10954_);
  nand (_10959_, _10958_, _01964_);
  or (_10960_, _10959_, _10953_);
  nand (_10961_, _10947_, _01963_);
  and (_10962_, _10961_, _10960_);
  and (_10963_, _10962_, _06229_);
  and (_10964_, _08324_, _05174_);
  nor (_10965_, _10964_, _10940_);
  nor (_10966_, _10965_, _06229_);
  or (_10967_, _10966_, _10963_);
  and (_10968_, _10967_, _04885_);
  nor (_10969_, _10940_, _08357_);
  or (_10970_, _10956_, _04885_);
  nor (_10971_, _10970_, _10969_);
  or (_10972_, _10971_, _01924_);
  or (_10973_, _10972_, _10968_);
  and (_10974_, _10973_, _10942_);
  nor (_10975_, _10974_, _04950_);
  nor (_10976_, _10975_, _10938_);
  nor (_10977_, _10976_, _04951_);
  and (_10978_, _04155_, _03516_);
  nor (_10979_, _10932_, _05513_);
  not (_10980_, _10979_);
  nor (_10981_, _10980_, _10978_);
  or (_10982_, _10981_, _01602_);
  nor (_10983_, _10982_, _10977_);
  nor (_10984_, _08425_, _06757_);
  nor (_10985_, _10984_, _10932_);
  nor (_10986_, _10985_, _01923_);
  or (_10987_, _10986_, _02019_);
  nor (_10988_, _10987_, _10983_);
  nor (_10989_, _10988_, _10935_);
  or (_10990_, _10989_, _02018_);
  and (_10991_, _08441_, _04155_);
  or (_10992_, _10991_, _10932_);
  or (_10993_, _10992_, _05049_);
  and (_10994_, _10993_, _02136_);
  and (_10995_, _10994_, _10990_);
  and (_10996_, _08304_, _04155_);
  nor (_10997_, _10996_, _10932_);
  nor (_10998_, _10997_, _02136_);
  nor (_10999_, _10998_, _10995_);
  nor (_11000_, _10999_, _02039_);
  nor (_11001_, _10932_, _05737_);
  not (_11002_, _11001_);
  nor (_11003_, _10934_, _05076_);
  and (_11004_, _11003_, _11002_);
  nor (_11005_, _11004_, _11000_);
  nor (_11006_, _11005_, _02130_);
  or (_11007_, _11001_, _02131_);
  nor (_11008_, _11007_, _10947_);
  or (_11009_, _11008_, _02016_);
  nor (_11010_, _11009_, _11006_);
  nor (_11011_, _08440_, _06757_);
  nor (_11012_, _11011_, _10932_);
  and (_11013_, _11012_, _02016_);
  nor (_11014_, _11013_, _11010_);
  and (_11015_, _11014_, _05474_);
  nor (_11016_, _08303_, _06757_);
  nor (_11017_, _11016_, _10932_);
  nor (_11018_, _11017_, _05474_);
  or (_11019_, _11018_, _11015_);
  and (_11020_, _11019_, _02168_);
  nor (_11021_, _10944_, _02168_);
  or (_11022_, _11021_, _02025_);
  or (_11023_, _11022_, _11020_);
  nand (_11024_, _10965_, _02025_);
  and (_11025_, _11024_, _11023_);
  nor (_11026_, _11025_, _01594_);
  and (_11027_, _08507_, _04155_);
  nor (_11028_, _11027_, _10932_);
  and (_11029_, _11028_, _01594_);
  nor (_11030_, _11029_, _11026_);
  or (_11031_, _11030_, _26506_);
  or (_11032_, _26505_, \oc8051_golden_model_1.IP [3]);
  and (_11033_, _11032_, _25964_);
  and (_27771_, _11033_, _11031_);
  not (_11034_, \oc8051_golden_model_1.IP [4]);
  nor (_11035_, _04155_, _11034_);
  and (_11036_, _04155_, _05524_);
  nor (_11037_, _11036_, _11035_);
  and (_11038_, _11037_, _02019_);
  nor (_11039_, _06757_, _04024_);
  nor (_11040_, _11039_, _11035_);
  and (_11041_, _11040_, _04950_);
  nor (_11042_, _08548_, _06757_);
  nor (_11043_, _11042_, _11035_);
  and (_11044_, _11043_, _01969_);
  and (_11045_, _04155_, \oc8051_golden_model_1.ACC [4]);
  nor (_11046_, _11045_, _11035_);
  nor (_11047_, _11046_, _05488_);
  nor (_11048_, _04571_, _11034_);
  or (_11049_, _11048_, _01969_);
  nor (_11050_, _11049_, _11047_);
  or (_11051_, _11050_, _06233_);
  nor (_11052_, _11051_, _11044_);
  nor (_11053_, _11040_, _05487_);
  nor (_11054_, _05174_, _11034_);
  and (_11055_, _08565_, _05174_);
  nor (_11056_, _11055_, _11054_);
  nor (_11057_, _11056_, _02223_);
  nor (_11058_, _11057_, _11053_);
  nand (_11059_, _11058_, _01964_);
  or (_11060_, _11059_, _11052_);
  nand (_11061_, _11046_, _01963_);
  and (_11062_, _11061_, _11060_);
  and (_11063_, _11062_, _06229_);
  and (_11064_, _08544_, _05174_);
  nor (_11065_, _11064_, _11054_);
  nor (_11066_, _11065_, _06229_);
  or (_11067_, _11066_, _11063_);
  and (_11068_, _11067_, _04885_);
  and (_11069_, _08582_, _05174_);
  nor (_11070_, _11069_, _11054_);
  nor (_11071_, _11070_, _04885_);
  nor (_11072_, _11071_, _11068_);
  nor (_11073_, _11072_, _01924_);
  nor (_11074_, _08607_, _06794_);
  nor (_11075_, _11074_, _11054_);
  nor (_11076_, _11075_, _01925_);
  nor (_11077_, _11076_, _04950_);
  not (_11078_, _11077_);
  nor (_11079_, _11078_, _11073_);
  nor (_11080_, _11079_, _11041_);
  nor (_11081_, _11080_, _04951_);
  and (_11082_, _04155_, _03903_);
  nor (_11083_, _11035_, _05513_);
  not (_11084_, _11083_);
  nor (_11085_, _11084_, _11082_);
  or (_11086_, _11085_, _01602_);
  nor (_11087_, _11086_, _11081_);
  nor (_11088_, _08663_, _06757_);
  nor (_11089_, _11088_, _11035_);
  nor (_11090_, _11089_, _01923_);
  or (_11091_, _11090_, _02019_);
  nor (_11092_, _11091_, _11087_);
  nor (_11093_, _11092_, _11038_);
  or (_11094_, _11093_, _02018_);
  and (_11095_, _08531_, _04155_);
  or (_11096_, _11095_, _11035_);
  or (_11097_, _11096_, _05049_);
  and (_11098_, _11097_, _02136_);
  and (_11099_, _11098_, _11094_);
  and (_11100_, _08527_, _04155_);
  nor (_11101_, _11100_, _11035_);
  nor (_11102_, _11101_, _02136_);
  nor (_11103_, _11102_, _11099_);
  nor (_11104_, _11103_, _02039_);
  nor (_11105_, _11035_, _08729_);
  not (_11106_, _11105_);
  nor (_11107_, _11037_, _05076_);
  and (_11108_, _11107_, _11106_);
  nor (_11109_, _11108_, _11104_);
  nor (_11110_, _11109_, _02130_);
  or (_11111_, _11105_, _02131_);
  nor (_11112_, _11111_, _11046_);
  or (_11113_, _11112_, _02016_);
  nor (_11114_, _11113_, _11110_);
  nor (_11115_, _08530_, _06757_);
  nor (_11116_, _11115_, _11035_);
  and (_11117_, _11116_, _02016_);
  nor (_11118_, _11117_, _11114_);
  and (_11119_, _11118_, _05474_);
  nor (_11120_, _08526_, _06757_);
  nor (_11121_, _11120_, _11035_);
  nor (_11122_, _11121_, _05474_);
  or (_11123_, _11122_, _11119_);
  and (_11124_, _11123_, _02168_);
  nor (_11125_, _11043_, _02168_);
  or (_11126_, _11125_, _02025_);
  or (_11127_, _11126_, _11124_);
  nand (_11128_, _11065_, _02025_);
  and (_11129_, _11128_, _11127_);
  nor (_11130_, _11129_, _01594_);
  and (_11131_, _08732_, _04155_);
  nor (_11132_, _11131_, _11035_);
  and (_11133_, _11132_, _01594_);
  nor (_11134_, _11133_, _11130_);
  or (_11135_, _11134_, _26506_);
  or (_11136_, _26505_, \oc8051_golden_model_1.IP [4]);
  and (_11137_, _11136_, _25964_);
  and (_27772_, _11137_, _11135_);
  not (_11138_, \oc8051_golden_model_1.IP [5]);
  nor (_11139_, _04155_, _11138_);
  and (_11140_, _04155_, _05548_);
  nor (_11141_, _11140_, _11139_);
  and (_11142_, _11141_, _02019_);
  nor (_11143_, _06757_, _03976_);
  nor (_11144_, _11143_, _11139_);
  and (_11145_, _11144_, _04950_);
  nor (_11146_, _05174_, _11138_);
  nor (_11147_, _11146_, _08801_);
  and (_11148_, _08785_, _05174_);
  nor (_11149_, _11148_, _11146_);
  or (_11150_, _11149_, _04885_);
  nor (_11151_, _11150_, _11147_);
  nor (_11152_, _08771_, _06757_);
  nor (_11153_, _11152_, _11139_);
  and (_11154_, _11153_, _01969_);
  and (_11155_, _04155_, \oc8051_golden_model_1.ACC [5]);
  nor (_11156_, _11155_, _11139_);
  nor (_11157_, _11156_, _05488_);
  nor (_11158_, _04571_, _11138_);
  or (_11159_, _11158_, _01969_);
  nor (_11160_, _11159_, _11157_);
  or (_11161_, _11160_, _06233_);
  nor (_11162_, _11161_, _11154_);
  nor (_11163_, _11144_, _05487_);
  nor (_11164_, _11149_, _02223_);
  nor (_11165_, _11164_, _11163_);
  nand (_11166_, _11165_, _01964_);
  or (_11167_, _11166_, _11162_);
  nand (_11168_, _11156_, _01963_);
  and (_11169_, _11168_, _11167_);
  and (_11170_, _11169_, _06229_);
  and (_11171_, _08768_, _05174_);
  nor (_11172_, _11171_, _11146_);
  nor (_11173_, _11172_, _06229_);
  or (_11174_, _11173_, _11170_);
  and (_11175_, _11174_, _04885_);
  nor (_11176_, _11175_, _11151_);
  nor (_11177_, _11176_, _01924_);
  nor (_11178_, _08754_, _06794_);
  nor (_11179_, _11178_, _11146_);
  nor (_11180_, _11179_, _01925_);
  nor (_11181_, _11180_, _04950_);
  not (_11182_, _11181_);
  nor (_11183_, _11182_, _11177_);
  nor (_11184_, _11183_, _11145_);
  nor (_11185_, _11184_, _04951_);
  and (_11186_, _04155_, _03850_);
  nor (_11187_, _11139_, _05513_);
  not (_11188_, _11187_);
  nor (_11189_, _11188_, _11186_);
  or (_11190_, _11189_, _01602_);
  nor (_11191_, _11190_, _11185_);
  nor (_11192_, _08874_, _06757_);
  nor (_11193_, _11192_, _11139_);
  nor (_11194_, _11193_, _01923_);
  or (_11195_, _11194_, _02019_);
  nor (_11196_, _11195_, _11191_);
  nor (_11197_, _11196_, _11142_);
  or (_11198_, _11197_, _02018_);
  and (_11199_, _08890_, _04155_);
  or (_11200_, _11199_, _11139_);
  or (_11201_, _11200_, _05049_);
  and (_11202_, _11201_, _02136_);
  and (_11203_, _11202_, _11198_);
  and (_11204_, _08750_, _04155_);
  nor (_11205_, _11204_, _11139_);
  nor (_11206_, _11205_, _02136_);
  nor (_11207_, _11206_, _11203_);
  nor (_11208_, _11207_, _02039_);
  nor (_11209_, _11139_, _08946_);
  not (_11210_, _11209_);
  nor (_11211_, _11141_, _05076_);
  and (_11212_, _11211_, _11210_);
  nor (_11213_, _11212_, _11208_);
  nor (_11214_, _11213_, _02130_);
  or (_11215_, _11209_, _02131_);
  nor (_11216_, _11215_, _11156_);
  or (_11217_, _11216_, _02016_);
  nor (_11218_, _11217_, _11214_);
  nor (_11219_, _08889_, _06757_);
  nor (_11220_, _11219_, _11139_);
  and (_11221_, _11220_, _02016_);
  nor (_11222_, _11221_, _11218_);
  and (_11223_, _11222_, _05474_);
  nor (_11224_, _08749_, _06757_);
  nor (_11225_, _11224_, _11139_);
  nor (_11226_, _11225_, _05474_);
  or (_11227_, _11226_, _11223_);
  and (_11228_, _11227_, _02168_);
  nor (_11229_, _11153_, _02168_);
  or (_11230_, _11229_, _02025_);
  or (_11231_, _11230_, _11228_);
  nand (_11232_, _11172_, _02025_);
  and (_11233_, _11232_, _11231_);
  nor (_11234_, _11233_, _01594_);
  and (_11235_, _08949_, _04155_);
  nor (_11236_, _11235_, _11139_);
  and (_11237_, _11236_, _01594_);
  nor (_11238_, _11237_, _11234_);
  or (_11239_, _11238_, _26506_);
  or (_11240_, _26505_, \oc8051_golden_model_1.IP [5]);
  and (_11241_, _11240_, _25964_);
  and (_27773_, _11241_, _11239_);
  not (_11242_, \oc8051_golden_model_1.IP [6]);
  nor (_11243_, _04155_, _11242_);
  and (_11244_, _04155_, _03748_);
  or (_11245_, _11244_, _11243_);
  and (_11246_, _11245_, _04951_);
  nor (_11247_, _05174_, _11242_);
  not (_11248_, _11247_);
  and (_11249_, _11248_, _09026_);
  and (_11250_, _09011_, _05174_);
  nor (_11251_, _11250_, _11247_);
  or (_11252_, _11251_, _04885_);
  nor (_11253_, _11252_, _11249_);
  nor (_11254_, _08995_, _06757_);
  nor (_11255_, _11254_, _11243_);
  and (_11256_, _11255_, _01969_);
  and (_11257_, _04155_, \oc8051_golden_model_1.ACC [6]);
  nor (_11258_, _11257_, _11243_);
  nor (_11259_, _11258_, _05488_);
  nor (_11260_, _04571_, _11242_);
  or (_11261_, _11260_, _01969_);
  nor (_11262_, _11261_, _11259_);
  or (_11263_, _11262_, _06233_);
  nor (_11264_, _11263_, _11256_);
  nor (_11265_, _06757_, _04074_);
  nor (_11266_, _11265_, _11243_);
  nor (_11267_, _11266_, _05487_);
  nor (_11268_, _11251_, _02223_);
  nor (_11269_, _11268_, _11267_);
  nand (_11270_, _11269_, _01964_);
  or (_11271_, _11270_, _11264_);
  nand (_11272_, _11258_, _01963_);
  and (_11273_, _11272_, _11271_);
  and (_11274_, _11273_, _06229_);
  and (_11275_, _08992_, _05174_);
  nor (_11276_, _11275_, _11247_);
  nor (_11277_, _11276_, _06229_);
  or (_11278_, _11277_, _11274_);
  and (_11279_, _11278_, _04885_);
  nor (_11280_, _11279_, _11253_);
  nor (_11281_, _11280_, _01924_);
  nor (_11282_, _08979_, _06794_);
  nor (_11283_, _11282_, _11247_);
  nor (_11284_, _11283_, _01925_);
  nor (_11285_, _11284_, _04950_);
  not (_11286_, _11285_);
  nor (_11287_, _11286_, _11281_);
  and (_11288_, _11266_, _04950_);
  or (_11289_, _11288_, _04951_);
  nor (_11290_, _11289_, _11287_);
  or (_11291_, _11290_, _11246_);
  and (_11292_, _11291_, _01923_);
  nor (_11293_, _09096_, _06757_);
  nor (_11294_, _11293_, _11243_);
  nor (_11295_, _11294_, _01923_);
  or (_11296_, _11295_, _06278_);
  or (_11297_, _11296_, _11292_);
  and (_11298_, _09112_, _04155_);
  or (_11299_, _11243_, _05049_);
  or (_11300_, _11299_, _11298_);
  and (_11301_, _04155_, _09103_);
  nor (_11302_, _11301_, _11243_);
  and (_11303_, _11302_, _02019_);
  nor (_11304_, _11303_, _02135_);
  and (_11305_, _11304_, _11300_);
  and (_11306_, _11305_, _11297_);
  and (_11307_, _08975_, _04155_);
  nor (_11308_, _11307_, _11243_);
  nor (_11309_, _11308_, _02136_);
  nor (_11310_, _11309_, _11306_);
  nor (_11311_, _11310_, _02039_);
  nor (_11312_, _11243_, _05735_);
  not (_11313_, _11312_);
  nor (_11314_, _11302_, _05076_);
  and (_11315_, _11314_, _11313_);
  nor (_11316_, _11315_, _11311_);
  nor (_11317_, _11316_, _02130_);
  or (_11318_, _11312_, _02131_);
  nor (_11319_, _11318_, _11258_);
  or (_11320_, _11319_, _02016_);
  nor (_11321_, _11320_, _11317_);
  nor (_11322_, _09111_, _06757_);
  nor (_11323_, _11322_, _11243_);
  and (_11324_, _11323_, _02016_);
  nor (_11325_, _11324_, _11321_);
  and (_11326_, _11325_, _05474_);
  nor (_11327_, _08974_, _06757_);
  nor (_11328_, _11327_, _11243_);
  nor (_11329_, _11328_, _05474_);
  or (_11330_, _11329_, _11326_);
  and (_11331_, _11330_, _02168_);
  nor (_11332_, _11255_, _02168_);
  or (_11333_, _11332_, _02025_);
  or (_11334_, _11333_, _11331_);
  nand (_11335_, _11276_, _02025_);
  and (_11336_, _11335_, _11334_);
  nor (_11337_, _11336_, _01594_);
  and (_11338_, _08965_, _04155_);
  nor (_11339_, _11338_, _11243_);
  and (_11340_, _11339_, _01594_);
  nor (_11341_, _11340_, _11337_);
  or (_11342_, _11341_, _26506_);
  or (_11343_, _26505_, \oc8051_golden_model_1.IP [6]);
  and (_11344_, _11343_, _25964_);
  and (_27774_, _11344_, _11342_);
  nor (_11345_, \oc8051_golden_model_1.P0 [0], rst);
  nor (_27777_, _11345_, _06750_);
  nor (_11346_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_27778_, _11346_, _06750_);
  nor (_11347_, \oc8051_golden_model_1.P0 [2], rst);
  nor (_27779_, _11347_, _06750_);
  nor (_11348_, \oc8051_golden_model_1.P0 [3], rst);
  nor (_27780_, _11348_, _06750_);
  nor (_11349_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_27781_, _11349_, _06750_);
  nor (_11350_, \oc8051_golden_model_1.P0 [5], rst);
  nor (_27782_, _11350_, _06750_);
  nor (_11351_, \oc8051_golden_model_1.P0 [6], rst);
  nor (_27783_, _11351_, _06750_);
  nor (_11352_, \oc8051_golden_model_1.P1 [0], rst);
  nor (_27786_, _11352_, _06750_);
  nor (_11353_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_27787_, _11353_, _06750_);
  nor (_11354_, \oc8051_golden_model_1.P1 [2], rst);
  nor (_27788_, _11354_, _06750_);
  nor (_11355_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_27789_, _11355_, _06750_);
  nor (_11356_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_27790_, _11356_, _06750_);
  nor (_11357_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_27791_, _11357_, _06750_);
  nor (_11358_, \oc8051_golden_model_1.P1 [6], rst);
  nor (_27792_, _11358_, _06750_);
  nor (_11359_, \oc8051_golden_model_1.P2 [0], rst);
  nor (_27797_, _11359_, _06750_);
  nor (_11360_, \oc8051_golden_model_1.P2 [1], rst);
  nor (_27798_, _11360_, _06750_);
  nor (_11361_, \oc8051_golden_model_1.P2 [2], rst);
  nor (_27799_, _11361_, _06750_);
  nor (_11362_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_27800_, _11362_, _06750_);
  nor (_11363_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_27801_, _11363_, _06750_);
  nor (_11364_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_27802_, _11364_, _06750_);
  nor (_11365_, \oc8051_golden_model_1.P2 [6], rst);
  nor (_27803_, _11365_, _06750_);
  nor (_11366_, \oc8051_golden_model_1.P3 [0], rst);
  nor (_27806_, _11366_, _06750_);
  nor (_11367_, \oc8051_golden_model_1.P3 [1], rst);
  nor (_27807_, _11367_, _06750_);
  nor (_11368_, \oc8051_golden_model_1.P3 [2], rst);
  nor (_27808_, _11368_, _06750_);
  nor (_11369_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_27809_, _11369_, _06750_);
  nor (_11370_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_27810_, _11370_, _06750_);
  nor (_11371_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_27811_, _11371_, _06750_);
  nor (_11372_, \oc8051_golden_model_1.P3 [6], rst);
  nor (_27812_, _11372_, _06750_);
  nand (_11373_, \oc8051_golden_model_1.PSW [0], _25964_);
  nor (_27815_, _11373_, _26505_);
  nand (_11374_, \oc8051_golden_model_1.PSW [1], _25964_);
  nor (_27816_, _11374_, _26505_);
  nand (_11375_, \oc8051_golden_model_1.PSW [2], _25964_);
  nor (_27817_, _11375_, _26505_);
  or (_11376_, _01974_, rst);
  nor (_27818_, _11376_, _26505_);
  nand (_11377_, \oc8051_golden_model_1.PSW [4], _25964_);
  nor (_27819_, _11377_, _26505_);
  nand (_11378_, \oc8051_golden_model_1.PSW [5], _25964_);
  nor (_27820_, _11378_, _26505_);
  nand (_11379_, \oc8051_golden_model_1.PSW [6], _25964_);
  nor (_27823_, _11379_, _26505_);
  not (_11380_, \oc8051_golden_model_1.PCON [0]);
  nor (_11381_, _04177_, _11380_);
  nor (_11382_, _04405_, _06680_);
  nor (_11383_, _11382_, _11381_);
  and (_11384_, _11383_, _02266_);
  and (_11385_, _04177_, _05531_);
  nor (_11386_, _11385_, _11381_);
  nor (_11387_, _11386_, _05076_);
  not (_11388_, _11387_);
  nor (_11389_, _11388_, _11382_);
  and (_11390_, _04177_, \oc8051_golden_model_1.ACC [0]);
  nor (_11391_, _11390_, _11381_);
  nor (_11392_, _11391_, _01964_);
  nor (_11393_, _11391_, _05488_);
  nor (_11394_, _04571_, _11380_);
  or (_11395_, _11394_, _11393_);
  and (_11396_, _11395_, _02438_);
  nor (_11397_, _11383_, _02438_);
  or (_11398_, _11397_, _11396_);
  and (_11399_, _11398_, _05487_);
  and (_11400_, _04177_, _03334_);
  nor (_11401_, _11400_, _11381_);
  nor (_11402_, _11401_, _05487_);
  nor (_11403_, _11402_, _11399_);
  nor (_11404_, _11403_, _01963_);
  or (_11405_, _11404_, _04950_);
  nor (_11406_, _11405_, _11392_);
  and (_11407_, _11401_, _04950_);
  nor (_11408_, _11407_, _11406_);
  nor (_11409_, _11408_, _04951_);
  and (_11410_, _04177_, _03677_);
  nor (_11411_, _11381_, _05513_);
  not (_11412_, _11411_);
  nor (_11413_, _11412_, _11410_);
  nor (_11414_, _11413_, _11409_);
  nor (_11415_, _11414_, _01602_);
  nor (_11416_, _07815_, _06680_);
  or (_11417_, _11381_, _01923_);
  nor (_11418_, _11417_, _11416_);
  or (_11419_, _11418_, _02019_);
  nor (_11420_, _11419_, _11415_);
  nand (_11421_, _11386_, _05049_);
  and (_11422_, _11421_, _06278_);
  nor (_11423_, _11422_, _11420_);
  and (_11424_, _07829_, _04177_);
  nor (_11425_, _11424_, _11381_);
  and (_11426_, _11425_, _02018_);
  nor (_11427_, _11426_, _11423_);
  and (_11428_, _11427_, _02136_);
  and (_11429_, _07834_, _04177_);
  nor (_11430_, _11429_, _11381_);
  nor (_11431_, _11430_, _02136_);
  or (_11432_, _11431_, _11428_);
  and (_11433_, _11432_, _05076_);
  nor (_11434_, _11433_, _11389_);
  nor (_11435_, _11434_, _02130_);
  and (_11436_, _07833_, _04177_);
  or (_11437_, _11436_, _11381_);
  and (_11438_, _11437_, _02130_);
  or (_11439_, _11438_, _11435_);
  and (_11440_, _11439_, _05104_);
  nor (_11441_, _07828_, _06680_);
  nor (_11442_, _11441_, _11381_);
  nor (_11443_, _11442_, _05104_);
  or (_11444_, _11443_, _11440_);
  and (_11445_, _11444_, _05474_);
  nor (_11446_, _07696_, _06680_);
  nor (_11447_, _11446_, _11381_);
  nor (_11448_, _11447_, _05474_);
  nor (_11449_, _11448_, _02266_);
  not (_11450_, _11449_);
  nor (_11451_, _11450_, _11445_);
  nor (_11452_, _11451_, _11384_);
  or (_11453_, _11452_, _26506_);
  or (_11454_, _26505_, \oc8051_golden_model_1.PCON [0]);
  and (_11455_, _11454_, _25964_);
  and (_27824_, _11455_, _11453_);
  nor (_11456_, _04177_, \oc8051_golden_model_1.PCON [1]);
  and (_11457_, _07909_, _04177_);
  nor (_11458_, _11457_, _11456_);
  nor (_11459_, _11458_, _02168_);
  not (_11460_, _11456_);
  nor (_11461_, _07893_, _06680_);
  nor (_11462_, _11461_, _05076_);
  and (_11463_, _11462_, _11460_);
  nor (_11464_, _08029_, _06680_);
  nor (_11465_, _11464_, _02136_);
  and (_11466_, _11465_, _11460_);
  and (_11467_, _04177_, _03613_);
  not (_11468_, \oc8051_golden_model_1.PCON [1]);
  nor (_11469_, _04177_, _11468_);
  nor (_11470_, _11469_, _05513_);
  not (_11471_, _11470_);
  nor (_11472_, _11471_, _11467_);
  not (_11473_, _11472_);
  nor (_11474_, _06680_, _03393_);
  nor (_11475_, _11474_, _11469_);
  and (_11476_, _11475_, _04950_);
  and (_11477_, _04177_, _01705_);
  nor (_11478_, _11477_, _11456_);
  and (_11479_, _11478_, _01963_);
  and (_11480_, _11478_, _04571_);
  nor (_11481_, _04571_, _11468_);
  or (_11482_, _11481_, _11480_);
  and (_11483_, _11482_, _02438_);
  and (_11484_, _11458_, _01969_);
  or (_11485_, _11484_, _11483_);
  and (_11486_, _11485_, _05487_);
  nor (_11487_, _11475_, _05487_);
  nor (_11488_, _11487_, _11486_);
  nor (_11489_, _11488_, _01963_);
  or (_11490_, _11489_, _04950_);
  nor (_11491_, _11490_, _11479_);
  nor (_11492_, _11491_, _11476_);
  nor (_11493_, _11492_, _04951_);
  nor (_11494_, _11493_, _01602_);
  and (_11495_, _11494_, _11473_);
  and (_11496_, _08009_, _04177_);
  nor (_11497_, _11496_, _01923_);
  and (_11498_, _11497_, _11460_);
  nor (_11499_, _11498_, _11495_);
  nor (_11500_, _11499_, _06278_);
  nor (_11501_, _08023_, _06680_);
  nor (_11502_, _11501_, _05049_);
  and (_11503_, _04177_, _02676_);
  nor (_11504_, _11503_, _04979_);
  or (_11505_, _11504_, _11502_);
  and (_11506_, _11505_, _11460_);
  nor (_11507_, _11506_, _11500_);
  nor (_11508_, _11507_, _02135_);
  nor (_11509_, _11508_, _11466_);
  nor (_11510_, _11509_, _02039_);
  nor (_11511_, _11510_, _11463_);
  nor (_11512_, _11511_, _02130_);
  nor (_11513_, _11469_, _05741_);
  nor (_11514_, _11513_, _02131_);
  and (_11515_, _11514_, _11478_);
  nor (_11516_, _11515_, _11512_);
  nor (_11517_, _11516_, _02128_);
  and (_11518_, _11503_, _04452_);
  nor (_11519_, _11518_, _05104_);
  nand (_11520_, _11477_, _04452_);
  and (_11521_, _11520_, _02126_);
  or (_11522_, _11521_, _11519_);
  and (_11523_, _11522_, _11460_);
  or (_11524_, _11523_, _02164_);
  nor (_11525_, _11524_, _11517_);
  nor (_11526_, _11525_, _11459_);
  nor (_11527_, _11526_, _01594_);
  nor (_11528_, _11469_, _11457_);
  and (_11529_, _11528_, _01594_);
  nor (_11530_, _11529_, _11527_);
  or (_11531_, _11530_, _26506_);
  or (_11532_, _26505_, \oc8051_golden_model_1.PCON [1]);
  and (_11533_, _11532_, _25964_);
  and (_27825_, _11533_, _11531_);
  not (_11534_, \oc8051_golden_model_1.PCON [2]);
  nor (_11535_, _04177_, _11534_);
  nor (_11536_, _11535_, _05739_);
  not (_11537_, _11536_);
  and (_11538_, _04177_, _05563_);
  nor (_11539_, _11538_, _11535_);
  nor (_11540_, _11539_, _05076_);
  and (_11541_, _11540_, _11537_);
  and (_11542_, _04177_, _03564_);
  nor (_11543_, _11542_, _11535_);
  or (_11544_, _11543_, _05513_);
  and (_11545_, _04177_, \oc8051_golden_model_1.ACC [2]);
  nor (_11546_, _11545_, _11535_);
  nor (_11547_, _11546_, _05488_);
  nor (_11548_, _04571_, _11534_);
  or (_11549_, _11548_, _11547_);
  and (_11550_, _11549_, _02438_);
  nor (_11551_, _08095_, _06680_);
  nor (_11552_, _11551_, _11535_);
  nor (_11553_, _11552_, _02438_);
  or (_11554_, _11553_, _11550_);
  and (_11555_, _11554_, _05487_);
  nor (_11556_, _06680_, _03272_);
  nor (_11557_, _11556_, _11535_);
  nor (_11558_, _11557_, _05487_);
  nor (_11559_, _11558_, _11555_);
  nor (_11560_, _11559_, _01963_);
  nor (_11561_, _11546_, _01964_);
  nor (_11562_, _11561_, _04950_);
  not (_11563_, _11562_);
  nor (_11564_, _11563_, _11560_);
  and (_11565_, _11557_, _04950_);
  or (_11566_, _11565_, _04951_);
  or (_11567_, _11566_, _11564_);
  and (_11568_, _11567_, _01923_);
  and (_11569_, _11568_, _11544_);
  nor (_11570_, _08216_, _06680_);
  or (_11571_, _11535_, _01923_);
  nor (_11572_, _11571_, _11570_);
  or (_11573_, _11572_, _02019_);
  nor (_11574_, _11573_, _11569_);
  nand (_11575_, _11539_, _05049_);
  and (_11576_, _11575_, _06278_);
  nor (_11577_, _11576_, _11574_);
  and (_11578_, _08230_, _04177_);
  nor (_11579_, _11578_, _11535_);
  and (_11580_, _11579_, _02018_);
  nor (_11581_, _11580_, _11577_);
  and (_11582_, _11581_, _02136_);
  and (_11583_, _08237_, _04177_);
  nor (_11584_, _11583_, _11535_);
  nor (_11585_, _11584_, _02136_);
  or (_11586_, _11585_, _11582_);
  and (_11587_, _11586_, _05076_);
  nor (_11588_, _11587_, _11541_);
  nor (_11589_, _11588_, _02130_);
  or (_11590_, _11536_, _02131_);
  nor (_11591_, _11590_, _11546_);
  or (_11592_, _11591_, _02016_);
  nor (_11593_, _11592_, _11589_);
  nor (_11594_, _08229_, _06680_);
  nor (_11595_, _11594_, _11535_);
  and (_11596_, _11595_, _02016_);
  nor (_11597_, _11596_, _11593_);
  and (_11598_, _11597_, _05474_);
  nor (_11599_, _08236_, _06680_);
  nor (_11600_, _11599_, _11535_);
  nor (_11601_, _11600_, _05474_);
  or (_11602_, _11601_, _11598_);
  and (_11603_, _11602_, _02168_);
  nor (_11604_, _11552_, _02168_);
  or (_11605_, _11604_, _01594_);
  nor (_11606_, _11605_, _11603_);
  and (_11607_, _08285_, _04177_);
  nor (_11608_, _11607_, _11535_);
  and (_11609_, _11608_, _01594_);
  nor (_11610_, _11609_, _11606_);
  or (_11611_, _11610_, _26506_);
  or (_11612_, _26505_, \oc8051_golden_model_1.PCON [2]);
  and (_11613_, _11612_, _25964_);
  and (_27828_, _11613_, _11611_);
  not (_11614_, \oc8051_golden_model_1.PCON [3]);
  nor (_11615_, _04177_, _11614_);
  nor (_11616_, _11615_, _05737_);
  not (_11617_, _11616_);
  and (_11618_, _04177_, _05529_);
  nor (_11619_, _11618_, _11615_);
  nor (_11620_, _11619_, _05076_);
  and (_11621_, _11620_, _11617_);
  and (_11622_, _04177_, \oc8051_golden_model_1.ACC [3]);
  nor (_11623_, _11622_, _11615_);
  nor (_11624_, _11623_, _05488_);
  nor (_11625_, _04571_, _11614_);
  or (_11626_, _11625_, _11624_);
  and (_11627_, _11626_, _02438_);
  nor (_11628_, _08337_, _06680_);
  nor (_11629_, _11628_, _11615_);
  nor (_11630_, _11629_, _02438_);
  or (_11631_, _11630_, _11627_);
  and (_11632_, _11631_, _05487_);
  nor (_11633_, _06680_, _03473_);
  nor (_11634_, _11633_, _11615_);
  nor (_11635_, _11634_, _05487_);
  nor (_11636_, _11635_, _11632_);
  nor (_11637_, _11636_, _01963_);
  nor (_11638_, _11623_, _01964_);
  nor (_11639_, _11638_, _04950_);
  not (_11640_, _11639_);
  nor (_11641_, _11640_, _11637_);
  and (_11642_, _11634_, _04950_);
  or (_11643_, _11642_, _04951_);
  or (_11644_, _11643_, _11641_);
  and (_11645_, _04177_, _03516_);
  nor (_11646_, _11645_, _11615_);
  or (_11647_, _11646_, _05513_);
  and (_11648_, _11647_, _01923_);
  and (_11649_, _11648_, _11644_);
  nor (_11650_, _08425_, _06680_);
  or (_11651_, _11615_, _01923_);
  nor (_11652_, _11651_, _11650_);
  or (_11653_, _11652_, _02019_);
  nor (_11654_, _11653_, _11649_);
  nand (_11655_, _11619_, _05049_);
  and (_11656_, _11655_, _06278_);
  nor (_11657_, _11656_, _11654_);
  and (_11658_, _08441_, _04177_);
  nor (_11659_, _11658_, _11615_);
  and (_11660_, _11659_, _02018_);
  nor (_11661_, _11660_, _11657_);
  and (_11662_, _11661_, _02136_);
  and (_11663_, _08304_, _04177_);
  nor (_11664_, _11663_, _11615_);
  nor (_11665_, _11664_, _02136_);
  or (_11666_, _11665_, _11662_);
  and (_11667_, _11666_, _05076_);
  nor (_11668_, _11667_, _11621_);
  nor (_11669_, _11668_, _02130_);
  or (_11670_, _11616_, _02131_);
  nor (_11671_, _11670_, _11623_);
  or (_11672_, _11671_, _02016_);
  nor (_11673_, _11672_, _11669_);
  nor (_11674_, _08440_, _06680_);
  nor (_11675_, _11674_, _11615_);
  and (_11676_, _11675_, _02016_);
  nor (_11677_, _11676_, _11673_);
  and (_11678_, _11677_, _05474_);
  nor (_11679_, _08303_, _06680_);
  nor (_11680_, _11679_, _11615_);
  nor (_11681_, _11680_, _05474_);
  or (_11682_, _11681_, _11678_);
  and (_11683_, _11682_, _02168_);
  nand (_11684_, _11629_, _01595_);
  and (_11685_, _11684_, _02266_);
  nor (_11686_, _11685_, _11683_);
  and (_11687_, _08507_, _04177_);
  nor (_11688_, _11687_, _11615_);
  and (_11689_, _11688_, _01594_);
  nor (_11690_, _11689_, _11686_);
  or (_11691_, _11690_, _26506_);
  or (_11692_, _26505_, \oc8051_golden_model_1.PCON [3]);
  and (_11693_, _11692_, _25964_);
  and (_27829_, _11693_, _11691_);
  not (_11694_, \oc8051_golden_model_1.PCON [4]);
  nor (_11695_, _04177_, _11694_);
  and (_11696_, _08527_, _04177_);
  nor (_11697_, _11696_, _11695_);
  nor (_11698_, _11697_, _02136_);
  and (_11699_, _04177_, _05524_);
  nor (_11700_, _11699_, _11695_);
  and (_11701_, _11700_, _02019_);
  nor (_11702_, _06680_, _04024_);
  nor (_11703_, _11702_, _11695_);
  and (_11704_, _11703_, _04950_);
  and (_11705_, _04177_, \oc8051_golden_model_1.ACC [4]);
  nor (_11706_, _11705_, _11695_);
  nor (_11707_, _11706_, _05488_);
  nor (_11708_, _04571_, _11694_);
  or (_11709_, _11708_, _11707_);
  and (_11710_, _11709_, _02438_);
  nor (_11711_, _08548_, _06680_);
  nor (_11712_, _11711_, _11695_);
  nor (_11713_, _11712_, _02438_);
  or (_11714_, _11713_, _11710_);
  and (_11715_, _11714_, _05487_);
  nor (_11716_, _11703_, _05487_);
  nor (_11717_, _11716_, _11715_);
  nor (_11718_, _11717_, _01963_);
  nor (_11719_, _11706_, _01964_);
  nor (_11720_, _11719_, _04950_);
  not (_11721_, _11720_);
  nor (_11722_, _11721_, _11718_);
  nor (_11723_, _11722_, _11704_);
  nor (_11724_, _11723_, _04951_);
  and (_11725_, _04177_, _03903_);
  nor (_11726_, _11695_, _05513_);
  not (_11727_, _11726_);
  nor (_11728_, _11727_, _11725_);
  or (_11729_, _11728_, _01602_);
  nor (_11730_, _11729_, _11724_);
  nor (_11731_, _08663_, _06680_);
  nor (_11732_, _11731_, _11695_);
  nor (_11733_, _11732_, _01923_);
  or (_11734_, _11733_, _02019_);
  nor (_11735_, _11734_, _11730_);
  nor (_11736_, _11735_, _11701_);
  or (_11737_, _11736_, _02018_);
  and (_11738_, _08531_, _04177_);
  or (_11739_, _11738_, _11695_);
  or (_11740_, _11739_, _05049_);
  and (_11741_, _11740_, _02136_);
  and (_11742_, _11741_, _11737_);
  nor (_11743_, _11742_, _11698_);
  nor (_11744_, _11743_, _02039_);
  nor (_11745_, _11695_, _08729_);
  not (_11746_, _11745_);
  nor (_11747_, _11700_, _05076_);
  and (_11748_, _11747_, _11746_);
  nor (_11749_, _11748_, _11744_);
  nor (_11750_, _11749_, _02130_);
  or (_11751_, _11745_, _02131_);
  nor (_11752_, _11751_, _11706_);
  or (_11753_, _11752_, _02016_);
  nor (_11754_, _11753_, _11750_);
  nor (_11755_, _08530_, _06680_);
  nor (_11756_, _11755_, _11695_);
  and (_11757_, _11756_, _02016_);
  nor (_11758_, _11757_, _11754_);
  and (_11759_, _11758_, _05474_);
  nor (_11760_, _08526_, _06680_);
  nor (_11761_, _11760_, _11695_);
  nor (_11762_, _11761_, _05474_);
  or (_11763_, _11762_, _11759_);
  and (_11764_, _11763_, _02168_);
  nor (_11765_, _11712_, _02168_);
  or (_11766_, _11765_, _01594_);
  nor (_11767_, _11766_, _11764_);
  and (_11768_, _08732_, _04177_);
  nor (_11769_, _11768_, _11695_);
  and (_11770_, _11769_, _01594_);
  nor (_11771_, _11770_, _11767_);
  or (_11772_, _11771_, _26506_);
  or (_11773_, _26505_, \oc8051_golden_model_1.PCON [4]);
  and (_11774_, _11773_, _25964_);
  and (_27830_, _11774_, _11772_);
  not (_11775_, \oc8051_golden_model_1.PCON [5]);
  nor (_11776_, _04177_, _11775_);
  and (_11777_, _08750_, _04177_);
  nor (_11778_, _11777_, _11776_);
  nor (_11779_, _11778_, _02136_);
  and (_11780_, _04177_, _05548_);
  nor (_11781_, _11780_, _11776_);
  and (_11782_, _11781_, _02019_);
  nor (_11783_, _06680_, _03976_);
  nor (_11784_, _11783_, _11776_);
  and (_11785_, _11784_, _04950_);
  and (_11786_, _04177_, \oc8051_golden_model_1.ACC [5]);
  nor (_11787_, _11786_, _11776_);
  nor (_11788_, _11787_, _01964_);
  nor (_11789_, _11787_, _05488_);
  nor (_11790_, _04571_, _11775_);
  or (_11791_, _11790_, _11789_);
  and (_11792_, _11791_, _02438_);
  nor (_11793_, _08771_, _06680_);
  nor (_11794_, _11793_, _11776_);
  nor (_11795_, _11794_, _02438_);
  or (_11796_, _11795_, _11792_);
  and (_11797_, _11796_, _05487_);
  nor (_11798_, _11784_, _05487_);
  nor (_11799_, _11798_, _11797_);
  nor (_11800_, _11799_, _01963_);
  or (_11801_, _11800_, _04950_);
  nor (_11802_, _11801_, _11788_);
  nor (_11803_, _11802_, _11785_);
  nor (_11804_, _11803_, _04951_);
  and (_11805_, _04177_, _03850_);
  nor (_11806_, _11776_, _05513_);
  not (_11807_, _11806_);
  nor (_11808_, _11807_, _11805_);
  or (_11809_, _11808_, _01602_);
  nor (_11810_, _11809_, _11804_);
  nor (_11811_, _08874_, _06680_);
  nor (_11812_, _11811_, _11776_);
  nor (_11813_, _11812_, _01923_);
  or (_11814_, _11813_, _02019_);
  nor (_11815_, _11814_, _11810_);
  nor (_11816_, _11815_, _11782_);
  or (_11817_, _11816_, _02018_);
  and (_11818_, _08890_, _04177_);
  or (_11819_, _11818_, _11776_);
  or (_11820_, _11819_, _05049_);
  and (_11821_, _11820_, _02136_);
  and (_11822_, _11821_, _11817_);
  nor (_11823_, _11822_, _11779_);
  nor (_11824_, _11823_, _02039_);
  nor (_11825_, _11776_, _08946_);
  not (_11826_, _11825_);
  nor (_11827_, _11781_, _05076_);
  and (_11828_, _11827_, _11826_);
  nor (_11829_, _11828_, _11824_);
  nor (_11830_, _11829_, _02130_);
  or (_11831_, _11825_, _02131_);
  nor (_11832_, _11831_, _11787_);
  or (_11833_, _11832_, _02016_);
  nor (_11834_, _11833_, _11830_);
  nor (_11835_, _08889_, _06680_);
  nor (_11836_, _11835_, _11776_);
  and (_11837_, _11836_, _02016_);
  nor (_11838_, _11837_, _11834_);
  and (_11839_, _11838_, _05474_);
  nor (_11840_, _08749_, _06680_);
  nor (_11841_, _11840_, _11776_);
  nor (_11842_, _11841_, _05474_);
  or (_11843_, _11842_, _11839_);
  and (_11844_, _11843_, _02168_);
  nor (_11845_, _11794_, _02168_);
  or (_11846_, _11845_, _01594_);
  nor (_11847_, _11846_, _11844_);
  and (_11848_, _08949_, _04177_);
  nor (_11849_, _11848_, _11776_);
  and (_11850_, _11849_, _01594_);
  nor (_11851_, _11850_, _11847_);
  or (_11852_, _11851_, _26506_);
  or (_11853_, _26505_, \oc8051_golden_model_1.PCON [5]);
  and (_11854_, _11853_, _25964_);
  and (_27831_, _11854_, _11852_);
  not (_11855_, \oc8051_golden_model_1.PCON [6]);
  nor (_11856_, _04177_, _11855_);
  and (_11857_, _08975_, _04177_);
  nor (_11858_, _11857_, _11856_);
  nor (_11859_, _11858_, _02136_);
  and (_11860_, _04177_, _03748_);
  or (_11861_, _11860_, _11856_);
  and (_11862_, _11861_, _04951_);
  and (_11863_, _04177_, \oc8051_golden_model_1.ACC [6]);
  nor (_11864_, _11863_, _11856_);
  nor (_11865_, _11864_, _01964_);
  nor (_11866_, _11864_, _05488_);
  nor (_11867_, _04571_, _11855_);
  or (_11868_, _11867_, _11866_);
  and (_11869_, _11868_, _02438_);
  nor (_11870_, _08995_, _06680_);
  nor (_11871_, _11870_, _11856_);
  nor (_11872_, _11871_, _02438_);
  or (_11873_, _11872_, _11869_);
  and (_11874_, _11873_, _05487_);
  nor (_11875_, _06680_, _04074_);
  nor (_11876_, _11875_, _11856_);
  nor (_11877_, _11876_, _05487_);
  nor (_11878_, _11877_, _11874_);
  nor (_11879_, _11878_, _01963_);
  or (_11880_, _11879_, _04950_);
  nor (_11881_, _11880_, _11865_);
  and (_11882_, _11876_, _04950_);
  or (_11883_, _11882_, _04951_);
  nor (_11884_, _11883_, _11881_);
  or (_11885_, _11884_, _11862_);
  and (_11886_, _11885_, _01923_);
  nor (_11887_, _09096_, _06680_);
  nor (_11888_, _11887_, _11856_);
  nor (_11889_, _11888_, _01923_);
  or (_11890_, _11889_, _06278_);
  or (_11891_, _11890_, _11886_);
  and (_11892_, _09112_, _04177_);
  or (_11893_, _11856_, _05049_);
  or (_11894_, _11893_, _11892_);
  and (_11895_, _04177_, _09103_);
  nor (_11896_, _11895_, _11856_);
  and (_11897_, _11896_, _02019_);
  nor (_11898_, _11897_, _02135_);
  and (_11899_, _11898_, _11894_);
  and (_11900_, _11899_, _11891_);
  nor (_11901_, _11900_, _11859_);
  nor (_11902_, _11901_, _02039_);
  nor (_11903_, _11856_, _05735_);
  not (_11904_, _11903_);
  nor (_11905_, _11896_, _05076_);
  and (_11906_, _11905_, _11904_);
  nor (_11907_, _11906_, _11902_);
  nor (_11908_, _11907_, _02130_);
  or (_11909_, _11903_, _02131_);
  nor (_11910_, _11909_, _11864_);
  or (_11911_, _11910_, _02016_);
  nor (_11912_, _11911_, _11908_);
  nor (_11913_, _09111_, _06680_);
  nor (_11914_, _11913_, _11856_);
  and (_11915_, _11914_, _02016_);
  nor (_11916_, _11915_, _11912_);
  and (_11917_, _11916_, _05474_);
  nor (_11918_, _08974_, _06680_);
  nor (_11919_, _11918_, _11856_);
  nor (_11920_, _11919_, _05474_);
  or (_11921_, _11920_, _11917_);
  and (_11922_, _11921_, _02168_);
  nor (_11923_, _11871_, _02168_);
  or (_11924_, _11923_, _01594_);
  nor (_11925_, _11924_, _11922_);
  and (_11926_, _08965_, _04177_);
  nor (_11927_, _11926_, _11856_);
  and (_11928_, _11927_, _01594_);
  nor (_11929_, _11928_, _11925_);
  or (_11930_, _11929_, _26506_);
  or (_11931_, _26505_, \oc8051_golden_model_1.PCON [6]);
  and (_11932_, _11931_, _25964_);
  and (_27832_, _11932_, _11930_);
  not (_11933_, \oc8051_golden_model_1.SBUF [0]);
  nor (_11934_, _04180_, _11933_);
  nor (_11935_, _04405_, _06599_);
  nor (_11936_, _11935_, _11934_);
  and (_11937_, _11936_, _02266_);
  and (_11938_, _04180_, \oc8051_golden_model_1.ACC [0]);
  nor (_11939_, _11938_, _11934_);
  nor (_11940_, _11939_, _01964_);
  nor (_11941_, _11940_, _04950_);
  nor (_11942_, _11936_, _02438_);
  nor (_11943_, _04571_, _11933_);
  nor (_11944_, _11939_, _05488_);
  nor (_11945_, _11944_, _11943_);
  nor (_11946_, _11945_, _01969_);
  or (_11947_, _11946_, _01967_);
  nor (_11948_, _11947_, _11942_);
  or (_11949_, _11948_, _01963_);
  and (_11950_, _11949_, _11941_);
  and (_11951_, _04180_, _03334_);
  nor (_11952_, _04950_, _01967_);
  or (_11953_, _11952_, _11934_);
  nor (_11954_, _11953_, _11951_);
  nor (_11955_, _11954_, _11950_);
  nor (_11956_, _11955_, _04951_);
  and (_11957_, _04180_, _03677_);
  nor (_11958_, _11934_, _05513_);
  not (_11959_, _11958_);
  nor (_11960_, _11959_, _11957_);
  nor (_11961_, _11960_, _11956_);
  nor (_11962_, _11961_, _01602_);
  nor (_11963_, _07815_, _06599_);
  or (_11964_, _11934_, _01923_);
  nor (_11965_, _11964_, _11963_);
  or (_11966_, _11965_, _02019_);
  nor (_11967_, _11966_, _11962_);
  and (_11968_, _04180_, _05531_);
  nor (_11969_, _11968_, _11934_);
  nand (_11970_, _11969_, _05049_);
  and (_11971_, _11970_, _06278_);
  nor (_11972_, _11971_, _11967_);
  and (_11973_, _07829_, _04180_);
  nor (_11974_, _11973_, _11934_);
  and (_11975_, _11974_, _02018_);
  nor (_11976_, _11975_, _11972_);
  and (_11977_, _11976_, _02136_);
  and (_11978_, _07834_, _04180_);
  nor (_11979_, _11978_, _11934_);
  nor (_11980_, _11979_, _02136_);
  or (_11981_, _11980_, _11977_);
  and (_11982_, _11981_, _05076_);
  or (_11983_, _11969_, _05076_);
  nor (_11984_, _11983_, _11935_);
  nor (_11985_, _11984_, _11982_);
  nor (_11986_, _11985_, _02130_);
  and (_11987_, _07833_, _04180_);
  or (_11988_, _11987_, _11934_);
  and (_11989_, _11988_, _02130_);
  or (_11990_, _11989_, _11986_);
  and (_11991_, _11990_, _05104_);
  nor (_11992_, _07828_, _06599_);
  nor (_11993_, _11992_, _11934_);
  nor (_11994_, _11993_, _05104_);
  or (_11995_, _11994_, _11991_);
  and (_11996_, _11995_, _05474_);
  nor (_11997_, _07696_, _06599_);
  nor (_11998_, _11997_, _11934_);
  nor (_11999_, _11998_, _05474_);
  nor (_12000_, _11999_, _02266_);
  not (_12001_, _12000_);
  nor (_12002_, _12001_, _11996_);
  nor (_12003_, _12002_, _11937_);
  or (_12004_, _12003_, _26506_);
  or (_12005_, _26505_, \oc8051_golden_model_1.SBUF [0]);
  and (_12006_, _12005_, _25964_);
  and (_27833_, _12006_, _12004_);
  nor (_12007_, _04180_, \oc8051_golden_model_1.SBUF [1]);
  and (_12008_, _07909_, _04180_);
  nor (_12009_, _12008_, _12007_);
  nor (_12010_, _12009_, _02168_);
  not (_12011_, _12007_);
  nor (_12012_, _08029_, _06599_);
  nor (_12013_, _12012_, _02136_);
  and (_12014_, _12013_, _12011_);
  and (_12015_, _04180_, _03613_);
  not (_12016_, \oc8051_golden_model_1.SBUF [1]);
  nor (_12017_, _04180_, _12016_);
  nor (_12018_, _12017_, _05513_);
  not (_12019_, _12018_);
  nor (_12020_, _12019_, _12015_);
  not (_12021_, _12020_);
  nor (_12022_, _06599_, _03393_);
  nor (_12023_, _12022_, _12017_);
  and (_12024_, _12023_, _04950_);
  and (_12025_, _04180_, _01705_);
  nor (_12026_, _12025_, _12007_);
  and (_12027_, _12026_, _01963_);
  and (_12028_, _12026_, _04571_);
  nor (_12029_, _04571_, _12016_);
  or (_12030_, _12029_, _12028_);
  and (_12031_, _12030_, _02438_);
  and (_12032_, _12009_, _01969_);
  or (_12033_, _12032_, _12031_);
  and (_12034_, _12033_, _05487_);
  nor (_12035_, _12023_, _05487_);
  nor (_12036_, _12035_, _12034_);
  nor (_12037_, _12036_, _01963_);
  or (_12038_, _12037_, _04950_);
  nor (_12039_, _12038_, _12027_);
  nor (_12040_, _12039_, _12024_);
  nor (_12041_, _12040_, _04951_);
  nor (_12042_, _12041_, _01602_);
  and (_12043_, _12042_, _12021_);
  and (_12044_, _08009_, _04180_);
  nor (_12045_, _12044_, _01923_);
  and (_12046_, _12045_, _12011_);
  nor (_12047_, _12046_, _12043_);
  nor (_12048_, _12047_, _06278_);
  nor (_12049_, _08023_, _06599_);
  nor (_12050_, _12049_, _05049_);
  and (_12051_, _04180_, _02676_);
  nor (_12052_, _12051_, _04979_);
  or (_12053_, _12052_, _12050_);
  and (_12054_, _12053_, _12011_);
  nor (_12055_, _12054_, _12048_);
  nor (_12056_, _12055_, _02135_);
  nor (_12057_, _12056_, _12014_);
  nor (_12058_, _12057_, _02039_);
  nor (_12059_, _07893_, _06599_);
  nor (_12060_, _12059_, _05076_);
  and (_12061_, _12060_, _12011_);
  nor (_12062_, _12061_, _12058_);
  nor (_12063_, _12062_, _02130_);
  nor (_12064_, _12017_, _05741_);
  nor (_12065_, _12064_, _02131_);
  and (_12066_, _12065_, _12026_);
  nor (_12067_, _12066_, _12063_);
  nor (_12068_, _12067_, _02128_);
  and (_12069_, _12051_, _04452_);
  nor (_12070_, _12069_, _05104_);
  and (_12071_, _12025_, _04452_);
  nor (_12072_, _12071_, _05474_);
  or (_12073_, _12072_, _12070_);
  and (_12074_, _12073_, _12011_);
  or (_12075_, _12074_, _02164_);
  nor (_12076_, _12075_, _12068_);
  nor (_12077_, _12076_, _12010_);
  nor (_12078_, _12077_, _01594_);
  nor (_12079_, _12017_, _12008_);
  and (_12080_, _12079_, _01594_);
  nor (_12081_, _12080_, _12078_);
  or (_12082_, _12081_, _26506_);
  or (_12083_, _26505_, \oc8051_golden_model_1.SBUF [1]);
  and (_12084_, _12083_, _25964_);
  and (_27834_, _12084_, _12082_);
  not (_12085_, \oc8051_golden_model_1.SBUF [2]);
  nor (_12086_, _04180_, _12085_);
  and (_12087_, _04180_, _03564_);
  nor (_12088_, _12087_, _12086_);
  or (_12089_, _12088_, _05513_);
  and (_12090_, _04180_, \oc8051_golden_model_1.ACC [2]);
  nor (_12091_, _12090_, _12086_);
  nor (_12092_, _12091_, _01964_);
  nor (_12093_, _12091_, _05488_);
  nor (_12094_, _04571_, _12085_);
  or (_12095_, _12094_, _12093_);
  and (_12096_, _12095_, _02438_);
  nor (_12097_, _08095_, _06599_);
  nor (_12098_, _12097_, _12086_);
  nor (_12099_, _12098_, _02438_);
  or (_12100_, _12099_, _12096_);
  and (_12101_, _12100_, _05487_);
  nor (_12102_, _06599_, _03272_);
  nor (_12103_, _12102_, _12086_);
  nor (_12104_, _12103_, _05487_);
  nor (_12105_, _12104_, _12101_);
  nor (_12106_, _12105_, _01963_);
  or (_12107_, _12106_, _04950_);
  nor (_12108_, _12107_, _12092_);
  and (_12109_, _12103_, _04950_);
  or (_12110_, _12109_, _04951_);
  or (_12111_, _12110_, _12108_);
  and (_12112_, _12111_, _01923_);
  and (_12113_, _12112_, _12089_);
  nor (_12114_, _08216_, _06599_);
  or (_12115_, _12086_, _01923_);
  nor (_12116_, _12115_, _12114_);
  or (_12117_, _12116_, _02019_);
  nor (_12118_, _12117_, _12113_);
  and (_12119_, _04180_, _05563_);
  nor (_12120_, _12119_, _12086_);
  nand (_12121_, _12120_, _05049_);
  and (_12122_, _12121_, _06278_);
  nor (_12123_, _12122_, _12118_);
  and (_12125_, _08230_, _04180_);
  nor (_12126_, _12125_, _12086_);
  and (_12128_, _12126_, _02018_);
  nor (_12129_, _12128_, _12123_);
  and (_12131_, _12129_, _02136_);
  and (_12132_, _08237_, _04180_);
  nor (_12134_, _12132_, _12086_);
  nor (_12135_, _12134_, _02136_);
  or (_12137_, _12135_, _12131_);
  and (_12138_, _12137_, _05076_);
  nor (_12140_, _12086_, _05739_);
  not (_12141_, _12140_);
  nor (_12143_, _12120_, _05076_);
  and (_12144_, _12143_, _12141_);
  nor (_12146_, _12144_, _12138_);
  nor (_12147_, _12146_, _02130_);
  or (_12149_, _12140_, _02131_);
  nor (_12150_, _12149_, _12091_);
  or (_12152_, _12150_, _02016_);
  nor (_12153_, _12152_, _12147_);
  nor (_12155_, _08229_, _06599_);
  nor (_12156_, _12155_, _12086_);
  and (_12158_, _12156_, _02016_);
  nor (_12159_, _12158_, _12153_);
  and (_12161_, _12159_, _05474_);
  nor (_12162_, _08236_, _06599_);
  nor (_12163_, _12162_, _12086_);
  nor (_12164_, _12163_, _05474_);
  or (_12165_, _12164_, _12161_);
  and (_12166_, _12165_, _02168_);
  nor (_12167_, _12098_, _02168_);
  or (_12168_, _12167_, _01594_);
  nor (_12169_, _12168_, _12166_);
  and (_12170_, _08285_, _04180_);
  nor (_12171_, _12170_, _12086_);
  and (_12172_, _12171_, _01594_);
  nor (_12173_, _12172_, _12169_);
  or (_12174_, _12173_, _26506_);
  or (_12175_, _26505_, \oc8051_golden_model_1.SBUF [2]);
  and (_12176_, _12175_, _25964_);
  and (_27835_, _12176_, _12174_);
  not (_12177_, \oc8051_golden_model_1.SBUF [3]);
  nor (_12178_, _04180_, _12177_);
  nor (_12179_, _12178_, _05737_);
  not (_12180_, _12179_);
  and (_12181_, _04180_, _05529_);
  nor (_12182_, _12181_, _12178_);
  nor (_12183_, _12182_, _05076_);
  and (_12184_, _12183_, _12180_);
  and (_12185_, _08304_, _04180_);
  nor (_12186_, _12185_, _12178_);
  nor (_12187_, _12186_, _02136_);
  and (_12188_, _04180_, _03516_);
  or (_12189_, _12188_, _12178_);
  and (_12190_, _12189_, _04951_);
  and (_12191_, _04180_, \oc8051_golden_model_1.ACC [3]);
  nor (_12192_, _12191_, _12178_);
  nor (_12193_, _12192_, _01964_);
  nor (_12194_, _12192_, _05488_);
  nor (_12195_, _04571_, _12177_);
  or (_12196_, _12195_, _12194_);
  and (_12197_, _12196_, _02438_);
  nor (_12198_, _08337_, _06599_);
  nor (_12199_, _12198_, _12178_);
  nor (_12200_, _12199_, _02438_);
  or (_12201_, _12200_, _12197_);
  and (_12202_, _12201_, _05487_);
  nor (_12203_, _06599_, _03473_);
  nor (_12204_, _12203_, _12178_);
  nor (_12205_, _12204_, _05487_);
  nor (_12206_, _12205_, _12202_);
  nor (_12207_, _12206_, _01963_);
  or (_12209_, _12207_, _04950_);
  nor (_12211_, _12209_, _12193_);
  and (_12212_, _12204_, _04950_);
  or (_12214_, _12212_, _04951_);
  nor (_12215_, _12214_, _12211_);
  or (_12217_, _12215_, _12190_);
  and (_12218_, _12217_, _01923_);
  nor (_12220_, _08425_, _06599_);
  nor (_12221_, _12220_, _12178_);
  nor (_12223_, _12221_, _01923_);
  or (_12224_, _12223_, _06278_);
  or (_12226_, _12224_, _12218_);
  and (_12227_, _08441_, _04180_);
  or (_12229_, _12178_, _05049_);
  or (_12230_, _12229_, _12227_);
  and (_12232_, _12182_, _02019_);
  nor (_12233_, _12232_, _02135_);
  and (_12235_, _12233_, _12230_);
  and (_12236_, _12235_, _12226_);
  nor (_12238_, _12236_, _12187_);
  nor (_12239_, _12238_, _02039_);
  nor (_12241_, _12239_, _12184_);
  nor (_12242_, _12241_, _02130_);
  or (_12243_, _12179_, _02131_);
  nor (_12244_, _12243_, _12192_);
  or (_12245_, _12244_, _02016_);
  nor (_12246_, _12245_, _12242_);
  nor (_12247_, _08440_, _06599_);
  nor (_12248_, _12247_, _12178_);
  and (_12249_, _12248_, _02016_);
  nor (_12250_, _12249_, _12246_);
  and (_12251_, _12250_, _05474_);
  nor (_12252_, _08303_, _06599_);
  nor (_12253_, _12252_, _12178_);
  nor (_12254_, _12253_, _05474_);
  or (_12255_, _12254_, _12251_);
  and (_12256_, _12255_, _02168_);
  nor (_12257_, _12199_, _02168_);
  or (_12258_, _12257_, _01594_);
  nor (_12259_, _12258_, _12256_);
  and (_12260_, _08507_, _04180_);
  nor (_12261_, _12260_, _12178_);
  and (_12262_, _12261_, _01594_);
  nor (_12263_, _12262_, _12259_);
  or (_12264_, _12263_, _26506_);
  or (_12265_, _26505_, \oc8051_golden_model_1.SBUF [3]);
  and (_12266_, _12265_, _25964_);
  and (_27836_, _12266_, _12264_);
  not (_12267_, \oc8051_golden_model_1.SBUF [4]);
  nor (_12268_, _04180_, _12267_);
  and (_12269_, _08527_, _04180_);
  nor (_12270_, _12269_, _12268_);
  nor (_12271_, _12270_, _02136_);
  and (_12272_, _04180_, _05524_);
  nor (_12273_, _12272_, _12268_);
  and (_12274_, _12273_, _02019_);
  and (_12275_, _04180_, \oc8051_golden_model_1.ACC [4]);
  nor (_12276_, _12275_, _12268_);
  nor (_12277_, _12276_, _01964_);
  nor (_12278_, _12276_, _05488_);
  nor (_12279_, _04571_, _12267_);
  or (_12280_, _12279_, _12278_);
  and (_12281_, _12280_, _02438_);
  nor (_12282_, _08548_, _06599_);
  nor (_12283_, _12282_, _12268_);
  nor (_12284_, _12283_, _02438_);
  or (_12285_, _12284_, _12281_);
  and (_12286_, _12285_, _05487_);
  nor (_12287_, _06599_, _04024_);
  nor (_12288_, _12287_, _12268_);
  nor (_12289_, _12288_, _05487_);
  nor (_12290_, _12289_, _12286_);
  nor (_12291_, _12290_, _01963_);
  or (_12292_, _12291_, _04950_);
  nor (_12293_, _12292_, _12277_);
  and (_12294_, _12288_, _04950_);
  nor (_12295_, _12294_, _12293_);
  nor (_12296_, _12295_, _04951_);
  and (_12297_, _04180_, _03903_);
  nor (_12298_, _12268_, _05513_);
  not (_12299_, _12298_);
  nor (_12300_, _12299_, _12297_);
  or (_12301_, _12300_, _01602_);
  nor (_12302_, _12301_, _12296_);
  nor (_12303_, _08663_, _06599_);
  nor (_12304_, _12303_, _12268_);
  nor (_12305_, _12304_, _01923_);
  or (_12306_, _12305_, _02019_);
  nor (_12307_, _12306_, _12302_);
  nor (_12308_, _12307_, _12274_);
  or (_12309_, _12308_, _02018_);
  and (_12310_, _08531_, _04180_);
  or (_12311_, _12310_, _12268_);
  or (_12312_, _12311_, _05049_);
  and (_12313_, _12312_, _02136_);
  and (_12314_, _12313_, _12309_);
  nor (_12315_, _12314_, _12271_);
  nor (_12316_, _12315_, _02039_);
  nor (_12317_, _12268_, _08729_);
  not (_12318_, _12317_);
  nor (_12319_, _12273_, _05076_);
  and (_12320_, _12319_, _12318_);
  nor (_12321_, _12320_, _12316_);
  nor (_12322_, _12321_, _02130_);
  or (_12323_, _12317_, _02131_);
  nor (_12324_, _12323_, _12276_);
  or (_12325_, _12324_, _02016_);
  nor (_12326_, _12325_, _12322_);
  nor (_12327_, _08530_, _06599_);
  nor (_12328_, _12327_, _12268_);
  and (_12329_, _12328_, _02016_);
  nor (_12330_, _12329_, _12326_);
  and (_12331_, _12330_, _05474_);
  nor (_12332_, _08526_, _06599_);
  nor (_12333_, _12332_, _12268_);
  nor (_12334_, _12333_, _05474_);
  or (_12335_, _12334_, _12331_);
  and (_12336_, _12335_, _02168_);
  nor (_12337_, _12283_, _02168_);
  or (_12338_, _12337_, _01594_);
  nor (_12339_, _12338_, _12336_);
  and (_12340_, _08732_, _04180_);
  nor (_12341_, _12340_, _12268_);
  and (_12342_, _12341_, _01594_);
  nor (_12343_, _12342_, _12339_);
  or (_12344_, _12343_, _26506_);
  or (_12345_, _26505_, \oc8051_golden_model_1.SBUF [4]);
  and (_12346_, _12345_, _25964_);
  and (_27837_, _12346_, _12344_);
  not (_12347_, \oc8051_golden_model_1.SBUF [5]);
  nor (_12348_, _04180_, _12347_);
  nor (_12349_, _12348_, _08946_);
  not (_12350_, _12349_);
  and (_12351_, _04180_, _05548_);
  nor (_12352_, _12351_, _12348_);
  nor (_12353_, _12352_, _05076_);
  and (_12354_, _12353_, _12350_);
  and (_12355_, _08750_, _04180_);
  nor (_12356_, _12355_, _12348_);
  nor (_12357_, _12356_, _02136_);
  nor (_12358_, _08874_, _06599_);
  or (_12359_, _12348_, _01923_);
  or (_12360_, _12359_, _12358_);
  nor (_12361_, _08771_, _06599_);
  nor (_12362_, _12361_, _12348_);
  nor (_12363_, _12362_, _02438_);
  nor (_12364_, _04571_, _12347_);
  and (_12365_, _04180_, \oc8051_golden_model_1.ACC [5]);
  nor (_12366_, _12365_, _12348_);
  nor (_12367_, _12366_, _05488_);
  nor (_12368_, _12367_, _12364_);
  nor (_12369_, _12368_, _01969_);
  or (_12370_, _12369_, _12363_);
  and (_12371_, _12370_, _05487_);
  nor (_12372_, _06599_, _03976_);
  nor (_12373_, _12372_, _12348_);
  nor (_12374_, _12373_, _05487_);
  or (_12375_, _12374_, _12371_);
  and (_12376_, _12375_, _01964_);
  nor (_12377_, _12366_, _01964_);
  nor (_12378_, _12377_, _04950_);
  not (_12379_, _12378_);
  nor (_12380_, _12379_, _12376_);
  and (_12381_, _12373_, _04950_);
  or (_12382_, _12381_, _04951_);
  nor (_12383_, _12382_, _12380_);
  and (_12384_, _04180_, _03850_);
  or (_12385_, _12384_, _12348_);
  and (_12386_, _12385_, _04951_);
  or (_12387_, _12386_, _01602_);
  or (_12388_, _12387_, _12383_);
  and (_12389_, _12388_, _12360_);
  and (_12390_, _12389_, _04979_);
  nor (_12391_, _12352_, _04979_);
  or (_12392_, _12391_, _12390_);
  or (_12393_, _12392_, _02018_);
  and (_12394_, _08890_, _04180_);
  or (_12395_, _12394_, _12348_);
  or (_12396_, _12395_, _05049_);
  and (_12397_, _12396_, _02136_);
  and (_12398_, _12397_, _12393_);
  nor (_12399_, _12398_, _12357_);
  nor (_12400_, _12399_, _02039_);
  nor (_12401_, _12400_, _12354_);
  nor (_12402_, _12401_, _02130_);
  or (_12403_, _12349_, _02131_);
  nor (_12404_, _12403_, _12366_);
  or (_12405_, _12404_, _02016_);
  nor (_12406_, _12405_, _12402_);
  nor (_12407_, _08889_, _06599_);
  nor (_12408_, _12407_, _12348_);
  and (_12409_, _12408_, _02016_);
  nor (_12410_, _12409_, _12406_);
  and (_12411_, _12410_, _05474_);
  nor (_12412_, _08749_, _06599_);
  nor (_12413_, _12412_, _12348_);
  nor (_12414_, _12413_, _05474_);
  or (_12415_, _12414_, _12411_);
  and (_12416_, _12415_, _02168_);
  nor (_12417_, _12362_, _02168_);
  or (_12418_, _12417_, _01594_);
  nor (_12419_, _12418_, _12416_);
  and (_12420_, _08949_, _04180_);
  nor (_12421_, _12420_, _12348_);
  and (_12422_, _12421_, _01594_);
  nor (_12423_, _12422_, _12419_);
  or (_12424_, _12423_, _26506_);
  or (_12425_, _26505_, \oc8051_golden_model_1.SBUF [5]);
  and (_12426_, _12425_, _25964_);
  and (_27838_, _12426_, _12424_);
  not (_12427_, \oc8051_golden_model_1.SBUF [6]);
  nor (_12428_, _04180_, _12427_);
  and (_12429_, _08975_, _04180_);
  nor (_12430_, _12429_, _12428_);
  nor (_12431_, _12430_, _02136_);
  and (_12432_, _04180_, _03748_);
  or (_12433_, _12432_, _12428_);
  and (_12434_, _12433_, _04951_);
  and (_12435_, _04180_, \oc8051_golden_model_1.ACC [6]);
  nor (_12436_, _12435_, _12428_);
  nor (_12437_, _12436_, _01964_);
  nor (_12438_, _12436_, _05488_);
  nor (_12439_, _04571_, _12427_);
  or (_12440_, _12439_, _12438_);
  and (_12441_, _12440_, _02438_);
  nor (_12442_, _08995_, _06599_);
  nor (_12443_, _12442_, _12428_);
  nor (_12444_, _12443_, _02438_);
  or (_12445_, _12444_, _12441_);
  and (_12446_, _12445_, _05487_);
  nor (_12447_, _06599_, _04074_);
  nor (_12448_, _12447_, _12428_);
  nor (_12449_, _12448_, _05487_);
  nor (_12450_, _12449_, _12446_);
  nor (_12451_, _12450_, _01963_);
  or (_12452_, _12451_, _04950_);
  nor (_12453_, _12452_, _12437_);
  and (_12454_, _12448_, _04950_);
  or (_12455_, _12454_, _04951_);
  nor (_12456_, _12455_, _12453_);
  or (_12457_, _12456_, _12434_);
  and (_12458_, _12457_, _01923_);
  nor (_12459_, _09096_, _06599_);
  nor (_12460_, _12459_, _12428_);
  nor (_12461_, _12460_, _01923_);
  or (_12462_, _12461_, _06278_);
  or (_12463_, _12462_, _12458_);
  and (_12464_, _09112_, _04180_);
  or (_12465_, _12428_, _05049_);
  or (_12466_, _12465_, _12464_);
  and (_12467_, _04180_, _09103_);
  nor (_12468_, _12467_, _12428_);
  and (_12469_, _12468_, _02019_);
  nor (_12470_, _12469_, _02135_);
  and (_12471_, _12470_, _12466_);
  and (_12472_, _12471_, _12463_);
  nor (_12473_, _12472_, _12431_);
  nor (_12474_, _12473_, _02039_);
  nor (_12475_, _12428_, _05735_);
  not (_12476_, _12475_);
  nor (_12477_, _12468_, _05076_);
  and (_12478_, _12477_, _12476_);
  nor (_12479_, _12478_, _12474_);
  nor (_12480_, _12479_, _02130_);
  or (_12481_, _12475_, _02131_);
  nor (_12482_, _12481_, _12436_);
  or (_12483_, _12482_, _02016_);
  nor (_12484_, _12483_, _12480_);
  nor (_12485_, _09111_, _06599_);
  nor (_12486_, _12485_, _12428_);
  and (_12487_, _12486_, _02016_);
  nor (_12488_, _12487_, _12484_);
  and (_12489_, _12488_, _05474_);
  nor (_12490_, _08974_, _06599_);
  nor (_12491_, _12490_, _12428_);
  nor (_12492_, _12491_, _05474_);
  or (_12493_, _12492_, _12489_);
  and (_12494_, _12493_, _02168_);
  nor (_12495_, _12443_, _02168_);
  or (_12496_, _12495_, _01594_);
  nor (_12497_, _12496_, _12494_);
  and (_12498_, _08965_, _04180_);
  nor (_12499_, _12498_, _12428_);
  and (_12500_, _12499_, _01594_);
  nor (_12501_, _12500_, _12497_);
  or (_12502_, _12501_, _26506_);
  or (_12503_, _26505_, \oc8051_golden_model_1.SBUF [6]);
  and (_12504_, _12503_, _25964_);
  and (_27839_, _12504_, _12502_);
  not (_12505_, \oc8051_golden_model_1.SCON [0]);
  nor (_12506_, _04129_, _12505_);
  nor (_12507_, _04405_, _06482_);
  nor (_12508_, _12507_, _12506_);
  nor (_12509_, _12508_, _01595_);
  and (_12510_, _07834_, _04129_);
  nor (_12511_, _12510_, _12506_);
  nor (_12512_, _12511_, _02136_);
  and (_12513_, _04129_, _05531_);
  nor (_12514_, _12513_, _12506_);
  and (_12515_, _12514_, _02019_);
  and (_12516_, _04129_, _03334_);
  nor (_12517_, _12516_, _12506_);
  and (_12518_, _12517_, _04950_);
  and (_12519_, _04129_, \oc8051_golden_model_1.ACC [0]);
  nor (_12520_, _12519_, _12506_);
  and (_12521_, _12520_, _01963_);
  and (_12522_, _12508_, _01969_);
  nor (_12523_, _12520_, _05488_);
  nor (_12524_, _04571_, _12505_);
  or (_12525_, _12524_, _01969_);
  nor (_12526_, _12525_, _12523_);
  or (_12527_, _12526_, _06233_);
  nor (_12528_, _12527_, _12522_);
  nor (_12529_, _12517_, _05487_);
  nor (_12530_, _12529_, _12528_);
  nor (_12531_, _05184_, _12505_);
  and (_12532_, _07725_, _05184_);
  nor (_12533_, _12532_, _12531_);
  nor (_12534_, _12533_, _02223_);
  nor (_12535_, _12534_, _01963_);
  and (_12536_, _12535_, _12530_);
  nor (_12537_, _12536_, _12521_);
  nor (_12538_, _12537_, _01957_);
  nor (_12539_, _12506_, _06229_);
  or (_12540_, _12539_, _01946_);
  nor (_12541_, _12540_, _12538_);
  nor (_12542_, _12508_, _04885_);
  or (_12543_, _12542_, _12541_);
  and (_12544_, _12543_, _01925_);
  nor (_12545_, _07759_, _06519_);
  nor (_12546_, _12545_, _12531_);
  nor (_12547_, _12546_, _01925_);
  or (_12548_, _12547_, _04950_);
  nor (_12549_, _12548_, _12544_);
  nor (_12550_, _12549_, _12518_);
  nor (_12551_, _12550_, _04951_);
  and (_12552_, _04129_, _03677_);
  nor (_12553_, _12506_, _05513_);
  not (_12554_, _12553_);
  nor (_12555_, _12554_, _12552_);
  or (_12556_, _12555_, _01602_);
  nor (_12557_, _12556_, _12551_);
  nor (_12558_, _07815_, _06482_);
  nor (_12559_, _12558_, _12506_);
  nor (_12560_, _12559_, _01923_);
  or (_12561_, _12560_, _02019_);
  nor (_12562_, _12561_, _12557_);
  nor (_12563_, _12562_, _12515_);
  or (_12564_, _12563_, _02018_);
  and (_12565_, _07829_, _04129_);
  or (_12566_, _12565_, _12506_);
  or (_12567_, _12566_, _05049_);
  and (_12568_, _12567_, _02136_);
  and (_12569_, _12568_, _12564_);
  nor (_12570_, _12569_, _12512_);
  nor (_12571_, _12570_, _02039_);
  or (_12572_, _12514_, _05076_);
  nor (_12573_, _12572_, _12507_);
  nor (_12574_, _12573_, _12571_);
  nor (_12575_, _12574_, _02130_);
  nor (_12576_, _12506_, _04405_);
  or (_12577_, _12576_, _02131_);
  nor (_12578_, _12577_, _12520_);
  or (_12579_, _12578_, _02016_);
  nor (_12580_, _12579_, _12575_);
  nor (_12581_, _07828_, _06482_);
  nor (_12582_, _12581_, _12506_);
  and (_12583_, _12582_, _02016_);
  nor (_12584_, _12583_, _12580_);
  and (_12585_, _12584_, _05474_);
  nor (_12586_, _07696_, _06482_);
  nor (_12587_, _12586_, _12506_);
  nor (_12588_, _12587_, _05474_);
  or (_12589_, _12588_, _12585_);
  and (_12590_, _12589_, _02168_);
  nor (_12591_, _12508_, _02168_);
  nor (_12592_, _12591_, _02025_);
  not (_12593_, _12592_);
  nor (_12594_, _12593_, _12590_);
  nor (_12595_, _12506_, _02377_);
  nor (_12596_, _12595_, _12594_);
  and (_12597_, _12596_, _01595_);
  nor (_12598_, _12597_, _12509_);
  nand (_12599_, _12598_, _26505_);
  or (_12600_, _26505_, \oc8051_golden_model_1.SCON [0]);
  and (_12601_, _12600_, _25964_);
  and (_27842_, _12601_, _12599_);
  nor (_12602_, _04129_, \oc8051_golden_model_1.SCON [1]);
  not (_12603_, _12602_);
  nor (_12604_, _08029_, _06482_);
  nor (_12605_, _12604_, _02136_);
  and (_12606_, _12605_, _12603_);
  not (_12607_, \oc8051_golden_model_1.SCON [1]);
  nor (_12608_, _04129_, _12607_);
  and (_12609_, _04129_, _03613_);
  or (_12610_, _12609_, _12608_);
  and (_12611_, _12610_, _04951_);
  nor (_12612_, _07953_, _06519_);
  nor (_12613_, _05184_, _12607_);
  or (_12614_, _12613_, _01925_);
  or (_12615_, _12614_, _12612_);
  and (_12616_, _07909_, _04129_);
  nor (_12617_, _12616_, _12602_);
  nor (_12618_, _12617_, _02438_);
  and (_12619_, _04129_, _01705_);
  nor (_12620_, _12619_, _12602_);
  and (_12621_, _12620_, _04571_);
  nor (_12622_, _04571_, _12607_);
  or (_12623_, _12622_, _01969_);
  nor (_12624_, _12623_, _12621_);
  or (_12625_, _12624_, _06233_);
  nor (_12626_, _12625_, _12618_);
  nor (_12627_, _06482_, _03393_);
  nor (_12628_, _12627_, _12608_);
  nor (_12629_, _12628_, _05487_);
  and (_12630_, _07920_, _05184_);
  nor (_12631_, _12630_, _12613_);
  nor (_12632_, _12631_, _02223_);
  nor (_12633_, _12632_, _12629_);
  nand (_12634_, _12633_, _01964_);
  or (_12635_, _12634_, _12626_);
  or (_12636_, _12620_, _01964_);
  and (_12637_, _12636_, _12635_);
  and (_12638_, _12637_, _06229_);
  and (_12639_, _07907_, _05184_);
  nor (_12640_, _12639_, _12613_);
  nor (_12641_, _12640_, _06229_);
  or (_12642_, _12641_, _12638_);
  and (_12643_, _12642_, _04885_);
  nor (_12644_, _12613_, _07935_);
  or (_12645_, _12644_, _04885_);
  nor (_12646_, _12645_, _12631_);
  or (_12647_, _12646_, _01924_);
  or (_12648_, _12647_, _12643_);
  and (_12649_, _12648_, _12615_);
  nor (_12650_, _12649_, _04950_);
  and (_12651_, _12628_, _04950_);
  or (_12652_, _12651_, _04951_);
  nor (_12653_, _12652_, _12650_);
  or (_12654_, _12653_, _12611_);
  and (_12655_, _12654_, _01923_);
  nor (_12656_, _08009_, _06482_);
  nor (_12657_, _12656_, _12608_);
  nor (_12658_, _12657_, _01923_);
  nor (_12659_, _12658_, _12655_);
  nor (_12660_, _12659_, _06278_);
  nor (_12661_, _08023_, _06482_);
  nor (_12662_, _12661_, _05049_);
  and (_12663_, _04129_, _02676_);
  nor (_12664_, _12663_, _04979_);
  or (_12665_, _12664_, _12662_);
  and (_12666_, _12665_, _12603_);
  nor (_12667_, _12666_, _12660_);
  nor (_12668_, _12667_, _02135_);
  nor (_12669_, _12668_, _12606_);
  nor (_12670_, _12669_, _02039_);
  nor (_12671_, _07893_, _06482_);
  nor (_12672_, _12671_, _05076_);
  and (_12673_, _12672_, _12603_);
  nor (_12674_, _12673_, _12670_);
  nor (_12675_, _12674_, _02130_);
  nor (_12676_, _12608_, _05741_);
  nor (_12677_, _12676_, _02131_);
  and (_12678_, _12677_, _12620_);
  nor (_12679_, _12678_, _12675_);
  nor (_12680_, _12679_, _02128_);
  and (_12681_, _12663_, _04452_);
  nor (_12682_, _12681_, _05104_);
  nand (_12683_, _12619_, _04452_);
  and (_12684_, _12683_, _02126_);
  or (_12685_, _12684_, _12682_);
  and (_12686_, _12685_, _12603_);
  or (_12687_, _12686_, _02164_);
  nor (_12688_, _12687_, _12680_);
  nor (_12689_, _12617_, _02168_);
  or (_12690_, _12689_, _02025_);
  nor (_12691_, _12690_, _12688_);
  nor (_12692_, _12640_, _02377_);
  or (_12693_, _12692_, _01594_);
  nor (_12694_, _12693_, _12691_);
  nor (_12695_, _12616_, _12608_);
  and (_12696_, _12695_, _01594_);
  nor (_12697_, _12696_, _12694_);
  or (_12698_, _12697_, _26506_);
  or (_12699_, _26505_, \oc8051_golden_model_1.SCON [1]);
  and (_12700_, _12699_, _25964_);
  and (_27843_, _12700_, _12698_);
  not (_12701_, \oc8051_golden_model_1.SCON [2]);
  nor (_12702_, _04129_, _12701_);
  and (_12703_, _04129_, _05563_);
  nor (_12704_, _12703_, _12702_);
  and (_12705_, _12704_, _02019_);
  nor (_12706_, _06482_, _03272_);
  nor (_12707_, _12706_, _12702_);
  and (_12708_, _12707_, _04950_);
  nor (_12709_, _08095_, _06482_);
  nor (_12710_, _12709_, _12702_);
  and (_12711_, _12710_, _01969_);
  and (_12712_, _04129_, \oc8051_golden_model_1.ACC [2]);
  nor (_12713_, _12712_, _12702_);
  nor (_12714_, _12713_, _05488_);
  nor (_12715_, _04571_, _12701_);
  or (_12716_, _12715_, _01969_);
  nor (_12717_, _12716_, _12714_);
  or (_12718_, _12717_, _06233_);
  nor (_12719_, _12718_, _12711_);
  nor (_12720_, _12707_, _05487_);
  nor (_12721_, _05184_, _12701_);
  and (_12722_, _08111_, _05184_);
  nor (_12723_, _12722_, _12721_);
  nor (_12724_, _12723_, _02223_);
  nor (_12725_, _12724_, _12720_);
  nand (_12726_, _12725_, _01964_);
  or (_12727_, _12726_, _12719_);
  nand (_12728_, _12713_, _01963_);
  and (_12729_, _12728_, _12727_);
  nor (_12730_, _12729_, _01957_);
  and (_12731_, _08109_, _05184_);
  nor (_12732_, _12731_, _12721_);
  and (_12733_, _12732_, _01957_);
  or (_12734_, _12733_, _01946_);
  nor (_12735_, _12734_, _12730_);
  nor (_12736_, _12721_, _08139_);
  or (_12737_, _12736_, _04885_);
  nor (_12738_, _12737_, _12723_);
  or (_12739_, _12738_, _12735_);
  and (_12740_, _12739_, _01925_);
  nor (_12741_, _08158_, _06519_);
  nor (_12742_, _12721_, _12741_);
  nor (_12743_, _12742_, _01925_);
  or (_12744_, _12743_, _04950_);
  nor (_12745_, _12744_, _12740_);
  nor (_12746_, _12745_, _12708_);
  nor (_12747_, _12746_, _04951_);
  and (_12748_, _04129_, _03564_);
  nor (_12749_, _12702_, _05513_);
  not (_12750_, _12749_);
  nor (_12751_, _12750_, _12748_);
  or (_12752_, _12751_, _01602_);
  nor (_12753_, _12752_, _12747_);
  nor (_12754_, _08216_, _06482_);
  nor (_12755_, _12754_, _12702_);
  nor (_12756_, _12755_, _01923_);
  or (_12757_, _12756_, _02019_);
  nor (_12758_, _12757_, _12753_);
  nor (_12759_, _12758_, _12705_);
  or (_12760_, _12759_, _02018_);
  and (_12761_, _08230_, _04129_);
  or (_12762_, _12761_, _12702_);
  or (_12763_, _12762_, _05049_);
  and (_12764_, _12763_, _02136_);
  and (_12765_, _12764_, _12760_);
  and (_12766_, _08237_, _04129_);
  nor (_12767_, _12766_, _12702_);
  nor (_12768_, _12767_, _02136_);
  nor (_12769_, _12768_, _12765_);
  nor (_12770_, _12769_, _02039_);
  nor (_12771_, _12702_, _05739_);
  not (_12772_, _12771_);
  nor (_12773_, _12704_, _05076_);
  and (_12774_, _12773_, _12772_);
  nor (_12775_, _12774_, _12770_);
  nor (_12776_, _12775_, _02130_);
  or (_12777_, _12771_, _02131_);
  nor (_12778_, _12777_, _12713_);
  or (_12779_, _12778_, _02016_);
  nor (_12780_, _12779_, _12776_);
  nor (_12781_, _08229_, _06482_);
  nor (_12782_, _12781_, _12702_);
  and (_12783_, _12782_, _02016_);
  nor (_12784_, _12783_, _12780_);
  and (_12785_, _12784_, _05474_);
  nor (_12786_, _08236_, _06482_);
  nor (_12787_, _12786_, _12702_);
  nor (_12788_, _12787_, _05474_);
  or (_12789_, _12788_, _12785_);
  and (_12790_, _12789_, _02168_);
  nor (_12791_, _12710_, _02168_);
  or (_12792_, _12791_, _02025_);
  or (_12793_, _12792_, _12790_);
  nand (_12794_, _12732_, _02025_);
  and (_12795_, _12794_, _12793_);
  nor (_12796_, _12795_, _01594_);
  and (_12797_, _08285_, _04129_);
  nor (_12798_, _12797_, _12702_);
  and (_12799_, _12798_, _01594_);
  nor (_12800_, _12799_, _12796_);
  or (_12801_, _12800_, _26506_);
  or (_12802_, _26505_, \oc8051_golden_model_1.SCON [2]);
  and (_12803_, _12802_, _25964_);
  and (_27844_, _12803_, _12801_);
  not (_12804_, \oc8051_golden_model_1.SCON [3]);
  nor (_12805_, _04129_, _12804_);
  and (_12806_, _04129_, _05529_);
  nor (_12807_, _12806_, _12805_);
  and (_12808_, _12807_, _02019_);
  nor (_12809_, _06482_, _03473_);
  nor (_12810_, _12809_, _12805_);
  and (_12811_, _12810_, _04950_);
  nor (_12812_, _08308_, _06519_);
  nor (_12813_, _05184_, _12804_);
  or (_12814_, _12813_, _01925_);
  or (_12815_, _12814_, _12812_);
  nor (_12816_, _08337_, _06482_);
  nor (_12817_, _12816_, _12805_);
  and (_12818_, _12817_, _01969_);
  and (_12819_, _04129_, \oc8051_golden_model_1.ACC [3]);
  nor (_12820_, _12819_, _12805_);
  nor (_12821_, _12820_, _05488_);
  nor (_12822_, _04571_, _12804_);
  or (_12823_, _12822_, _01969_);
  nor (_12824_, _12823_, _12821_);
  or (_12825_, _12824_, _06233_);
  nor (_12826_, _12825_, _12818_);
  nor (_12827_, _12810_, _05487_);
  and (_12828_, _08341_, _05184_);
  nor (_12829_, _12828_, _12813_);
  nor (_12830_, _12829_, _02223_);
  nor (_12831_, _12830_, _12827_);
  nand (_12832_, _12831_, _01964_);
  or (_12833_, _12832_, _12826_);
  nand (_12834_, _12820_, _01963_);
  and (_12835_, _12834_, _12833_);
  and (_12836_, _12835_, _06229_);
  and (_12837_, _08324_, _05184_);
  nor (_12838_, _12837_, _12813_);
  nor (_12839_, _12838_, _06229_);
  or (_12840_, _12839_, _12836_);
  and (_12841_, _12840_, _04885_);
  nor (_12842_, _12813_, _08357_);
  or (_12843_, _12829_, _04885_);
  nor (_12844_, _12843_, _12842_);
  or (_12845_, _12844_, _01924_);
  or (_12846_, _12845_, _12841_);
  and (_12847_, _12846_, _12815_);
  nor (_12848_, _12847_, _04950_);
  nor (_12849_, _12848_, _12811_);
  nor (_12850_, _12849_, _04951_);
  and (_12851_, _04129_, _03516_);
  nor (_12852_, _12805_, _05513_);
  not (_12853_, _12852_);
  nor (_12854_, _12853_, _12851_);
  or (_12855_, _12854_, _01602_);
  nor (_12856_, _12855_, _12850_);
  nor (_12857_, _08425_, _06482_);
  nor (_12858_, _12857_, _12805_);
  nor (_12859_, _12858_, _01923_);
  or (_12860_, _12859_, _02019_);
  nor (_12861_, _12860_, _12856_);
  nor (_12862_, _12861_, _12808_);
  or (_12863_, _12862_, _02018_);
  and (_12864_, _08441_, _04129_);
  or (_12865_, _12864_, _12805_);
  or (_12866_, _12865_, _05049_);
  and (_12867_, _12866_, _02136_);
  and (_12868_, _12867_, _12863_);
  and (_12869_, _08304_, _04129_);
  nor (_12870_, _12869_, _12805_);
  nor (_12871_, _12870_, _02136_);
  nor (_12872_, _12871_, _12868_);
  nor (_12873_, _12872_, _02039_);
  nor (_12874_, _12805_, _05737_);
  not (_12875_, _12874_);
  nor (_12876_, _12807_, _05076_);
  and (_12877_, _12876_, _12875_);
  nor (_12878_, _12877_, _12873_);
  nor (_12879_, _12878_, _02130_);
  or (_12880_, _12874_, _02131_);
  nor (_12881_, _12880_, _12820_);
  or (_12882_, _12881_, _02016_);
  nor (_12883_, _12882_, _12879_);
  nor (_12884_, _08440_, _06482_);
  nor (_12885_, _12884_, _12805_);
  and (_12886_, _12885_, _02016_);
  nor (_12887_, _12886_, _12883_);
  and (_12888_, _12887_, _05474_);
  nor (_12889_, _08303_, _06482_);
  nor (_12890_, _12889_, _12805_);
  nor (_12891_, _12890_, _05474_);
  or (_12892_, _12891_, _12888_);
  and (_12893_, _12892_, _02168_);
  nor (_12894_, _12817_, _02168_);
  or (_12895_, _12894_, _02025_);
  or (_12896_, _12895_, _12893_);
  nand (_12897_, _12838_, _02025_);
  and (_12898_, _12897_, _12896_);
  nor (_12899_, _12898_, _01594_);
  and (_12900_, _08507_, _04129_);
  nor (_12901_, _12900_, _12805_);
  and (_12902_, _12901_, _01594_);
  nor (_12903_, _12902_, _12899_);
  or (_12904_, _12903_, _26506_);
  or (_12905_, _26505_, \oc8051_golden_model_1.SCON [3]);
  and (_12906_, _12905_, _25964_);
  and (_27845_, _12906_, _12904_);
  not (_12907_, \oc8051_golden_model_1.SCON [4]);
  nor (_12908_, _04129_, _12907_);
  and (_12909_, _04129_, _05524_);
  nor (_12910_, _12909_, _12908_);
  and (_12911_, _12910_, _02019_);
  nor (_12912_, _06482_, _04024_);
  nor (_12913_, _12912_, _12908_);
  and (_12914_, _12913_, _04950_);
  nor (_12915_, _05184_, _12907_);
  nor (_12916_, _12915_, _08581_);
  and (_12917_, _08565_, _05184_);
  nor (_12918_, _12917_, _12915_);
  or (_12919_, _12918_, _04885_);
  nor (_12920_, _12919_, _12916_);
  nor (_12921_, _08548_, _06482_);
  nor (_12922_, _12921_, _12908_);
  and (_12923_, _12922_, _01969_);
  and (_12924_, _04129_, \oc8051_golden_model_1.ACC [4]);
  nor (_12925_, _12924_, _12908_);
  nor (_12926_, _12925_, _05488_);
  nor (_12927_, _04571_, _12907_);
  or (_12928_, _12927_, _01969_);
  nor (_12929_, _12928_, _12926_);
  or (_12930_, _12929_, _06233_);
  nor (_12931_, _12930_, _12923_);
  nor (_12932_, _12913_, _05487_);
  nor (_12933_, _12918_, _02223_);
  nor (_12934_, _12933_, _12932_);
  nand (_12935_, _12934_, _01964_);
  or (_12936_, _12935_, _12931_);
  nand (_12937_, _12925_, _01963_);
  and (_12938_, _12937_, _12936_);
  and (_12939_, _12938_, _06229_);
  and (_12940_, _08544_, _05184_);
  nor (_12941_, _12940_, _12915_);
  nor (_12942_, _12941_, _06229_);
  or (_12943_, _12942_, _12939_);
  and (_12944_, _12943_, _04885_);
  nor (_12945_, _12944_, _12920_);
  nor (_12946_, _12945_, _01924_);
  nor (_12947_, _08607_, _06519_);
  nor (_12948_, _12947_, _12915_);
  nor (_12949_, _12948_, _01925_);
  nor (_12950_, _12949_, _04950_);
  not (_12951_, _12950_);
  nor (_12952_, _12951_, _12946_);
  nor (_12953_, _12952_, _12914_);
  nor (_12954_, _12953_, _04951_);
  and (_12955_, _04129_, _03903_);
  nor (_12956_, _12908_, _05513_);
  not (_12957_, _12956_);
  nor (_12958_, _12957_, _12955_);
  or (_12959_, _12958_, _01602_);
  nor (_12960_, _12959_, _12954_);
  nor (_12961_, _08663_, _06482_);
  nor (_12962_, _12961_, _12908_);
  nor (_12963_, _12962_, _01923_);
  or (_12964_, _12963_, _02019_);
  nor (_12965_, _12964_, _12960_);
  nor (_12966_, _12965_, _12911_);
  or (_12967_, _12966_, _02018_);
  and (_12968_, _08531_, _04129_);
  or (_12969_, _12968_, _12908_);
  or (_12970_, _12969_, _05049_);
  and (_12971_, _12970_, _02136_);
  and (_12972_, _12971_, _12967_);
  and (_12973_, _08527_, _04129_);
  nor (_12974_, _12973_, _12908_);
  nor (_12975_, _12974_, _02136_);
  nor (_12976_, _12975_, _12972_);
  nor (_12977_, _12976_, _02039_);
  nor (_12978_, _12908_, _08729_);
  not (_12979_, _12978_);
  nor (_12980_, _12910_, _05076_);
  and (_12981_, _12980_, _12979_);
  nor (_12982_, _12981_, _12977_);
  nor (_12983_, _12982_, _02130_);
  or (_12984_, _12978_, _02131_);
  nor (_12985_, _12984_, _12925_);
  or (_12986_, _12985_, _02016_);
  nor (_12987_, _12986_, _12983_);
  nor (_12988_, _08530_, _06482_);
  nor (_12989_, _12988_, _12908_);
  and (_12990_, _12989_, _02016_);
  nor (_12991_, _12990_, _12987_);
  and (_12992_, _12991_, _05474_);
  nor (_12993_, _08526_, _06482_);
  nor (_12994_, _12993_, _12908_);
  nor (_12995_, _12994_, _05474_);
  or (_12996_, _12995_, _12992_);
  and (_12997_, _12996_, _02168_);
  nor (_12998_, _12922_, _02168_);
  or (_12999_, _12998_, _02025_);
  or (_13000_, _12999_, _12997_);
  nand (_13001_, _12941_, _02025_);
  and (_13002_, _13001_, _13000_);
  nor (_13003_, _13002_, _01594_);
  and (_13004_, _08732_, _04129_);
  nor (_13005_, _13004_, _12908_);
  and (_13006_, _13005_, _01594_);
  nor (_13007_, _13006_, _13003_);
  or (_13008_, _13007_, _26506_);
  or (_13009_, _26505_, \oc8051_golden_model_1.SCON [4]);
  and (_13010_, _13009_, _25964_);
  and (_27848_, _13010_, _13008_);
  not (_13011_, \oc8051_golden_model_1.SCON [5]);
  nor (_13012_, _04129_, _13011_);
  and (_13013_, _04129_, _05548_);
  nor (_13014_, _13013_, _13012_);
  and (_13015_, _13014_, _02019_);
  nor (_13016_, _06482_, _03976_);
  nor (_13017_, _13016_, _13012_);
  and (_13018_, _13017_, _04950_);
  and (_13019_, _04129_, \oc8051_golden_model_1.ACC [5]);
  nor (_13020_, _13019_, _13012_);
  and (_13021_, _13020_, _01963_);
  nor (_13022_, _08771_, _06482_);
  nor (_13023_, _13022_, _13012_);
  and (_13024_, _13023_, _01969_);
  nor (_13025_, _13020_, _05488_);
  nor (_13026_, _04571_, _13011_);
  or (_13027_, _13026_, _01969_);
  nor (_13028_, _13027_, _13025_);
  or (_13029_, _13028_, _06233_);
  nor (_13030_, _13029_, _13024_);
  nor (_13031_, _13017_, _05487_);
  nor (_13032_, _13031_, _13030_);
  nor (_13033_, _05184_, _13011_);
  and (_13034_, _08785_, _05184_);
  nor (_13035_, _13034_, _13033_);
  nor (_13036_, _13035_, _02223_);
  nor (_13037_, _13036_, _01963_);
  and (_13038_, _13037_, _13032_);
  nor (_13039_, _13038_, _13021_);
  and (_13040_, _13039_, _06229_);
  and (_13041_, _08768_, _05184_);
  nor (_13042_, _13041_, _13033_);
  nor (_13043_, _13042_, _06229_);
  or (_13044_, _13043_, _13040_);
  and (_13045_, _13044_, _04885_);
  nor (_13046_, _13033_, _08801_);
  or (_13047_, _13035_, _04885_);
  nor (_13048_, _13047_, _13046_);
  nor (_13049_, _13048_, _13045_);
  nor (_13050_, _13049_, _01924_);
  nor (_13051_, _08754_, _06519_);
  nor (_13052_, _13051_, _13033_);
  nor (_13053_, _13052_, _01925_);
  nor (_13054_, _13053_, _04950_);
  not (_13055_, _13054_);
  nor (_13056_, _13055_, _13050_);
  nor (_13057_, _13056_, _13018_);
  nor (_13058_, _13057_, _04951_);
  and (_13059_, _04129_, _03850_);
  nor (_13060_, _13012_, _05513_);
  not (_13061_, _13060_);
  nor (_13062_, _13061_, _13059_);
  or (_13063_, _13062_, _01602_);
  nor (_13064_, _13063_, _13058_);
  nor (_13065_, _08874_, _06482_);
  nor (_13066_, _13065_, _13012_);
  nor (_13067_, _13066_, _01923_);
  or (_13068_, _13067_, _02019_);
  nor (_13069_, _13068_, _13064_);
  nor (_13070_, _13069_, _13015_);
  or (_13071_, _13070_, _02018_);
  and (_13072_, _08890_, _04129_);
  or (_13073_, _13072_, _13012_);
  or (_13074_, _13073_, _05049_);
  and (_13075_, _13074_, _02136_);
  and (_13076_, _13075_, _13071_);
  and (_13077_, _08750_, _04129_);
  nor (_13078_, _13077_, _13012_);
  nor (_13079_, _13078_, _02136_);
  nor (_13080_, _13079_, _13076_);
  nor (_13081_, _13080_, _02039_);
  nor (_13082_, _13012_, _08946_);
  not (_13083_, _13082_);
  nor (_13084_, _13014_, _05076_);
  and (_13085_, _13084_, _13083_);
  nor (_13086_, _13085_, _13081_);
  nor (_13087_, _13086_, _02130_);
  or (_13088_, _13082_, _02131_);
  nor (_13089_, _13088_, _13020_);
  or (_13090_, _13089_, _02016_);
  nor (_13091_, _13090_, _13087_);
  nor (_13092_, _08889_, _06482_);
  nor (_13093_, _13092_, _13012_);
  and (_13094_, _13093_, _02016_);
  nor (_13095_, _13094_, _13091_);
  and (_13096_, _13095_, _05474_);
  nor (_13097_, _08749_, _06482_);
  nor (_13098_, _13097_, _13012_);
  nor (_13099_, _13098_, _05474_);
  or (_13100_, _13099_, _13096_);
  and (_13101_, _13100_, _02168_);
  nor (_13102_, _13023_, _02168_);
  or (_13103_, _13102_, _02025_);
  or (_13104_, _13103_, _13101_);
  nand (_13105_, _13042_, _02025_);
  and (_13106_, _13105_, _13104_);
  nor (_13107_, _13106_, _01594_);
  and (_13108_, _08949_, _04129_);
  nor (_13109_, _13108_, _13012_);
  and (_13110_, _13109_, _01594_);
  nor (_13111_, _13110_, _13107_);
  or (_13112_, _13111_, _26506_);
  or (_13113_, _26505_, \oc8051_golden_model_1.SCON [5]);
  and (_13114_, _13113_, _25964_);
  and (_27849_, _13114_, _13112_);
  not (_13115_, \oc8051_golden_model_1.SCON [6]);
  nor (_13116_, _04129_, _13115_);
  and (_13117_, _04129_, _03748_);
  or (_13118_, _13117_, _13116_);
  and (_13119_, _13118_, _04951_);
  nor (_13120_, _05184_, _13115_);
  not (_13121_, _13120_);
  and (_13122_, _13121_, _09026_);
  and (_13123_, _09011_, _05184_);
  nor (_13124_, _13123_, _13120_);
  or (_13125_, _13124_, _04885_);
  nor (_13126_, _13125_, _13122_);
  nor (_13127_, _08995_, _06482_);
  nor (_13128_, _13127_, _13116_);
  and (_13129_, _13128_, _01969_);
  and (_13130_, _04129_, \oc8051_golden_model_1.ACC [6]);
  nor (_13131_, _13130_, _13116_);
  nor (_13132_, _13131_, _05488_);
  nor (_13133_, _04571_, _13115_);
  or (_13134_, _13133_, _01969_);
  nor (_13135_, _13134_, _13132_);
  or (_13136_, _13135_, _06233_);
  nor (_13137_, _13136_, _13129_);
  nor (_13138_, _06482_, _04074_);
  nor (_13139_, _13138_, _13116_);
  nor (_13140_, _13139_, _05487_);
  nor (_13141_, _13124_, _02223_);
  nor (_13142_, _13141_, _13140_);
  nand (_13143_, _13142_, _01964_);
  or (_13144_, _13143_, _13137_);
  nand (_13145_, _13131_, _01963_);
  and (_13146_, _13145_, _13144_);
  and (_13147_, _13146_, _06229_);
  and (_13148_, _08992_, _05184_);
  nor (_13149_, _13148_, _13120_);
  nor (_13150_, _13149_, _06229_);
  or (_13151_, _13150_, _13147_);
  and (_13152_, _13151_, _04885_);
  nor (_13153_, _13152_, _13126_);
  nor (_13154_, _13153_, _01924_);
  nor (_13155_, _08979_, _06519_);
  nor (_13156_, _13155_, _13120_);
  nor (_13157_, _13156_, _01925_);
  nor (_13158_, _13157_, _04950_);
  not (_13159_, _13158_);
  nor (_13160_, _13159_, _13154_);
  and (_13161_, _13139_, _04950_);
  or (_13162_, _13161_, _04951_);
  nor (_13163_, _13162_, _13160_);
  or (_13164_, _13163_, _13119_);
  and (_13165_, _13164_, _01923_);
  nor (_13166_, _09096_, _06482_);
  nor (_13167_, _13166_, _13116_);
  nor (_13168_, _13167_, _01923_);
  or (_13169_, _13168_, _06278_);
  or (_13170_, _13169_, _13165_);
  and (_13171_, _09112_, _04129_);
  or (_13172_, _13116_, _05049_);
  or (_13173_, _13172_, _13171_);
  and (_13174_, _04129_, _09103_);
  nor (_13175_, _13174_, _13116_);
  and (_13176_, _13175_, _02019_);
  nor (_13177_, _13176_, _02135_);
  and (_13178_, _13177_, _13173_);
  and (_13179_, _13178_, _13170_);
  and (_13180_, _08975_, _04129_);
  nor (_13181_, _13180_, _13116_);
  nor (_13182_, _13181_, _02136_);
  nor (_13183_, _13182_, _13179_);
  nor (_13184_, _13183_, _02039_);
  nor (_13185_, _13116_, _05735_);
  not (_13186_, _13185_);
  nor (_13187_, _13175_, _05076_);
  and (_13188_, _13187_, _13186_);
  nor (_13189_, _13188_, _13184_);
  nor (_13190_, _13189_, _02130_);
  or (_13191_, _13185_, _02131_);
  nor (_13192_, _13191_, _13131_);
  or (_13193_, _13192_, _02016_);
  nor (_13194_, _13193_, _13190_);
  nor (_13195_, _09111_, _06482_);
  nor (_13196_, _13195_, _13116_);
  and (_13197_, _13196_, _02016_);
  nor (_13198_, _13197_, _13194_);
  and (_13199_, _13198_, _05474_);
  nor (_13200_, _08974_, _06482_);
  nor (_13201_, _13200_, _13116_);
  nor (_13202_, _13201_, _05474_);
  or (_13203_, _13202_, _13199_);
  and (_13204_, _13203_, _02168_);
  nor (_13205_, _13128_, _02168_);
  or (_13206_, _13205_, _02025_);
  or (_13207_, _13206_, _13204_);
  nand (_13208_, _13149_, _02025_);
  and (_13209_, _13208_, _13207_);
  nor (_13210_, _13209_, _01594_);
  and (_13211_, _08965_, _04129_);
  nor (_13212_, _13211_, _13116_);
  and (_13213_, _13212_, _01594_);
  nor (_13214_, _13213_, _13210_);
  or (_13215_, _13214_, _26506_);
  or (_13216_, _26505_, \oc8051_golden_model_1.SCON [6]);
  and (_13217_, _13216_, _25964_);
  and (_27850_, _13217_, _13215_);
  nor (_13218_, _04111_, _02441_);
  nor (_13219_, _04405_, _06336_);
  or (_13220_, _13219_, _13218_);
  or (_13221_, _13220_, _02438_);
  and (_13222_, _04396_, \oc8051_golden_model_1.ACC [0]);
  or (_13223_, _13222_, _13218_);
  and (_13224_, _13223_, _04571_);
  nor (_13225_, _04571_, _02441_);
  or (_13226_, _13225_, _01969_);
  or (_13227_, _13226_, _13224_);
  and (_13228_, _13227_, _05487_);
  and (_13229_, _13228_, _13221_);
  or (_13230_, _13229_, _02443_);
  or (_13231_, _13223_, _01964_);
  and (_13232_, _13231_, _02457_);
  and (_13233_, _13232_, _13230_);
  or (_13234_, _06978_, _04950_);
  or (_13235_, _13234_, _13233_);
  and (_13236_, _04111_, _03334_);
  or (_13237_, _13218_, _06397_);
  or (_13238_, _13237_, _13236_);
  and (_13239_, _13238_, _13235_);
  or (_13240_, _13239_, _04951_);
  or (_13241_, _13218_, _05513_);
  and (_13242_, _04396_, _03677_);
  or (_13243_, _13242_, _13241_);
  and (_13244_, _13243_, _13240_);
  or (_13245_, _13244_, _01602_);
  nor (_13246_, _07815_, _06442_);
  or (_13247_, _13246_, _13218_);
  or (_13248_, _13247_, _01923_);
  and (_13249_, _13248_, _04979_);
  and (_13250_, _13249_, _13245_);
  and (_13251_, _04396_, _05531_);
  or (_13252_, _13251_, _13218_);
  and (_13253_, _13252_, _02019_);
  or (_13254_, _13253_, _02018_);
  or (_13255_, _13254_, _13250_);
  and (_13256_, _07829_, _04396_);
  or (_13257_, _13256_, _13218_);
  or (_13258_, _13257_, _05049_);
  and (_13259_, _13258_, _13255_);
  or (_13260_, _13259_, _02135_);
  and (_13261_, _07834_, _04111_);
  or (_13262_, _13218_, _02136_);
  or (_13263_, _13262_, _13261_);
  and (_13264_, _13263_, _05076_);
  and (_13265_, _13264_, _13260_);
  nand (_13266_, _13252_, _02039_);
  nor (_13267_, _13266_, _13219_);
  or (_13268_, _13267_, _13265_);
  and (_13269_, _13268_, _02131_);
  or (_13270_, _13218_, _04405_);
  and (_13271_, _13223_, _02130_);
  and (_13272_, _13271_, _13270_);
  or (_13273_, _13272_, _02016_);
  or (_13274_, _13273_, _13269_);
  nor (_13275_, _07828_, _06336_);
  or (_13276_, _13218_, _05104_);
  or (_13277_, _13276_, _13275_);
  and (_13278_, _13277_, _05474_);
  and (_13279_, _13278_, _13274_);
  nor (_13280_, _07696_, _06336_);
  or (_13281_, _13280_, _13218_);
  and (_13282_, _13281_, _02126_);
  or (_13283_, _13282_, _02266_);
  or (_13284_, _13283_, _13279_);
  or (_13285_, _13220_, _02265_);
  and (_13286_, _13285_, _26505_);
  and (_13287_, _13286_, _13284_);
  nor (_13288_, _26505_, _02441_);
  or (_13289_, _13288_, rst);
  or (_27852_, _13289_, _13287_);
  nor (_13290_, _04111_, _02717_);
  and (_13291_, _07909_, _04111_);
  or (_13292_, _13291_, _13290_);
  and (_13293_, _13292_, _01594_);
  nand (_13294_, _02146_, \oc8051_golden_model_1.SP [1]);
  or (_13295_, _08029_, _06336_);
  or (_13296_, _04111_, \oc8051_golden_model_1.SP [1]);
  and (_13297_, _13296_, _02135_);
  and (_13298_, _13297_, _13295_);
  not (_13299_, _13291_);
  and (_13300_, _13296_, _13299_);
  or (_13301_, _13300_, _02438_);
  or (_13302_, _01625_, _02717_);
  nand (_13303_, _04111_, _01705_);
  and (_13304_, _13303_, _13296_);
  and (_13305_, _13304_, _04571_);
  nor (_13306_, _04571_, _02717_);
  or (_13307_, _13306_, _04568_);
  or (_13308_, _13307_, _13305_);
  and (_13309_, _13308_, _13302_);
  or (_13310_, _13309_, _01969_);
  and (_13311_, _13310_, _01621_);
  and (_13312_, _13311_, _13301_);
  nor (_13313_, _01621_, \oc8051_golden_model_1.SP [1]);
  or (_13314_, _13313_, _01967_);
  or (_13315_, _13314_, _13312_);
  nand (_13316_, _03400_, _01967_);
  and (_13317_, _13316_, _13315_);
  or (_13318_, _13317_, _01963_);
  or (_13319_, _13304_, _01964_);
  and (_13320_, _13319_, _02457_);
  and (_13321_, _13320_, _13318_);
  not (_13322_, _06394_);
  or (_13323_, _07210_, _13322_);
  or (_13324_, _13323_, _13321_);
  or (_13325_, _06394_, _02717_);
  and (_13326_, _13325_, _06397_);
  and (_13327_, _13326_, _13324_);
  nand (_13328_, _04111_, _03393_);
  and (_13329_, _13296_, _04950_);
  and (_13330_, _13329_, _13328_);
  or (_13331_, _13330_, _04951_);
  or (_13332_, _13331_, _13327_);
  or (_13333_, _13290_, _05513_);
  and (_13334_, _04396_, _03613_);
  or (_13335_, _13334_, _13333_);
  and (_13336_, _13335_, _01923_);
  and (_13337_, _13336_, _13332_);
  and (_13338_, _13296_, _01602_);
  nand (_13339_, _08009_, _04111_);
  and (_13340_, _13339_, _13338_);
  or (_13341_, _13340_, _13337_);
  and (_13342_, _13341_, _04979_);
  and (_13343_, _13296_, _02019_);
  nand (_13344_, _04396_, _02676_);
  and (_13345_, _13344_, _13343_);
  or (_13346_, _13345_, _01650_);
  or (_13347_, _13346_, _13342_);
  nand (_13348_, _01650_, \oc8051_golden_model_1.SP [1]);
  and (_13349_, _13348_, _05049_);
  and (_13350_, _13349_, _13347_);
  or (_13351_, _08023_, _06336_);
  and (_13352_, _13296_, _02018_);
  and (_13353_, _13352_, _13351_);
  or (_13354_, _13353_, _13350_);
  and (_13355_, _13354_, _02136_);
  or (_13356_, _13355_, _13298_);
  and (_13357_, _13356_, _05076_);
  or (_13358_, _07893_, _06336_);
  and (_13359_, _13296_, _02039_);
  and (_13360_, _13359_, _13358_);
  or (_13361_, _13360_, _13357_);
  and (_13362_, _13361_, _05082_);
  and (_13363_, _01666_, _02717_);
  or (_13364_, _13290_, _05741_);
  and (_13365_, _13304_, _02130_);
  and (_13366_, _13365_, _13364_);
  or (_13367_, _13366_, _13363_);
  or (_13368_, _13367_, _13362_);
  and (_13369_, _13368_, _02127_);
  or (_13370_, _13303_, _05741_);
  and (_13371_, _13370_, _02126_);
  and (_13372_, _13371_, _13296_);
  or (_13373_, _13372_, _02146_);
  or (_13374_, _13344_, _05741_);
  and (_13375_, _13374_, _02016_);
  and (_13376_, _13375_, _13296_);
  or (_13377_, _13376_, _13373_);
  or (_13378_, _13377_, _13369_);
  nand (_13379_, _13378_, _13294_);
  nor (_13380_, _01660_, _01585_);
  nand (_13381_, _13380_, _13379_);
  or (_13382_, _13380_, _02717_);
  and (_13383_, _13382_, _02168_);
  and (_13384_, _13383_, _13381_);
  and (_13385_, _13300_, _02164_);
  or (_13386_, _13385_, _06467_);
  or (_13387_, _13386_, _13384_);
  or (_13388_, _06466_, _02717_);
  and (_13389_, _13388_, _01595_);
  and (_13390_, _13389_, _13387_);
  or (_13391_, _13390_, _13293_);
  and (_13392_, _13391_, _26505_);
  nor (_13393_, _26505_, _02717_);
  or (_13394_, _13393_, rst);
  or (_27853_, _13394_, _13392_);
  nor (_13395_, _26505_, _02334_);
  or (_13396_, _13395_, rst);
  nor (_13397_, _04111_, _02334_);
  and (_13398_, _08237_, _04111_);
  or (_13399_, _13398_, _13397_);
  and (_13400_, _13399_, _02135_);
  nand (_13401_, _09521_, _01650_);
  nor (_13402_, _06336_, _03272_);
  or (_13403_, _13397_, _06397_);
  or (_13404_, _13403_, _13402_);
  nor (_13405_, _08095_, _06336_);
  or (_13406_, _13405_, _13397_);
  or (_13407_, _13406_, _02438_);
  and (_13408_, _04396_, \oc8051_golden_model_1.ACC [2]);
  or (_13409_, _13408_, _13397_);
  or (_13410_, _13409_, _05488_);
  or (_13411_, _04571_, \oc8051_golden_model_1.SP [2]);
  and (_13412_, _13411_, _01625_);
  and (_13413_, _13412_, _13410_);
  nor (_13414_, _09521_, _01625_);
  or (_13415_, _13414_, _01969_);
  or (_13416_, _13415_, _13413_);
  and (_13417_, _13416_, _01621_);
  and (_13418_, _13417_, _13407_);
  nor (_13419_, _09521_, _01621_);
  or (_13420_, _13419_, _01967_);
  or (_13421_, _13420_, _13418_);
  nand (_13422_, _03195_, _01967_);
  and (_13423_, _13422_, _13421_);
  or (_13424_, _13423_, _01963_);
  or (_13425_, _13409_, _01964_);
  and (_13426_, _13425_, _02457_);
  and (_13427_, _13426_, _13424_);
  or (_13428_, _13427_, _07415_);
  and (_13429_, _13428_, _06394_);
  nor (_13430_, _09521_, _06394_);
  or (_13431_, _13430_, _04950_);
  or (_13432_, _13431_, _13429_);
  and (_13433_, _13432_, _13404_);
  or (_13434_, _13433_, _04951_);
  or (_13435_, _13397_, _05513_);
  and (_13436_, _04396_, _03564_);
  or (_13437_, _13436_, _13435_);
  and (_13438_, _13437_, _01923_);
  and (_13439_, _13438_, _13434_);
  nor (_13440_, _08216_, _06442_);
  or (_13441_, _13440_, _13397_);
  and (_13442_, _13441_, _01602_);
  or (_13443_, _13442_, _02019_);
  or (_13444_, _13443_, _13439_);
  and (_13445_, _04396_, _05563_);
  or (_13446_, _13445_, _13397_);
  or (_13447_, _13446_, _04979_);
  and (_13448_, _13447_, _13444_);
  or (_13449_, _13448_, _01650_);
  and (_13450_, _13449_, _13401_);
  or (_13451_, _13450_, _02018_);
  and (_13452_, _08230_, _04111_);
  or (_13453_, _13397_, _05049_);
  or (_13454_, _13453_, _13452_);
  and (_13455_, _13454_, _02136_);
  and (_13456_, _13455_, _13451_);
  or (_13457_, _13456_, _13400_);
  and (_13458_, _13457_, _05076_);
  or (_13459_, _13397_, _05739_);
  and (_13460_, _13446_, _02039_);
  and (_13461_, _13460_, _13459_);
  or (_13462_, _13461_, _13458_);
  and (_13463_, _13462_, _05082_);
  and (_13464_, _07481_, _01666_);
  or (_13465_, _13464_, _02016_);
  and (_13466_, _13409_, _02130_);
  and (_13467_, _13466_, _13459_);
  or (_13468_, _13467_, _13465_);
  or (_13469_, _13468_, _13463_);
  nor (_13470_, _08229_, _06442_);
  or (_13471_, _13470_, _13397_);
  or (_13472_, _13471_, _05104_);
  and (_13473_, _13472_, _13469_);
  or (_13474_, _13473_, _02126_);
  nor (_13475_, _08236_, _06336_);
  or (_13476_, _13397_, _05474_);
  or (_13477_, _13476_, _13475_);
  and (_13478_, _13477_, _02718_);
  and (_13479_, _13478_, _13474_);
  and (_13480_, _09521_, _02146_);
  or (_13481_, _13480_, _01660_);
  or (_13482_, _13481_, _13479_);
  nand (_13483_, _09521_, _01660_);
  and (_13484_, _13483_, _01596_);
  and (_13485_, _13484_, _13482_);
  and (_13486_, _09521_, _01585_);
  or (_13487_, _13486_, _02164_);
  or (_13488_, _13487_, _13485_);
  or (_13489_, _13406_, _02168_);
  and (_13490_, _13489_, _06466_);
  and (_13491_, _13490_, _13488_);
  nor (_13492_, _09521_, _06466_);
  or (_13493_, _13492_, _01594_);
  or (_13494_, _13493_, _13491_);
  and (_13495_, _08285_, _04111_);
  or (_13496_, _13397_, _01595_);
  or (_13497_, _13496_, _13495_);
  and (_13498_, _13497_, _26505_);
  and (_13499_, _13498_, _13494_);
  or (_27854_, _13499_, _13396_);
  nor (_13500_, _26505_, _02160_);
  or (_13501_, _07484_, _06466_);
  nor (_13502_, _04111_, _02160_);
  and (_13503_, _08304_, _04111_);
  or (_13504_, _13503_, _13502_);
  and (_13505_, _13504_, _02135_);
  nand (_13506_, _09338_, _01650_);
  nor (_13507_, _06336_, _03473_);
  or (_13508_, _13502_, _04951_);
  or (_13509_, _13508_, _13507_);
  and (_13510_, _13509_, _04953_);
  nor (_13511_, _08337_, _06336_);
  or (_13512_, _13511_, _13502_);
  or (_13513_, _13512_, _02438_);
  and (_13514_, _04396_, \oc8051_golden_model_1.ACC [3]);
  or (_13515_, _13514_, _13502_);
  and (_13516_, _13515_, _04571_);
  nor (_13517_, _04571_, _02160_);
  or (_13518_, _13517_, _04568_);
  or (_13519_, _13518_, _13516_);
  or (_13520_, _07484_, _01625_);
  and (_13521_, _13520_, _13519_);
  or (_13522_, _13521_, _01969_);
  and (_13523_, _13522_, _01621_);
  and (_13524_, _13523_, _13513_);
  nor (_13525_, _09338_, _01621_);
  or (_13526_, _13525_, _01967_);
  or (_13527_, _13526_, _13524_);
  nand (_13528_, _03420_, _01967_);
  and (_13529_, _13528_, _13527_);
  or (_13530_, _13529_, _01963_);
  or (_13531_, _13515_, _01964_);
  and (_13532_, _13531_, _02457_);
  and (_13533_, _13532_, _13530_);
  or (_13534_, _07314_, _13322_);
  or (_13535_, _13534_, _13533_);
  or (_13536_, _07484_, _06394_);
  and (_13537_, _13536_, _06397_);
  and (_13538_, _13537_, _13535_);
  or (_13539_, _13538_, _13510_);
  or (_13540_, _13502_, _05513_);
  and (_13541_, _04396_, _03516_);
  or (_13542_, _13541_, _13540_);
  and (_13543_, _13542_, _01923_);
  and (_13544_, _13543_, _13539_);
  nor (_13545_, _08425_, _06442_);
  or (_13546_, _13545_, _13502_);
  and (_13547_, _13546_, _01602_);
  or (_13548_, _13547_, _02019_);
  or (_13549_, _13548_, _13544_);
  and (_13550_, _04396_, _05529_);
  or (_13551_, _13550_, _13502_);
  or (_13552_, _13551_, _04979_);
  and (_13553_, _13552_, _13549_);
  or (_13554_, _13553_, _01650_);
  and (_13555_, _13554_, _13506_);
  or (_13556_, _13555_, _02018_);
  and (_13557_, _08441_, _04111_);
  or (_13558_, _13502_, _05049_);
  or (_13559_, _13558_, _13557_);
  and (_13560_, _13559_, _02136_);
  and (_13561_, _13560_, _13556_);
  or (_13562_, _13561_, _13505_);
  and (_13563_, _13562_, _05076_);
  or (_13564_, _13502_, _05737_);
  and (_13565_, _13551_, _02039_);
  and (_13566_, _13565_, _13564_);
  or (_13567_, _13566_, _13563_);
  and (_13568_, _13567_, _05082_);
  and (_13569_, _13515_, _02130_);
  and (_13570_, _13569_, _13564_);
  and (_13571_, _07484_, _01666_);
  or (_13572_, _13571_, _02016_);
  or (_13573_, _13572_, _13570_);
  or (_13574_, _13573_, _13568_);
  nor (_13575_, _08440_, _06442_);
  or (_13576_, _13575_, _13502_);
  or (_13577_, _13576_, _05104_);
  and (_13578_, _13577_, _13574_);
  or (_13579_, _13578_, _02126_);
  nor (_13580_, _08303_, _06336_);
  or (_13581_, _13502_, _05474_);
  or (_13582_, _13581_, _13580_);
  and (_13583_, _13582_, _02718_);
  and (_13584_, _13583_, _13579_);
  nor (_13585_, _03417_, _02160_);
  or (_13586_, _13585_, _03418_);
  and (_13587_, _13586_, _02146_);
  or (_13588_, _13587_, _01660_);
  or (_13589_, _13588_, _13584_);
  nand (_13590_, _09338_, _01660_);
  and (_13591_, _13590_, _13589_);
  or (_13592_, _13591_, _01585_);
  or (_13593_, _13586_, _01596_);
  and (_13594_, _13593_, _02168_);
  and (_13595_, _13594_, _13592_);
  and (_13596_, _13512_, _02164_);
  or (_13597_, _13596_, _06467_);
  or (_13598_, _13597_, _13595_);
  and (_13599_, _13598_, _13501_);
  or (_13600_, _13599_, _01594_);
  and (_13601_, _08507_, _04111_);
  or (_13602_, _13502_, _01595_);
  or (_13603_, _13602_, _13601_);
  and (_13604_, _13603_, _26505_);
  and (_13605_, _13604_, _13600_);
  or (_13606_, _13605_, _13500_);
  and (_27855_, _13606_, _25964_);
  nor (_13607_, _04111_, _06369_);
  and (_13608_, _08527_, _04111_);
  or (_13609_, _13608_, _13607_);
  and (_13610_, _13609_, _02135_);
  nor (_13611_, _06336_, _04024_);
  or (_13612_, _13607_, _04951_);
  or (_13613_, _13612_, _13611_);
  and (_13614_, _13613_, _04953_);
  nor (_13615_, _08548_, _06336_);
  or (_13616_, _13615_, _13607_);
  or (_13617_, _13616_, _02438_);
  and (_13618_, _04396_, \oc8051_golden_model_1.ACC [4]);
  or (_13619_, _13618_, _13607_);
  and (_13620_, _13619_, _04571_);
  nor (_13621_, _04571_, _06369_);
  or (_13622_, _13621_, _04568_);
  or (_13623_, _13622_, _13620_);
  nor (_13624_, _06351_, \oc8051_golden_model_1.SP [4]);
  nor (_13625_, _13624_, _06352_);
  or (_13626_, _13625_, _01625_);
  and (_13627_, _13626_, _13623_);
  or (_13628_, _13627_, _01969_);
  and (_13629_, _13628_, _01621_);
  and (_13630_, _13629_, _13617_);
  and (_13631_, _13625_, _06363_);
  or (_13632_, _13631_, _01967_);
  or (_13633_, _13632_, _13630_);
  and (_13634_, _06370_, _02441_);
  nor (_13635_, _03419_, _06369_);
  nor (_13636_, _13635_, _13634_);
  nand (_13637_, _13636_, _01967_);
  and (_13638_, _13637_, _13633_);
  or (_13639_, _13638_, _01963_);
  or (_13640_, _13619_, _01964_);
  and (_13641_, _13640_, _02457_);
  and (_13642_, _13641_, _13639_);
  nor (_13643_, _06384_, \oc8051_golden_model_1.SP [4]);
  nor (_13644_, _13643_, _06385_);
  nand (_13645_, _13644_, _01953_);
  nand (_13646_, _13645_, _06394_);
  or (_13647_, _13646_, _13642_);
  or (_13648_, _13625_, _06394_);
  and (_13649_, _13648_, _06397_);
  and (_13650_, _13649_, _13647_);
  or (_13651_, _13650_, _13614_);
  or (_13652_, _13607_, _05513_);
  and (_13653_, _04396_, _03903_);
  or (_13654_, _13653_, _13652_);
  and (_13655_, _13654_, _01923_);
  and (_13656_, _13655_, _13651_);
  nor (_13657_, _08663_, _06442_);
  or (_13658_, _13657_, _13607_);
  and (_13659_, _13658_, _01602_);
  or (_13660_, _13659_, _02019_);
  or (_13661_, _13660_, _13656_);
  and (_13662_, _04396_, _05524_);
  or (_13663_, _13662_, _13607_);
  or (_13664_, _13663_, _04979_);
  and (_13665_, _13664_, _13661_);
  or (_13666_, _13665_, _01650_);
  or (_13667_, _13625_, _01651_);
  and (_13668_, _13667_, _13666_);
  or (_13669_, _13668_, _02018_);
  and (_13670_, _08531_, _04111_);
  or (_13671_, _13607_, _05049_);
  or (_13672_, _13671_, _13670_);
  and (_13673_, _13672_, _02136_);
  and (_13674_, _13673_, _13669_);
  or (_13675_, _13674_, _13610_);
  and (_13676_, _13675_, _05076_);
  or (_13677_, _13607_, _08729_);
  and (_13678_, _13663_, _02039_);
  and (_13679_, _13678_, _13677_);
  or (_13680_, _13679_, _13676_);
  and (_13681_, _13680_, _05082_);
  and (_13682_, _13625_, _01666_);
  or (_13683_, _13682_, _02016_);
  and (_13684_, _13619_, _02130_);
  and (_13685_, _13684_, _13677_);
  or (_13686_, _13685_, _13683_);
  or (_13687_, _13686_, _13681_);
  nor (_13688_, _08530_, _06442_);
  or (_13689_, _13688_, _13607_);
  or (_13690_, _13689_, _05104_);
  and (_13691_, _13690_, _13687_);
  or (_13692_, _13691_, _02126_);
  nor (_13693_, _08526_, _06336_);
  or (_13694_, _13607_, _05474_);
  or (_13695_, _13694_, _13693_);
  and (_13696_, _13695_, _02718_);
  and (_13697_, _13696_, _13692_);
  nor (_13698_, _03418_, _06369_);
  or (_13699_, _13698_, _06370_);
  and (_13700_, _13699_, _02146_);
  or (_13701_, _13700_, _01660_);
  or (_13702_, _13701_, _13697_);
  or (_13703_, _13625_, _05157_);
  and (_13704_, _13703_, _13702_);
  or (_13705_, _13704_, _01585_);
  or (_13706_, _13699_, _01596_);
  and (_13707_, _13706_, _02168_);
  and (_13708_, _13707_, _13705_);
  and (_13709_, _13616_, _02164_);
  or (_13710_, _13709_, _06467_);
  or (_13711_, _13710_, _13708_);
  or (_13712_, _13625_, _06466_);
  and (_13713_, _13712_, _01595_);
  and (_13714_, _13713_, _13711_);
  and (_13715_, _08732_, _04111_);
  or (_13716_, _13715_, _13607_);
  and (_13717_, _13716_, _01594_);
  or (_13718_, _13717_, _26506_);
  or (_13719_, _13718_, _13714_);
  or (_13720_, _26505_, \oc8051_golden_model_1.SP [4]);
  and (_13721_, _13720_, _25964_);
  and (_27856_, _13721_, _13719_);
  nor (_13722_, _04111_, _06368_);
  and (_13723_, _08750_, _04111_);
  or (_13724_, _13723_, _13722_);
  and (_13725_, _13724_, _02135_);
  nor (_13726_, _06336_, _03976_);
  or (_13727_, _13722_, _04951_);
  or (_13728_, _13727_, _13726_);
  and (_13729_, _13728_, _04953_);
  nor (_13730_, _08771_, _06336_);
  or (_13731_, _13730_, _13722_);
  or (_13732_, _13731_, _02438_);
  and (_13733_, _04396_, \oc8051_golden_model_1.ACC [5]);
  or (_13734_, _13733_, _13722_);
  and (_13735_, _13734_, _04571_);
  nor (_13736_, _04571_, _06368_);
  or (_13737_, _13736_, _04568_);
  or (_13738_, _13737_, _13735_);
  nor (_13739_, _06352_, \oc8051_golden_model_1.SP [5]);
  nor (_13740_, _13739_, _06353_);
  or (_13741_, _13740_, _01625_);
  and (_13742_, _13741_, _13738_);
  or (_13743_, _13742_, _01969_);
  and (_13744_, _13743_, _13732_);
  and (_13745_, _13744_, _01621_);
  and (_13746_, _13740_, _06363_);
  or (_13747_, _13746_, _01967_);
  or (_13748_, _13747_, _13745_);
  and (_13749_, _06371_, _02441_);
  nor (_13750_, _13634_, _06368_);
  nor (_13751_, _13750_, _13749_);
  nand (_13752_, _13751_, _01967_);
  and (_13753_, _13752_, _13748_);
  or (_13754_, _13753_, _01963_);
  or (_13755_, _13734_, _01964_);
  and (_13756_, _13755_, _02457_);
  and (_13757_, _13756_, _13754_);
  nor (_13758_, _06385_, \oc8051_golden_model_1.SP [5]);
  nor (_13759_, _13758_, _06386_);
  nand (_13760_, _13759_, _01953_);
  nand (_13761_, _13760_, _06394_);
  or (_13762_, _13761_, _13757_);
  or (_13763_, _13740_, _06394_);
  and (_13764_, _13763_, _06397_);
  and (_13765_, _13764_, _13762_);
  or (_13766_, _13765_, _13729_);
  or (_13767_, _13722_, _05513_);
  and (_13768_, _04396_, _03850_);
  or (_13769_, _13768_, _13767_);
  and (_13770_, _13769_, _01923_);
  and (_13771_, _13770_, _13766_);
  nor (_13772_, _08874_, _06442_);
  or (_13773_, _13772_, _13722_);
  and (_13774_, _13773_, _01602_);
  or (_13775_, _13774_, _02019_);
  or (_13776_, _13775_, _13771_);
  and (_13777_, _04396_, _05548_);
  or (_13778_, _13777_, _13722_);
  or (_13779_, _13778_, _04979_);
  and (_13780_, _13779_, _13776_);
  or (_13781_, _13780_, _01650_);
  or (_13782_, _13740_, _01651_);
  and (_13783_, _13782_, _13781_);
  or (_13784_, _13783_, _02018_);
  and (_13785_, _08890_, _04111_);
  or (_13786_, _13722_, _05049_);
  or (_13787_, _13786_, _13785_);
  and (_13788_, _13787_, _02136_);
  and (_13789_, _13788_, _13784_);
  or (_13790_, _13789_, _13725_);
  and (_13791_, _13790_, _05076_);
  or (_13792_, _13722_, _08946_);
  and (_13793_, _13778_, _02039_);
  and (_13794_, _13793_, _13792_);
  or (_13795_, _13794_, _13791_);
  and (_13796_, _13795_, _05082_);
  and (_13797_, _13740_, _01666_);
  or (_13798_, _13797_, _02016_);
  and (_13799_, _13734_, _02130_);
  and (_13800_, _13799_, _13792_);
  or (_13801_, _13800_, _13798_);
  or (_13802_, _13801_, _13796_);
  nor (_13803_, _08889_, _06442_);
  or (_13804_, _13803_, _13722_);
  or (_13805_, _13804_, _05104_);
  and (_13806_, _13805_, _13802_);
  or (_13807_, _13806_, _02126_);
  nor (_13808_, _08749_, _06336_);
  or (_13809_, _13722_, _05474_);
  or (_13810_, _13809_, _13808_);
  and (_13811_, _13810_, _02718_);
  and (_13812_, _13811_, _13807_);
  nor (_13813_, _06370_, _06368_);
  or (_13814_, _13813_, _06371_);
  and (_13815_, _13814_, _02146_);
  or (_13816_, _13815_, _01660_);
  or (_13817_, _13816_, _13812_);
  or (_13818_, _13740_, _05157_);
  and (_13819_, _13818_, _13817_);
  or (_13820_, _13819_, _01585_);
  or (_13821_, _13814_, _01596_);
  and (_13822_, _13821_, _02168_);
  and (_13823_, _13822_, _13820_);
  and (_13824_, _13731_, _02164_);
  or (_13825_, _13824_, _06467_);
  or (_13826_, _13825_, _13823_);
  or (_13827_, _13740_, _06466_);
  and (_13828_, _13827_, _01595_);
  and (_13829_, _13828_, _13826_);
  and (_13830_, _08949_, _04111_);
  or (_13831_, _13830_, _13722_);
  and (_13832_, _13831_, _01594_);
  or (_13833_, _13832_, _26506_);
  or (_13834_, _13833_, _13829_);
  or (_13835_, _26505_, \oc8051_golden_model_1.SP [5]);
  and (_13836_, _13835_, _25964_);
  and (_27857_, _13836_, _13834_);
  nor (_13837_, _26505_, _06367_);
  nor (_13838_, _04111_, _06367_);
  and (_13839_, _08975_, _04111_);
  or (_13840_, _13839_, _13838_);
  and (_13841_, _13840_, _02135_);
  nor (_13842_, _08995_, _06336_);
  or (_13843_, _13842_, _13838_);
  or (_13844_, _13843_, _02438_);
  and (_13845_, _04396_, \oc8051_golden_model_1.ACC [6]);
  or (_13846_, _13845_, _13838_);
  or (_13847_, _13846_, _05488_);
  or (_13848_, _04571_, \oc8051_golden_model_1.SP [6]);
  and (_13849_, _13848_, _01625_);
  and (_13850_, _13849_, _13847_);
  nor (_13851_, _06353_, \oc8051_golden_model_1.SP [6]);
  nor (_13852_, _13851_, _06354_);
  and (_13853_, _13852_, _04568_);
  or (_13854_, _13853_, _01969_);
  or (_13855_, _13854_, _13850_);
  and (_13856_, _13855_, _01621_);
  and (_13857_, _13856_, _13844_);
  and (_13858_, _13852_, _06363_);
  or (_13859_, _13858_, _01967_);
  or (_13860_, _13859_, _13857_);
  nor (_13861_, _13749_, _06367_);
  nor (_13862_, _13861_, _06373_);
  nand (_13863_, _13862_, _01967_);
  and (_13864_, _13863_, _13860_);
  or (_13865_, _13864_, _01963_);
  or (_13866_, _13846_, _01964_);
  and (_13867_, _13866_, _02457_);
  and (_13868_, _13867_, _13865_);
  nor (_13869_, _06386_, \oc8051_golden_model_1.SP [6]);
  nor (_13870_, _13869_, _06387_);
  and (_13871_, _13870_, _01953_);
  or (_13872_, _13871_, _13868_);
  and (_13873_, _13872_, _06394_);
  and (_13874_, _13852_, _13322_);
  or (_13875_, _13874_, _04950_);
  or (_13876_, _13875_, _13873_);
  nor (_13877_, _06336_, _04074_);
  or (_13878_, _13838_, _06397_);
  or (_13879_, _13878_, _13877_);
  and (_13880_, _13879_, _13876_);
  or (_13881_, _13880_, _04951_);
  and (_13882_, _04396_, _03748_);
  or (_13883_, _13838_, _05513_);
  or (_13884_, _13883_, _13882_);
  and (_13885_, _13884_, _01923_);
  and (_13886_, _13885_, _13881_);
  nor (_13887_, _09096_, _06336_);
  or (_13888_, _13887_, _13838_);
  and (_13889_, _13888_, _01602_);
  or (_13890_, _13889_, _02019_);
  or (_13891_, _13890_, _13886_);
  and (_13892_, _04396_, _09103_);
  or (_13893_, _13892_, _13838_);
  or (_13894_, _13893_, _04979_);
  and (_13895_, _13894_, _13891_);
  or (_13896_, _13895_, _01650_);
  or (_13897_, _13852_, _01651_);
  and (_13898_, _13897_, _13896_);
  or (_13899_, _13898_, _02018_);
  and (_13900_, _09112_, _04111_);
  or (_13901_, _13838_, _05049_);
  or (_13902_, _13901_, _13900_);
  and (_13903_, _13902_, _02136_);
  and (_13904_, _13903_, _13899_);
  or (_13905_, _13904_, _13841_);
  and (_13906_, _13905_, _05076_);
  or (_13907_, _13838_, _05735_);
  and (_13908_, _13893_, _02039_);
  and (_13909_, _13908_, _13907_);
  or (_13910_, _13909_, _13906_);
  and (_13911_, _13910_, _05082_);
  and (_13912_, _13846_, _02130_);
  and (_13913_, _13912_, _13907_);
  and (_13914_, _13852_, _01666_);
  or (_13915_, _13914_, _02016_);
  or (_13916_, _13915_, _13913_);
  or (_13917_, _13916_, _13911_);
  nor (_13918_, _09111_, _06442_);
  or (_13919_, _13918_, _13838_);
  or (_13920_, _13919_, _05104_);
  and (_13921_, _13920_, _13917_);
  or (_13922_, _13921_, _02126_);
  nor (_13923_, _08974_, _06336_);
  or (_13924_, _13838_, _05474_);
  or (_13925_, _13924_, _13923_);
  and (_13926_, _13925_, _02718_);
  and (_13927_, _13926_, _13922_);
  nor (_13928_, _06371_, _06367_);
  or (_13929_, _13928_, _06372_);
  and (_13930_, _13929_, _02146_);
  or (_13931_, _13930_, _01660_);
  or (_13932_, _13931_, _13927_);
  or (_13933_, _13852_, _05157_);
  and (_13934_, _13933_, _13932_);
  or (_13935_, _13934_, _01585_);
  or (_13936_, _13929_, _01596_);
  and (_13937_, _13936_, _13935_);
  or (_13938_, _13937_, _02164_);
  or (_13939_, _13843_, _02168_);
  and (_13940_, _13939_, _06466_);
  and (_13941_, _13940_, _13938_);
  and (_13942_, _13852_, _06467_);
  or (_13943_, _13942_, _01594_);
  or (_13944_, _13943_, _13941_);
  and (_13945_, _08965_, _04111_);
  or (_13946_, _13838_, _01595_);
  or (_13947_, _13946_, _13945_);
  and (_13948_, _13947_, _26505_);
  and (_13949_, _13948_, _13944_);
  or (_13950_, _13949_, _13837_);
  and (_27858_, _13950_, _25964_);
  not (_13951_, \oc8051_golden_model_1.TCON [0]);
  nor (_13952_, _04119_, _13951_);
  nor (_13953_, _04405_, _06206_);
  nor (_13954_, _13953_, _13952_);
  nor (_13955_, _13954_, _01595_);
  and (_13956_, _04119_, _05531_);
  nor (_13957_, _13956_, _13952_);
  nor (_13958_, _13957_, _05076_);
  not (_13959_, _13958_);
  nor (_13960_, _13959_, _13953_);
  and (_13961_, _04119_, _03677_);
  nor (_13962_, _13952_, _05513_);
  not (_13963_, _13962_);
  nor (_13964_, _13963_, _13961_);
  nor (_13965_, _05167_, _13951_);
  and (_13966_, _07725_, _05167_);
  nor (_13967_, _13966_, _13965_);
  nor (_13968_, _13967_, _02223_);
  and (_13969_, _13954_, _01969_);
  and (_13970_, _04119_, \oc8051_golden_model_1.ACC [0]);
  nor (_13971_, _13970_, _13952_);
  nor (_13972_, _13971_, _05488_);
  nor (_13973_, _04571_, _13951_);
  or (_13974_, _13973_, _01969_);
  nor (_13975_, _13974_, _13972_);
  or (_13976_, _13975_, _06233_);
  nor (_13977_, _13976_, _13969_);
  and (_13978_, _04119_, _03334_);
  nor (_13979_, _13978_, _13952_);
  nor (_13980_, _13979_, _05487_);
  or (_13981_, _13980_, _01963_);
  or (_13982_, _13981_, _13977_);
  nor (_13983_, _13982_, _13968_);
  and (_13984_, _13971_, _01963_);
  nor (_13985_, _13984_, _01957_);
  not (_13986_, _13985_);
  nor (_13987_, _13986_, _13983_);
  and (_13988_, _13952_, _01957_);
  or (_13989_, _13988_, _13987_);
  and (_13990_, _13989_, _04885_);
  nor (_13991_, _13954_, _04885_);
  or (_13992_, _13991_, _13990_);
  nor (_13993_, _13992_, _01924_);
  nor (_13994_, _07759_, _06258_);
  or (_13995_, _13965_, _01925_);
  nor (_13996_, _13995_, _13994_);
  or (_13997_, _13996_, _04950_);
  or (_13998_, _13997_, _13993_);
  or (_13999_, _13979_, _06397_);
  and (_14000_, _13999_, _05513_);
  and (_14001_, _14000_, _13998_);
  nor (_14002_, _14001_, _13964_);
  nor (_14003_, _14002_, _01602_);
  nor (_14004_, _07815_, _06206_);
  or (_14005_, _13952_, _01923_);
  nor (_14006_, _14005_, _14004_);
  or (_14007_, _14006_, _02019_);
  nor (_14008_, _14007_, _14003_);
  nand (_14009_, _13957_, _05049_);
  and (_14010_, _14009_, _06278_);
  nor (_14011_, _14010_, _14008_);
  and (_14012_, _07829_, _04119_);
  nor (_14013_, _14012_, _13952_);
  and (_14014_, _14013_, _02018_);
  nor (_14015_, _14014_, _14011_);
  and (_14016_, _14015_, _02136_);
  and (_14017_, _07834_, _04119_);
  nor (_14018_, _14017_, _13952_);
  nor (_14019_, _14018_, _02136_);
  or (_14020_, _14019_, _14016_);
  and (_14021_, _14020_, _05076_);
  nor (_14022_, _14021_, _13960_);
  nor (_14023_, _14022_, _02130_);
  nor (_14024_, _13952_, _04405_);
  or (_14025_, _14024_, _02131_);
  nor (_14026_, _14025_, _13971_);
  or (_14027_, _14026_, _02016_);
  nor (_14028_, _14027_, _14023_);
  nor (_14029_, _07828_, _06206_);
  nor (_14030_, _14029_, _13952_);
  and (_14031_, _14030_, _02016_);
  nor (_14032_, _14031_, _14028_);
  and (_14033_, _14032_, _05474_);
  nor (_14034_, _07696_, _06206_);
  nor (_14035_, _14034_, _13952_);
  nor (_14036_, _14035_, _05474_);
  or (_14037_, _14036_, _14033_);
  and (_14038_, _14037_, _02168_);
  nor (_14039_, _13954_, _02168_);
  nor (_14040_, _14039_, _02025_);
  not (_14041_, _14040_);
  nor (_14042_, _14041_, _14038_);
  nor (_14043_, _13952_, _02377_);
  nor (_14044_, _14043_, _14042_);
  and (_14045_, _14044_, _01595_);
  nor (_14046_, _14045_, _13955_);
  nand (_14047_, _14046_, _26505_);
  or (_14048_, _26505_, \oc8051_golden_model_1.TCON [0]);
  and (_14049_, _14048_, _25964_);
  and (_27861_, _14049_, _14047_);
  or (_14050_, _08029_, _06206_);
  or (_14051_, _04119_, \oc8051_golden_model_1.TCON [1]);
  and (_14052_, _14051_, _02135_);
  and (_14053_, _14052_, _14050_);
  nor (_14054_, _07953_, _06258_);
  and (_14055_, _06258_, \oc8051_golden_model_1.TCON [1]);
  or (_14056_, _14055_, _01925_);
  or (_14057_, _14056_, _14054_);
  and (_14058_, _07909_, _04119_);
  not (_14059_, _14058_);
  and (_14060_, _14059_, _14051_);
  or (_14061_, _14060_, _02438_);
  nand (_14062_, _04119_, _01705_);
  and (_14063_, _14062_, _14051_);
  and (_14064_, _14063_, _04571_);
  and (_14065_, _05488_, \oc8051_golden_model_1.TCON [1]);
  or (_14066_, _14065_, _01969_);
  or (_14067_, _14066_, _14064_);
  and (_14068_, _14067_, _01968_);
  and (_14069_, _14068_, _14061_);
  and (_14070_, _06206_, \oc8051_golden_model_1.TCON [1]);
  nor (_14071_, _06206_, _03393_);
  or (_14072_, _14071_, _14070_);
  and (_14073_, _14072_, _01967_);
  and (_14074_, _07920_, _05167_);
  or (_14075_, _14074_, _14055_);
  and (_14076_, _14075_, _01959_);
  or (_14077_, _14076_, _14073_);
  or (_14078_, _14077_, _01963_);
  or (_14079_, _14078_, _14069_);
  or (_14080_, _14063_, _01964_);
  and (_14081_, _14080_, _14079_);
  or (_14082_, _14081_, _01957_);
  and (_14083_, _07907_, _05167_);
  or (_14084_, _14083_, _14055_);
  or (_14085_, _14084_, _06229_);
  and (_14086_, _14085_, _04885_);
  and (_14087_, _14086_, _14082_);
  and (_14088_, _07936_, _05167_);
  or (_14089_, _14088_, _14055_);
  and (_14090_, _14089_, _01946_);
  or (_14091_, _14090_, _01924_);
  or (_14092_, _14091_, _14087_);
  and (_14093_, _14092_, _14057_);
  or (_14094_, _14093_, _04950_);
  or (_14095_, _14072_, _06397_);
  and (_14096_, _14095_, _14094_);
  or (_14097_, _14096_, _04951_);
  and (_14098_, _04119_, _03613_);
  or (_14099_, _14070_, _05513_);
  or (_14100_, _14099_, _14098_);
  and (_14101_, _14100_, _01923_);
  and (_14102_, _14101_, _14097_);
  nor (_14103_, _08009_, _06206_);
  or (_14104_, _14103_, _14070_);
  and (_14105_, _14104_, _01602_);
  or (_14106_, _14105_, _14102_);
  and (_14107_, _14106_, _02020_);
  or (_14108_, _08023_, _06206_);
  and (_14109_, _14108_, _02018_);
  nand (_14110_, _04119_, _02676_);
  and (_14111_, _14110_, _02019_);
  or (_14112_, _14111_, _14109_);
  and (_14113_, _14112_, _14051_);
  or (_14114_, _14113_, _14107_);
  and (_14115_, _14114_, _02136_);
  or (_14116_, _14115_, _14053_);
  and (_14117_, _14116_, _05076_);
  or (_14118_, _07893_, _06206_);
  and (_14119_, _14051_, _02039_);
  and (_14120_, _14119_, _14118_);
  or (_14121_, _14120_, _14117_);
  and (_14122_, _14121_, _02131_);
  or (_14123_, _14070_, _05741_);
  and (_14124_, _14063_, _02130_);
  and (_14125_, _14124_, _14123_);
  or (_14126_, _14125_, _14122_);
  and (_14127_, _14126_, _02127_);
  or (_14128_, _14110_, _05741_);
  and (_14129_, _14128_, _02016_);
  or (_14130_, _14062_, _05741_);
  and (_14131_, _14130_, _02126_);
  or (_14132_, _14131_, _14129_);
  and (_14133_, _14132_, _14051_);
  or (_14134_, _14133_, _02164_);
  or (_14135_, _14134_, _14127_);
  or (_14136_, _14060_, _02168_);
  and (_14137_, _14136_, _02377_);
  and (_14138_, _14137_, _14135_);
  and (_14139_, _14084_, _02025_);
  or (_14140_, _14139_, _01594_);
  or (_14141_, _14140_, _14138_);
  or (_14142_, _14058_, _14070_);
  or (_14143_, _14142_, _01595_);
  and (_14144_, _14143_, _14141_);
  and (_14145_, _14144_, _26505_);
  and (_14146_, _26506_, \oc8051_golden_model_1.TCON [1]);
  or (_14147_, _14146_, rst);
  or (_27862_, _14147_, _14145_);
  not (_14148_, \oc8051_golden_model_1.TCON [2]);
  nor (_14149_, _04119_, _14148_);
  and (_14150_, _04119_, _05563_);
  nor (_14151_, _14150_, _14149_);
  and (_14152_, _14151_, _02019_);
  nor (_14153_, _06206_, _03272_);
  nor (_14154_, _14153_, _14149_);
  and (_14155_, _14154_, _04950_);
  nor (_14156_, _08095_, _06206_);
  nor (_14157_, _14156_, _14149_);
  and (_14158_, _14157_, _01969_);
  and (_14159_, _04119_, \oc8051_golden_model_1.ACC [2]);
  nor (_14160_, _14159_, _14149_);
  nor (_14161_, _14160_, _05488_);
  nor (_14162_, _04571_, _14148_);
  or (_14163_, _14162_, _01969_);
  nor (_14164_, _14163_, _14161_);
  or (_14165_, _14164_, _06233_);
  nor (_14166_, _14165_, _14158_);
  nor (_14167_, _14154_, _05487_);
  nor (_14168_, _05167_, _14148_);
  and (_14169_, _08111_, _05167_);
  nor (_14170_, _14169_, _14168_);
  nor (_14171_, _14170_, _02223_);
  nor (_14172_, _14171_, _14167_);
  nand (_14173_, _14172_, _01964_);
  or (_14174_, _14173_, _14166_);
  nand (_14175_, _14160_, _01963_);
  and (_14176_, _14175_, _14174_);
  nor (_14177_, _14176_, _01957_);
  and (_14178_, _08109_, _05167_);
  nor (_14179_, _14178_, _14168_);
  and (_14180_, _14179_, _01957_);
  or (_14181_, _14180_, _01946_);
  nor (_14182_, _14181_, _14177_);
  and (_14183_, _08140_, _05167_);
  nor (_14184_, _14183_, _14168_);
  nor (_14185_, _14184_, _04885_);
  or (_14186_, _14185_, _14182_);
  and (_14187_, _14186_, _01925_);
  nor (_14188_, _08158_, _06258_);
  nor (_14189_, _14168_, _14188_);
  nor (_14190_, _14189_, _01925_);
  or (_14191_, _14190_, _04950_);
  nor (_14192_, _14191_, _14187_);
  nor (_14193_, _14192_, _14155_);
  nor (_14194_, _14193_, _04951_);
  and (_14195_, _04119_, _03564_);
  nor (_14196_, _14149_, _05513_);
  not (_14197_, _14196_);
  nor (_14198_, _14197_, _14195_);
  or (_14199_, _14198_, _01602_);
  nor (_14200_, _14199_, _14194_);
  nor (_14201_, _08216_, _06206_);
  nor (_14202_, _14201_, _14149_);
  nor (_14203_, _14202_, _01923_);
  or (_14204_, _14203_, _02019_);
  nor (_14205_, _14204_, _14200_);
  nor (_14206_, _14205_, _14152_);
  or (_14207_, _14206_, _02018_);
  and (_14208_, _08230_, _04119_);
  or (_14209_, _14208_, _14149_);
  or (_14210_, _14209_, _05049_);
  and (_14211_, _14210_, _02136_);
  and (_14212_, _14211_, _14207_);
  and (_14213_, _08237_, _04119_);
  nor (_14214_, _14213_, _14149_);
  nor (_14215_, _14214_, _02136_);
  nor (_14216_, _14215_, _14212_);
  nor (_14217_, _14216_, _02039_);
  nor (_14218_, _14149_, _05739_);
  not (_14219_, _14218_);
  nor (_14220_, _14151_, _05076_);
  and (_14221_, _14220_, _14219_);
  nor (_14222_, _14221_, _14217_);
  nor (_14223_, _14222_, _02130_);
  or (_14224_, _14218_, _02131_);
  nor (_14225_, _14224_, _14160_);
  or (_14226_, _14225_, _02016_);
  nor (_14227_, _14226_, _14223_);
  nor (_14228_, _08229_, _06206_);
  nor (_14229_, _14228_, _14149_);
  and (_14230_, _14229_, _02016_);
  nor (_14231_, _14230_, _14227_);
  and (_14232_, _14231_, _05474_);
  nor (_14233_, _08236_, _06206_);
  nor (_14234_, _14233_, _14149_);
  nor (_14235_, _14234_, _05474_);
  or (_14236_, _14235_, _14232_);
  and (_14237_, _14236_, _02168_);
  nor (_14238_, _14157_, _02168_);
  or (_14239_, _14238_, _02025_);
  or (_14240_, _14239_, _14237_);
  nand (_14241_, _14179_, _02025_);
  and (_14242_, _14241_, _14240_);
  nor (_14243_, _14242_, _01594_);
  and (_14244_, _08285_, _04119_);
  nor (_14245_, _14244_, _14149_);
  and (_14246_, _14245_, _01594_);
  nor (_14247_, _14246_, _14243_);
  or (_14248_, _14247_, _26506_);
  or (_14249_, _26505_, \oc8051_golden_model_1.TCON [2]);
  and (_14250_, _14249_, _25964_);
  and (_27863_, _14250_, _14248_);
  not (_14251_, \oc8051_golden_model_1.TCON [3]);
  nor (_14252_, _04119_, _14251_);
  and (_14253_, _04119_, _05529_);
  nor (_14254_, _14253_, _14252_);
  and (_14255_, _14254_, _02019_);
  nor (_14256_, _06206_, _03473_);
  nor (_14257_, _14256_, _14252_);
  and (_14258_, _14257_, _04950_);
  nor (_14259_, _08308_, _06258_);
  nor (_14260_, _05167_, _14251_);
  or (_14261_, _14260_, _01925_);
  or (_14262_, _14261_, _14259_);
  nor (_14263_, _08337_, _06206_);
  nor (_14264_, _14263_, _14252_);
  and (_14265_, _14264_, _01969_);
  and (_14266_, _04119_, \oc8051_golden_model_1.ACC [3]);
  nor (_14267_, _14266_, _14252_);
  nor (_14268_, _14267_, _05488_);
  nor (_14269_, _04571_, _14251_);
  or (_14270_, _14269_, _01969_);
  nor (_14271_, _14270_, _14268_);
  or (_14272_, _14271_, _06233_);
  nor (_14273_, _14272_, _14265_);
  nor (_14274_, _14257_, _05487_);
  and (_14275_, _08341_, _05167_);
  nor (_14276_, _14275_, _14260_);
  nor (_14277_, _14276_, _02223_);
  nor (_14278_, _14277_, _14274_);
  nand (_14279_, _14278_, _01964_);
  or (_14280_, _14279_, _14273_);
  nand (_14281_, _14267_, _01963_);
  and (_14282_, _14281_, _14280_);
  and (_14283_, _14282_, _06229_);
  and (_14284_, _08324_, _05167_);
  nor (_14285_, _14284_, _14260_);
  nor (_14286_, _14285_, _06229_);
  or (_14287_, _14286_, _14283_);
  and (_14288_, _14287_, _04885_);
  nor (_14289_, _14260_, _08357_);
  or (_14290_, _14276_, _04885_);
  nor (_14291_, _14290_, _14289_);
  or (_14292_, _14291_, _01924_);
  or (_14293_, _14292_, _14288_);
  and (_14294_, _14293_, _14262_);
  nor (_14295_, _14294_, _04950_);
  nor (_14296_, _14295_, _14258_);
  nor (_14297_, _14296_, _04951_);
  and (_14298_, _04119_, _03516_);
  nor (_14299_, _14252_, _05513_);
  not (_14300_, _14299_);
  nor (_14301_, _14300_, _14298_);
  or (_14302_, _14301_, _01602_);
  nor (_14303_, _14302_, _14297_);
  nor (_14304_, _08425_, _06206_);
  nor (_14305_, _14304_, _14252_);
  nor (_14306_, _14305_, _01923_);
  or (_14307_, _14306_, _02019_);
  nor (_14308_, _14307_, _14303_);
  nor (_14309_, _14308_, _14255_);
  or (_14310_, _14309_, _02018_);
  and (_14311_, _08441_, _04119_);
  or (_14312_, _14311_, _14252_);
  or (_14313_, _14312_, _05049_);
  and (_14314_, _14313_, _02136_);
  and (_14315_, _14314_, _14310_);
  and (_14316_, _08304_, _04119_);
  nor (_14317_, _14316_, _14252_);
  nor (_14318_, _14317_, _02136_);
  nor (_14319_, _14318_, _14315_);
  nor (_14320_, _14319_, _02039_);
  nor (_14321_, _14252_, _05737_);
  not (_14322_, _14321_);
  nor (_14323_, _14254_, _05076_);
  and (_14324_, _14323_, _14322_);
  nor (_14325_, _14324_, _14320_);
  nor (_14326_, _14325_, _02130_);
  or (_14327_, _14321_, _02131_);
  nor (_14328_, _14327_, _14267_);
  or (_14329_, _14328_, _02016_);
  nor (_14330_, _14329_, _14326_);
  nor (_14331_, _08440_, _06206_);
  nor (_14332_, _14331_, _14252_);
  and (_14333_, _14332_, _02016_);
  nor (_14334_, _14333_, _14330_);
  and (_14335_, _14334_, _05474_);
  nor (_14336_, _08303_, _06206_);
  nor (_14337_, _14336_, _14252_);
  nor (_14338_, _14337_, _05474_);
  or (_14339_, _14338_, _14335_);
  and (_14340_, _14339_, _02168_);
  nor (_14341_, _14264_, _02168_);
  or (_14342_, _14341_, _02025_);
  or (_14343_, _14342_, _14340_);
  nand (_14344_, _14285_, _02025_);
  and (_14345_, _14344_, _14343_);
  nor (_14346_, _14345_, _01594_);
  and (_14347_, _08507_, _04119_);
  nor (_14348_, _14347_, _14252_);
  and (_14349_, _14348_, _01594_);
  nor (_14350_, _14349_, _14346_);
  or (_14351_, _14350_, _26506_);
  or (_14352_, _26505_, \oc8051_golden_model_1.TCON [3]);
  and (_14353_, _14352_, _25964_);
  and (_27864_, _14353_, _14351_);
  not (_14354_, \oc8051_golden_model_1.TCON [4]);
  nor (_14355_, _04119_, _14354_);
  and (_14356_, _04119_, _05524_);
  nor (_14357_, _14356_, _14355_);
  and (_14358_, _14357_, _02019_);
  nor (_14359_, _06206_, _04024_);
  nor (_14360_, _14359_, _14355_);
  and (_14361_, _14360_, _04950_);
  nor (_14362_, _05167_, _14354_);
  nor (_14363_, _14362_, _08581_);
  and (_14364_, _08565_, _05167_);
  nor (_14365_, _14364_, _14362_);
  or (_14366_, _14365_, _04885_);
  nor (_14367_, _14366_, _14363_);
  nor (_14368_, _08548_, _06206_);
  nor (_14369_, _14368_, _14355_);
  and (_14370_, _14369_, _01969_);
  and (_14371_, _04119_, \oc8051_golden_model_1.ACC [4]);
  nor (_14372_, _14371_, _14355_);
  nor (_14373_, _14372_, _05488_);
  nor (_14374_, _04571_, _14354_);
  or (_14375_, _14374_, _01969_);
  nor (_14376_, _14375_, _14373_);
  or (_14377_, _14376_, _06233_);
  nor (_14378_, _14377_, _14370_);
  nor (_14379_, _14360_, _05487_);
  nor (_14380_, _14365_, _02223_);
  nor (_14381_, _14380_, _14379_);
  nand (_14382_, _14381_, _01964_);
  or (_14383_, _14382_, _14378_);
  nand (_14384_, _14372_, _01963_);
  and (_14385_, _14384_, _14383_);
  and (_14386_, _14385_, _06229_);
  and (_14387_, _08544_, _05167_);
  nor (_14388_, _14387_, _14362_);
  nor (_14389_, _14388_, _06229_);
  or (_14390_, _14389_, _14386_);
  and (_14391_, _14390_, _04885_);
  nor (_14392_, _14391_, _14367_);
  nor (_14393_, _14392_, _01924_);
  nor (_14394_, _08607_, _06258_);
  nor (_14395_, _14394_, _14362_);
  nor (_14396_, _14395_, _01925_);
  nor (_14397_, _14396_, _04950_);
  not (_14398_, _14397_);
  nor (_14399_, _14398_, _14393_);
  nor (_14400_, _14399_, _14361_);
  nor (_14401_, _14400_, _04951_);
  and (_14402_, _04119_, _03903_);
  nor (_14403_, _14355_, _05513_);
  not (_14404_, _14403_);
  nor (_14405_, _14404_, _14402_);
  or (_14406_, _14405_, _01602_);
  nor (_14407_, _14406_, _14401_);
  nor (_14408_, _08663_, _06206_);
  nor (_14409_, _14408_, _14355_);
  nor (_14410_, _14409_, _01923_);
  or (_14411_, _14410_, _02019_);
  nor (_14412_, _14411_, _14407_);
  nor (_14413_, _14412_, _14358_);
  or (_14414_, _14413_, _02018_);
  and (_14415_, _08531_, _04119_);
  or (_14416_, _14415_, _14355_);
  or (_14417_, _14416_, _05049_);
  and (_14418_, _14417_, _02136_);
  and (_14419_, _14418_, _14414_);
  and (_14420_, _08527_, _04119_);
  nor (_14421_, _14420_, _14355_);
  nor (_14422_, _14421_, _02136_);
  nor (_14423_, _14422_, _14419_);
  nor (_14424_, _14423_, _02039_);
  nor (_14425_, _14355_, _08729_);
  not (_14426_, _14425_);
  nor (_14427_, _14357_, _05076_);
  and (_14428_, _14427_, _14426_);
  nor (_14429_, _14428_, _14424_);
  nor (_14430_, _14429_, _02130_);
  or (_14431_, _14425_, _02131_);
  nor (_14432_, _14431_, _14372_);
  or (_14433_, _14432_, _02016_);
  nor (_14434_, _14433_, _14430_);
  nor (_14435_, _08530_, _06206_);
  nor (_14436_, _14435_, _14355_);
  and (_14437_, _14436_, _02016_);
  nor (_14438_, _14437_, _14434_);
  and (_14439_, _14438_, _05474_);
  nor (_14440_, _08526_, _06206_);
  nor (_14441_, _14440_, _14355_);
  nor (_14442_, _14441_, _05474_);
  or (_14443_, _14442_, _14439_);
  and (_14444_, _14443_, _02168_);
  nor (_14445_, _14369_, _02168_);
  or (_14446_, _14445_, _02025_);
  or (_14447_, _14446_, _14444_);
  nand (_14448_, _14388_, _02025_);
  and (_14449_, _14448_, _14447_);
  nor (_14450_, _14449_, _01594_);
  and (_14451_, _08732_, _04119_);
  nor (_14452_, _14451_, _14355_);
  and (_14453_, _14452_, _01594_);
  nor (_14454_, _14453_, _14450_);
  or (_14455_, _14454_, _26506_);
  or (_14456_, _26505_, \oc8051_golden_model_1.TCON [4]);
  and (_14457_, _14456_, _25964_);
  and (_27865_, _14457_, _14455_);
  not (_14458_, \oc8051_golden_model_1.TCON [5]);
  nor (_14459_, _04119_, _14458_);
  and (_14460_, _04119_, _05548_);
  nor (_14461_, _14460_, _14459_);
  and (_14462_, _14461_, _02019_);
  nor (_14463_, _06206_, _03976_);
  nor (_14464_, _14463_, _14459_);
  and (_14465_, _14464_, _04950_);
  nor (_14466_, _05167_, _14458_);
  nor (_14467_, _14466_, _08801_);
  and (_14468_, _08785_, _05167_);
  nor (_14469_, _14468_, _14466_);
  or (_14470_, _14469_, _04885_);
  nor (_14471_, _14470_, _14467_);
  nor (_14472_, _08771_, _06206_);
  nor (_14473_, _14472_, _14459_);
  and (_14474_, _14473_, _01969_);
  and (_14475_, _04119_, \oc8051_golden_model_1.ACC [5]);
  nor (_14476_, _14475_, _14459_);
  nor (_14477_, _14476_, _05488_);
  nor (_14478_, _04571_, _14458_);
  or (_14479_, _14478_, _01969_);
  nor (_14480_, _14479_, _14477_);
  or (_14481_, _14480_, _06233_);
  nor (_14482_, _14481_, _14474_);
  nor (_14483_, _14464_, _05487_);
  nor (_14484_, _14469_, _02223_);
  nor (_14485_, _14484_, _14483_);
  nand (_14486_, _14485_, _01964_);
  or (_14487_, _14486_, _14482_);
  nand (_14488_, _14476_, _01963_);
  and (_14489_, _14488_, _14487_);
  and (_14490_, _14489_, _06229_);
  and (_14491_, _08768_, _05167_);
  nor (_14492_, _14491_, _14466_);
  nor (_14493_, _14492_, _06229_);
  or (_14494_, _14493_, _14490_);
  and (_14495_, _14494_, _04885_);
  nor (_14496_, _14495_, _14471_);
  nor (_14497_, _14496_, _01924_);
  nor (_14498_, _08754_, _06258_);
  nor (_14499_, _14498_, _14466_);
  nor (_14500_, _14499_, _01925_);
  nor (_14501_, _14500_, _04950_);
  not (_14502_, _14501_);
  nor (_14503_, _14502_, _14497_);
  nor (_14504_, _14503_, _14465_);
  nor (_14505_, _14504_, _04951_);
  and (_14506_, _04119_, _03850_);
  nor (_14507_, _14459_, _05513_);
  not (_14508_, _14507_);
  nor (_14509_, _14508_, _14506_);
  or (_14510_, _14509_, _01602_);
  nor (_14511_, _14510_, _14505_);
  nor (_14512_, _08874_, _06206_);
  nor (_14513_, _14512_, _14459_);
  nor (_14514_, _14513_, _01923_);
  or (_14515_, _14514_, _02019_);
  nor (_14516_, _14515_, _14511_);
  nor (_14517_, _14516_, _14462_);
  or (_14518_, _14517_, _02018_);
  and (_14519_, _08890_, _04119_);
  or (_14520_, _14519_, _14459_);
  or (_14521_, _14520_, _05049_);
  and (_14522_, _14521_, _02136_);
  and (_14523_, _14522_, _14518_);
  and (_14524_, _08750_, _04119_);
  nor (_14525_, _14524_, _14459_);
  nor (_14526_, _14525_, _02136_);
  nor (_14527_, _14526_, _14523_);
  nor (_14528_, _14527_, _02039_);
  nor (_14529_, _14459_, _08946_);
  not (_14530_, _14529_);
  nor (_14531_, _14461_, _05076_);
  and (_14532_, _14531_, _14530_);
  nor (_14533_, _14532_, _14528_);
  nor (_14534_, _14533_, _02130_);
  or (_14535_, _14529_, _02131_);
  nor (_14536_, _14535_, _14476_);
  or (_14537_, _14536_, _02016_);
  nor (_14538_, _14537_, _14534_);
  nor (_14539_, _08889_, _06206_);
  nor (_14540_, _14539_, _14459_);
  and (_14541_, _14540_, _02016_);
  nor (_14542_, _14541_, _14538_);
  and (_14543_, _14542_, _05474_);
  nor (_14544_, _08749_, _06206_);
  nor (_14545_, _14544_, _14459_);
  nor (_14546_, _14545_, _05474_);
  or (_14547_, _14546_, _14543_);
  and (_14548_, _14547_, _02168_);
  nor (_14549_, _14473_, _02168_);
  or (_14550_, _14549_, _02025_);
  or (_14551_, _14550_, _14548_);
  nand (_14552_, _14492_, _02025_);
  and (_14553_, _14552_, _14551_);
  nor (_14554_, _14553_, _01594_);
  and (_14555_, _08949_, _04119_);
  nor (_14556_, _14555_, _14459_);
  and (_14557_, _14556_, _01594_);
  nor (_14558_, _14557_, _14554_);
  or (_14559_, _14558_, _26506_);
  or (_14560_, _26505_, \oc8051_golden_model_1.TCON [5]);
  and (_14561_, _14560_, _25964_);
  and (_27866_, _14561_, _14559_);
  not (_14562_, \oc8051_golden_model_1.TCON [6]);
  nor (_14563_, _04119_, _14562_);
  and (_14564_, _04119_, _03748_);
  or (_14565_, _14564_, _14563_);
  and (_14566_, _14565_, _04951_);
  nor (_14567_, _05167_, _14562_);
  not (_14568_, _14567_);
  and (_14569_, _14568_, _09026_);
  and (_14570_, _09011_, _05167_);
  nor (_14571_, _14570_, _14567_);
  or (_14572_, _14571_, _04885_);
  nor (_14573_, _14572_, _14569_);
  nor (_14574_, _08995_, _06206_);
  nor (_14575_, _14574_, _14563_);
  and (_14576_, _14575_, _01969_);
  and (_14577_, _04119_, \oc8051_golden_model_1.ACC [6]);
  nor (_14578_, _14577_, _14563_);
  nor (_14579_, _14578_, _05488_);
  nor (_14580_, _04571_, _14562_);
  or (_14581_, _14580_, _01969_);
  nor (_14582_, _14581_, _14579_);
  or (_14583_, _14582_, _06233_);
  nor (_14584_, _14583_, _14576_);
  nor (_14585_, _06206_, _04074_);
  nor (_14586_, _14585_, _14563_);
  nor (_14587_, _14586_, _05487_);
  nor (_14588_, _14571_, _02223_);
  nor (_14589_, _14588_, _14587_);
  nand (_14590_, _14589_, _01964_);
  or (_14591_, _14590_, _14584_);
  nand (_14592_, _14578_, _01963_);
  and (_14593_, _14592_, _14591_);
  and (_14594_, _14593_, _06229_);
  and (_14595_, _08992_, _05167_);
  nor (_14596_, _14595_, _14567_);
  nor (_14597_, _14596_, _06229_);
  or (_14598_, _14597_, _14594_);
  and (_14599_, _14598_, _04885_);
  nor (_14600_, _14599_, _14573_);
  nor (_14601_, _14600_, _01924_);
  nor (_14602_, _08979_, _06258_);
  nor (_14603_, _14602_, _14567_);
  nor (_14604_, _14603_, _01925_);
  nor (_14605_, _14604_, _04950_);
  not (_14606_, _14605_);
  nor (_14607_, _14606_, _14601_);
  and (_14608_, _14586_, _04950_);
  or (_14609_, _14608_, _04951_);
  nor (_14610_, _14609_, _14607_);
  or (_14611_, _14610_, _14566_);
  and (_14612_, _14611_, _01923_);
  nor (_14613_, _09096_, _06206_);
  nor (_14614_, _14613_, _14563_);
  nor (_14615_, _14614_, _01923_);
  or (_14616_, _14615_, _06278_);
  or (_14617_, _14616_, _14612_);
  and (_14618_, _09112_, _04119_);
  or (_14619_, _14563_, _05049_);
  or (_14620_, _14619_, _14618_);
  and (_14621_, _04119_, _09103_);
  nor (_14622_, _14621_, _14563_);
  and (_14623_, _14622_, _02019_);
  nor (_14624_, _14623_, _02135_);
  and (_14625_, _14624_, _14620_);
  and (_14626_, _14625_, _14617_);
  and (_14627_, _08975_, _04119_);
  nor (_14628_, _14627_, _14563_);
  nor (_14629_, _14628_, _02136_);
  nor (_14630_, _14629_, _14626_);
  nor (_14631_, _14630_, _02039_);
  nor (_14632_, _14563_, _05735_);
  not (_14633_, _14632_);
  nor (_14634_, _14622_, _05076_);
  and (_14635_, _14634_, _14633_);
  nor (_14636_, _14635_, _14631_);
  nor (_14637_, _14636_, _02130_);
  or (_14638_, _14632_, _02131_);
  nor (_14639_, _14638_, _14578_);
  or (_14640_, _14639_, _02016_);
  nor (_14641_, _14640_, _14637_);
  nor (_14642_, _09111_, _06206_);
  nor (_14643_, _14642_, _14563_);
  and (_14644_, _14643_, _02016_);
  nor (_14645_, _14644_, _14641_);
  and (_14646_, _14645_, _05474_);
  nor (_14647_, _08974_, _06206_);
  nor (_14648_, _14647_, _14563_);
  nor (_14649_, _14648_, _05474_);
  or (_14650_, _14649_, _14646_);
  and (_14651_, _14650_, _02168_);
  nor (_14652_, _14575_, _02168_);
  or (_14653_, _14652_, _02025_);
  or (_14654_, _14653_, _14651_);
  nand (_14655_, _14596_, _02025_);
  and (_14656_, _14655_, _14654_);
  nor (_14657_, _14656_, _01594_);
  and (_14658_, _08965_, _04119_);
  nor (_14659_, _14658_, _14563_);
  and (_14660_, _14659_, _01594_);
  nor (_14661_, _14660_, _14657_);
  or (_14662_, _14661_, _26506_);
  or (_14663_, _26505_, \oc8051_golden_model_1.TCON [6]);
  and (_14664_, _14663_, _25964_);
  and (_27868_, _14664_, _14662_);
  not (_14665_, \oc8051_golden_model_1.TH0 [0]);
  nor (_14666_, _04125_, _14665_);
  nor (_14667_, _04405_, _06128_);
  nor (_14668_, _14667_, _14666_);
  and (_14669_, _14668_, _02266_);
  and (_14670_, _04125_, \oc8051_golden_model_1.ACC [0]);
  nor (_14671_, _14670_, _14666_);
  nor (_14672_, _14671_, _01964_);
  nor (_14673_, _14671_, _05488_);
  nor (_14674_, _04571_, _14665_);
  or (_14675_, _14674_, _14673_);
  and (_14676_, _14675_, _02438_);
  nor (_14677_, _14668_, _02438_);
  or (_14678_, _14677_, _14676_);
  and (_14679_, _14678_, _05487_);
  and (_14680_, _04125_, _03334_);
  nor (_14681_, _14680_, _14666_);
  nor (_14682_, _14681_, _05487_);
  nor (_14683_, _14682_, _14679_);
  nor (_14684_, _14683_, _01963_);
  or (_14685_, _14684_, _04950_);
  nor (_14686_, _14685_, _14672_);
  and (_14687_, _14681_, _04950_);
  nor (_14688_, _14687_, _14686_);
  nor (_14689_, _14688_, _04951_);
  and (_14690_, _04125_, _03677_);
  nor (_14691_, _14666_, _05513_);
  not (_14692_, _14691_);
  nor (_14693_, _14692_, _14690_);
  nor (_14694_, _14693_, _14689_);
  nor (_14695_, _14694_, _01602_);
  nor (_14696_, _07815_, _06128_);
  or (_14697_, _14666_, _01923_);
  nor (_14698_, _14697_, _14696_);
  or (_14699_, _14698_, _02019_);
  nor (_14700_, _14699_, _14695_);
  and (_14701_, _04125_, _05531_);
  nor (_14702_, _14701_, _14666_);
  nand (_14703_, _14702_, _05049_);
  and (_14704_, _14703_, _06278_);
  nor (_14705_, _14704_, _14700_);
  and (_14706_, _07829_, _04125_);
  nor (_14707_, _14706_, _14666_);
  and (_14708_, _14707_, _02018_);
  nor (_14709_, _14708_, _14705_);
  and (_14710_, _14709_, _02136_);
  and (_14711_, _07834_, _04125_);
  nor (_14712_, _14711_, _14666_);
  nor (_14713_, _14712_, _02136_);
  or (_14714_, _14713_, _14710_);
  and (_14715_, _14714_, _05076_);
  or (_14716_, _14702_, _05076_);
  nor (_14717_, _14716_, _14667_);
  nor (_14718_, _14717_, _14715_);
  nor (_14719_, _14718_, _02130_);
  and (_14720_, _07833_, _04125_);
  or (_14721_, _14720_, _14666_);
  and (_14722_, _14721_, _02130_);
  or (_14723_, _14722_, _14719_);
  and (_14724_, _14723_, _05104_);
  nor (_14725_, _07828_, _06128_);
  nor (_14726_, _14725_, _14666_);
  nor (_14727_, _14726_, _05104_);
  or (_14728_, _14727_, _14724_);
  and (_14729_, _14728_, _05474_);
  nor (_14730_, _07696_, _06128_);
  nor (_14731_, _14730_, _14666_);
  nor (_14732_, _14731_, _05474_);
  nor (_14733_, _14732_, _02266_);
  not (_14734_, _14733_);
  nor (_14735_, _14734_, _14729_);
  nor (_14736_, _14735_, _14669_);
  or (_14737_, _14736_, _26506_);
  or (_14738_, _26505_, \oc8051_golden_model_1.TH0 [0]);
  and (_14739_, _14738_, _25964_);
  and (_27869_, _14739_, _14737_);
  nor (_14740_, _04125_, \oc8051_golden_model_1.TH0 [1]);
  and (_14741_, _07909_, _04125_);
  nor (_14742_, _14741_, _14740_);
  nor (_14743_, _14742_, _02168_);
  not (_14744_, _14740_);
  nor (_14745_, _07893_, _06128_);
  nor (_14746_, _14745_, _05076_);
  and (_14747_, _14746_, _14744_);
  nor (_14748_, _08029_, _06128_);
  nor (_14749_, _14748_, _02136_);
  and (_14750_, _14749_, _14744_);
  and (_14751_, _04125_, _03613_);
  not (_14752_, \oc8051_golden_model_1.TH0 [1]);
  nor (_14753_, _04125_, _14752_);
  nor (_14754_, _14753_, _05513_);
  not (_14755_, _14754_);
  nor (_14756_, _14755_, _14751_);
  not (_14757_, _14756_);
  nor (_14758_, _06128_, _03393_);
  nor (_14759_, _14758_, _14753_);
  and (_14760_, _14759_, _04950_);
  and (_14761_, _04125_, _01705_);
  nor (_14762_, _14761_, _14740_);
  and (_14763_, _14762_, _01963_);
  nor (_14764_, _14759_, _05487_);
  and (_14765_, _14762_, _04571_);
  nor (_14766_, _04571_, _14752_);
  or (_14767_, _14766_, _14765_);
  and (_14768_, _14767_, _02438_);
  and (_14769_, _14742_, _01969_);
  or (_14770_, _14769_, _14768_);
  and (_14771_, _14770_, _05487_);
  nor (_14772_, _14771_, _14764_);
  nor (_14773_, _14772_, _01963_);
  or (_14774_, _14773_, _04950_);
  nor (_14775_, _14774_, _14763_);
  nor (_14776_, _14775_, _14760_);
  nor (_14777_, _14776_, _04951_);
  nor (_14778_, _14777_, _01602_);
  and (_14779_, _14778_, _14757_);
  and (_14780_, _08009_, _04125_);
  nor (_14781_, _14780_, _01923_);
  and (_14782_, _14781_, _14744_);
  nor (_14783_, _14782_, _14779_);
  nor (_14784_, _14783_, _06278_);
  nor (_14785_, _08023_, _06128_);
  nor (_14786_, _14785_, _05049_);
  and (_14787_, _04125_, _02676_);
  nor (_14788_, _14787_, _04979_);
  or (_14789_, _14788_, _14786_);
  and (_14790_, _14789_, _14744_);
  nor (_14791_, _14790_, _14784_);
  nor (_14792_, _14791_, _02135_);
  nor (_14793_, _14792_, _14750_);
  nor (_14794_, _14793_, _02039_);
  nor (_14795_, _14794_, _14747_);
  nor (_14796_, _14795_, _02130_);
  nor (_14797_, _14753_, _05741_);
  nor (_14798_, _14797_, _02131_);
  and (_14799_, _14798_, _14762_);
  nor (_14800_, _14799_, _14796_);
  nor (_14801_, _14800_, _02128_);
  and (_14802_, _14787_, _04452_);
  nor (_14803_, _14802_, _05104_);
  nand (_14804_, _14761_, _04452_);
  and (_14805_, _14804_, _02126_);
  or (_14806_, _14805_, _14803_);
  and (_14807_, _14806_, _14744_);
  or (_14808_, _14807_, _02164_);
  nor (_14809_, _14808_, _14801_);
  nor (_14810_, _14809_, _14743_);
  nor (_14811_, _14810_, _01594_);
  nor (_14812_, _14753_, _14741_);
  and (_14813_, _14812_, _01594_);
  nor (_14814_, _14813_, _14811_);
  or (_14815_, _14814_, _26506_);
  or (_14816_, _26505_, \oc8051_golden_model_1.TH0 [1]);
  and (_14817_, _14816_, _25964_);
  and (_27870_, _14817_, _14815_);
  not (_14818_, \oc8051_golden_model_1.TH0 [2]);
  nor (_14819_, _04125_, _14818_);
  nor (_14820_, _14819_, _05739_);
  not (_14821_, _14820_);
  and (_14822_, _04125_, _05563_);
  nor (_14823_, _14822_, _14819_);
  nor (_14824_, _14823_, _05076_);
  and (_14825_, _14824_, _14821_);
  and (_14826_, _04125_, _03564_);
  nor (_14827_, _14826_, _14819_);
  or (_14828_, _14827_, _05513_);
  and (_14829_, _04125_, \oc8051_golden_model_1.ACC [2]);
  nor (_14830_, _14829_, _14819_);
  nor (_14831_, _14830_, _01964_);
  nor (_14832_, _14830_, _05488_);
  nor (_14833_, _04571_, _14818_);
  or (_14834_, _14833_, _14832_);
  and (_14835_, _14834_, _02438_);
  nor (_14836_, _08095_, _06128_);
  nor (_14837_, _14836_, _14819_);
  nor (_14838_, _14837_, _02438_);
  or (_14839_, _14838_, _14835_);
  and (_14840_, _14839_, _05487_);
  nor (_14841_, _06128_, _03272_);
  nor (_14842_, _14841_, _14819_);
  nor (_14843_, _14842_, _05487_);
  nor (_14844_, _14843_, _14840_);
  nor (_14845_, _14844_, _01963_);
  or (_14846_, _14845_, _04950_);
  nor (_14847_, _14846_, _14831_);
  and (_14848_, _14842_, _04950_);
  or (_14849_, _14848_, _04951_);
  or (_14850_, _14849_, _14847_);
  and (_14851_, _14850_, _01923_);
  and (_14852_, _14851_, _14828_);
  nor (_14853_, _08216_, _06128_);
  or (_14854_, _14819_, _01923_);
  nor (_14855_, _14854_, _14853_);
  or (_14856_, _14855_, _02019_);
  nor (_14857_, _14856_, _14852_);
  nand (_14858_, _14823_, _05049_);
  and (_14859_, _14858_, _06278_);
  nor (_14860_, _14859_, _14857_);
  and (_14861_, _08230_, _04125_);
  nor (_14862_, _14861_, _14819_);
  and (_14863_, _14862_, _02018_);
  nor (_14864_, _14863_, _14860_);
  and (_14865_, _14864_, _02136_);
  and (_14866_, _08237_, _04125_);
  nor (_14867_, _14866_, _14819_);
  nor (_14868_, _14867_, _02136_);
  or (_14869_, _14868_, _14865_);
  and (_14870_, _14869_, _05076_);
  nor (_14871_, _14870_, _14825_);
  nor (_14872_, _14871_, _02130_);
  or (_14873_, _14820_, _02131_);
  nor (_14874_, _14873_, _14830_);
  or (_14875_, _14874_, _02016_);
  nor (_14876_, _14875_, _14872_);
  nor (_14877_, _08229_, _06128_);
  nor (_14878_, _14877_, _14819_);
  and (_14879_, _14878_, _02016_);
  nor (_14880_, _14879_, _14876_);
  and (_14881_, _14880_, _05474_);
  nor (_14882_, _08236_, _06128_);
  nor (_14883_, _14882_, _14819_);
  nor (_14884_, _14883_, _05474_);
  or (_14885_, _14884_, _14881_);
  and (_14886_, _14885_, _02168_);
  nor (_14887_, _14837_, _02168_);
  or (_14888_, _14887_, _01594_);
  nor (_14889_, _14888_, _14886_);
  and (_14890_, _08285_, _04125_);
  nor (_14891_, _14890_, _14819_);
  and (_14892_, _14891_, _01594_);
  nor (_14893_, _14892_, _14889_);
  or (_14894_, _14893_, _26506_);
  or (_14895_, _26505_, \oc8051_golden_model_1.TH0 [2]);
  and (_14896_, _14895_, _25964_);
  and (_27871_, _14896_, _14894_);
  not (_14897_, \oc8051_golden_model_1.TH0 [3]);
  nor (_14898_, _04125_, _14897_);
  nor (_14899_, _14898_, _05737_);
  not (_14900_, _14899_);
  and (_14901_, _04125_, _05529_);
  nor (_14902_, _14901_, _14898_);
  nor (_14903_, _14902_, _05076_);
  and (_14904_, _14903_, _14900_);
  and (_14905_, _08304_, _04125_);
  nor (_14906_, _14905_, _14898_);
  nor (_14907_, _14906_, _02136_);
  and (_14908_, _04125_, _03516_);
  or (_14909_, _14908_, _14898_);
  and (_14910_, _14909_, _04951_);
  and (_14911_, _04125_, \oc8051_golden_model_1.ACC [3]);
  nor (_14912_, _14911_, _14898_);
  nor (_14913_, _14912_, _01964_);
  nor (_14914_, _14912_, _05488_);
  nor (_14915_, _04571_, _14897_);
  or (_14916_, _14915_, _14914_);
  and (_14917_, _14916_, _02438_);
  nor (_14918_, _08337_, _06128_);
  nor (_14919_, _14918_, _14898_);
  nor (_14920_, _14919_, _02438_);
  or (_14921_, _14920_, _14917_);
  and (_14922_, _14921_, _05487_);
  nor (_14923_, _06128_, _03473_);
  nor (_14924_, _14923_, _14898_);
  nor (_14925_, _14924_, _05487_);
  nor (_14926_, _14925_, _14922_);
  nor (_14927_, _14926_, _01963_);
  or (_14928_, _14927_, _04950_);
  nor (_14929_, _14928_, _14913_);
  and (_14930_, _14924_, _04950_);
  or (_14931_, _14930_, _04951_);
  nor (_14932_, _14931_, _14929_);
  or (_14933_, _14932_, _14910_);
  and (_14934_, _14933_, _01923_);
  nor (_14935_, _08425_, _06128_);
  nor (_14936_, _14935_, _14898_);
  nor (_14937_, _14936_, _01923_);
  or (_14938_, _14937_, _06278_);
  or (_14939_, _14938_, _14934_);
  and (_14940_, _08441_, _04125_);
  or (_14941_, _14898_, _05049_);
  or (_14942_, _14941_, _14940_);
  and (_14943_, _14902_, _02019_);
  nor (_14944_, _14943_, _02135_);
  and (_14945_, _14944_, _14942_);
  and (_14946_, _14945_, _14939_);
  nor (_14947_, _14946_, _14907_);
  nor (_14948_, _14947_, _02039_);
  nor (_14949_, _14948_, _14904_);
  nor (_14950_, _14949_, _02130_);
  or (_14951_, _14899_, _02131_);
  nor (_14952_, _14951_, _14912_);
  or (_14953_, _14952_, _02016_);
  nor (_14954_, _14953_, _14950_);
  nor (_14955_, _08440_, _06128_);
  nor (_14956_, _14955_, _14898_);
  and (_14957_, _14956_, _02016_);
  nor (_14958_, _14957_, _14954_);
  and (_14959_, _14958_, _05474_);
  nor (_14960_, _08303_, _06128_);
  nor (_14961_, _14960_, _14898_);
  nor (_14962_, _14961_, _05474_);
  or (_14963_, _14962_, _14959_);
  and (_14964_, _14963_, _02168_);
  nor (_14965_, _14919_, _02168_);
  or (_14966_, _14965_, _01594_);
  nor (_14967_, _14966_, _14964_);
  and (_14968_, _08507_, _04125_);
  nor (_14969_, _14968_, _14898_);
  and (_14970_, _14969_, _01594_);
  nor (_14971_, _14970_, _14967_);
  or (_14972_, _14971_, _26506_);
  or (_14973_, _26505_, \oc8051_golden_model_1.TH0 [3]);
  and (_14974_, _14973_, _25964_);
  and (_27872_, _14974_, _14972_);
  not (_14975_, \oc8051_golden_model_1.TH0 [4]);
  nor (_14976_, _04125_, _14975_);
  and (_14977_, _08527_, _04125_);
  nor (_14978_, _14977_, _14976_);
  nor (_14979_, _14978_, _02136_);
  and (_14980_, _04125_, _05524_);
  nor (_14981_, _14980_, _14976_);
  and (_14982_, _14981_, _02019_);
  nor (_14983_, _06128_, _04024_);
  nor (_14984_, _14983_, _14976_);
  and (_14985_, _14984_, _04950_);
  and (_14986_, _04125_, \oc8051_golden_model_1.ACC [4]);
  nor (_14987_, _14986_, _14976_);
  nor (_14988_, _14987_, _01964_);
  nor (_14989_, _14987_, _05488_);
  nor (_14990_, _04571_, _14975_);
  or (_14991_, _14990_, _14989_);
  and (_14992_, _14991_, _02438_);
  nor (_14993_, _08548_, _06128_);
  nor (_14994_, _14993_, _14976_);
  nor (_14995_, _14994_, _02438_);
  or (_14996_, _14995_, _14992_);
  and (_14997_, _14996_, _05487_);
  nor (_14998_, _14984_, _05487_);
  nor (_14999_, _14998_, _14997_);
  nor (_15000_, _14999_, _01963_);
  or (_15001_, _15000_, _04950_);
  nor (_15002_, _15001_, _14988_);
  nor (_15003_, _15002_, _14985_);
  nor (_15004_, _15003_, _04951_);
  and (_15005_, _04125_, _03903_);
  nor (_15006_, _14976_, _05513_);
  not (_15007_, _15006_);
  nor (_15008_, _15007_, _15005_);
  or (_15009_, _15008_, _01602_);
  nor (_15010_, _15009_, _15004_);
  nor (_15011_, _08663_, _06128_);
  nor (_15012_, _15011_, _14976_);
  nor (_15013_, _15012_, _01923_);
  or (_15014_, _15013_, _02019_);
  nor (_15015_, _15014_, _15010_);
  nor (_15016_, _15015_, _14982_);
  or (_15017_, _15016_, _02018_);
  and (_15018_, _08531_, _04125_);
  or (_15019_, _15018_, _14976_);
  or (_15020_, _15019_, _05049_);
  and (_15021_, _15020_, _02136_);
  and (_15022_, _15021_, _15017_);
  nor (_15023_, _15022_, _14979_);
  nor (_15024_, _15023_, _02039_);
  nor (_15025_, _14976_, _08729_);
  not (_15026_, _15025_);
  nor (_15027_, _14981_, _05076_);
  and (_15028_, _15027_, _15026_);
  nor (_15029_, _15028_, _15024_);
  nor (_15030_, _15029_, _02130_);
  or (_15031_, _15025_, _02131_);
  nor (_15032_, _15031_, _14987_);
  or (_15033_, _15032_, _02016_);
  nor (_15034_, _15033_, _15030_);
  nor (_15035_, _08530_, _06128_);
  nor (_15036_, _15035_, _14976_);
  and (_15037_, _15036_, _02016_);
  nor (_15038_, _15037_, _15034_);
  and (_15039_, _15038_, _05474_);
  nor (_15040_, _08526_, _06128_);
  nor (_15041_, _15040_, _14976_);
  nor (_15042_, _15041_, _05474_);
  or (_15043_, _15042_, _15039_);
  and (_15044_, _15043_, _02168_);
  nor (_15045_, _14994_, _02168_);
  or (_15046_, _15045_, _01594_);
  nor (_15047_, _15046_, _15044_);
  and (_15048_, _08732_, _04125_);
  nor (_15049_, _15048_, _14976_);
  and (_15050_, _15049_, _01594_);
  nor (_15051_, _15050_, _15047_);
  or (_15052_, _15051_, _26506_);
  or (_15053_, _26505_, \oc8051_golden_model_1.TH0 [4]);
  and (_15054_, _15053_, _25964_);
  and (_27873_, _15054_, _15052_);
  not (_15055_, \oc8051_golden_model_1.TH0 [5]);
  nor (_15056_, _04125_, _15055_);
  and (_15057_, _08750_, _04125_);
  nor (_15058_, _15057_, _15056_);
  nor (_15059_, _15058_, _02136_);
  nor (_15060_, _08874_, _06128_);
  or (_15061_, _15056_, _01923_);
  or (_15062_, _15061_, _15060_);
  nor (_15063_, _08771_, _06128_);
  nor (_15064_, _15063_, _15056_);
  nor (_15065_, _15064_, _02438_);
  nor (_15066_, _04571_, _15055_);
  and (_15067_, _04125_, \oc8051_golden_model_1.ACC [5]);
  nor (_15068_, _15067_, _15056_);
  nor (_15069_, _15068_, _05488_);
  nor (_15070_, _15069_, _15066_);
  nor (_15071_, _15070_, _01969_);
  or (_15072_, _15071_, _15065_);
  and (_15073_, _15072_, _05487_);
  nor (_15074_, _06128_, _03976_);
  nor (_15075_, _15074_, _15056_);
  nor (_15076_, _15075_, _05487_);
  or (_15077_, _15076_, _15073_);
  and (_15078_, _15077_, _01964_);
  nor (_15079_, _15068_, _01964_);
  nor (_15080_, _15079_, _04950_);
  not (_15081_, _15080_);
  nor (_15082_, _15081_, _15078_);
  and (_15083_, _15075_, _04950_);
  or (_15084_, _15083_, _04951_);
  nor (_15085_, _15084_, _15082_);
  and (_15086_, _04125_, _03850_);
  or (_15087_, _15086_, _15056_);
  and (_15088_, _15087_, _04951_);
  or (_15089_, _15088_, _01602_);
  or (_15090_, _15089_, _15085_);
  and (_15091_, _15090_, _15062_);
  and (_15092_, _15091_, _04979_);
  and (_15093_, _04125_, _05548_);
  nor (_15094_, _15093_, _15056_);
  nor (_15095_, _15094_, _04979_);
  or (_15096_, _15095_, _15092_);
  or (_15097_, _15096_, _02018_);
  and (_15098_, _08890_, _04125_);
  or (_15099_, _15098_, _15056_);
  or (_15100_, _15099_, _05049_);
  and (_15101_, _15100_, _02136_);
  and (_15102_, _15101_, _15097_);
  nor (_15103_, _15102_, _15059_);
  nor (_15104_, _15103_, _02039_);
  nor (_15105_, _15056_, _08946_);
  not (_15106_, _15105_);
  nor (_15107_, _15094_, _05076_);
  and (_15108_, _15107_, _15106_);
  nor (_15109_, _15108_, _15104_);
  nor (_15110_, _15109_, _02130_);
  or (_15111_, _15105_, _02131_);
  nor (_15112_, _15111_, _15068_);
  or (_15113_, _15112_, _02016_);
  nor (_15114_, _15113_, _15110_);
  nor (_15115_, _08889_, _06128_);
  nor (_15116_, _15115_, _15056_);
  and (_15117_, _15116_, _02016_);
  nor (_15118_, _15117_, _15114_);
  and (_15119_, _15118_, _05474_);
  nor (_15120_, _08749_, _06128_);
  nor (_15121_, _15120_, _15056_);
  nor (_15122_, _15121_, _05474_);
  or (_15123_, _15122_, _15119_);
  and (_15124_, _15123_, _02168_);
  nor (_15125_, _15064_, _02168_);
  or (_15126_, _15125_, _01594_);
  nor (_15127_, _15126_, _15124_);
  and (_15128_, _08949_, _04125_);
  nor (_15129_, _15128_, _15056_);
  and (_15130_, _15129_, _01594_);
  nor (_15131_, _15130_, _15127_);
  or (_15132_, _15131_, _26506_);
  or (_15133_, _26505_, \oc8051_golden_model_1.TH0 [5]);
  and (_15134_, _15133_, _25964_);
  and (_27874_, _15134_, _15132_);
  not (_15135_, \oc8051_golden_model_1.TH0 [6]);
  nor (_15136_, _04125_, _15135_);
  nor (_15137_, _15136_, _05735_);
  not (_15138_, _15137_);
  and (_15139_, _04125_, _09103_);
  nor (_15140_, _15139_, _15136_);
  nor (_15141_, _15140_, _05076_);
  and (_15142_, _15141_, _15138_);
  and (_15143_, _08975_, _04125_);
  nor (_15144_, _15143_, _15136_);
  nor (_15145_, _15144_, _02136_);
  and (_15146_, _04125_, _03748_);
  or (_15147_, _15146_, _15136_);
  and (_15148_, _15147_, _04951_);
  and (_15149_, _04125_, \oc8051_golden_model_1.ACC [6]);
  nor (_15150_, _15149_, _15136_);
  nor (_15151_, _15150_, _01964_);
  nor (_15152_, _15150_, _05488_);
  nor (_15153_, _04571_, _15135_);
  or (_15154_, _15153_, _15152_);
  and (_15155_, _15154_, _02438_);
  nor (_15156_, _08995_, _06128_);
  nor (_15157_, _15156_, _15136_);
  nor (_15158_, _15157_, _02438_);
  or (_15159_, _15158_, _15155_);
  and (_15160_, _15159_, _05487_);
  nor (_15161_, _06128_, _04074_);
  nor (_15162_, _15161_, _15136_);
  nor (_15163_, _15162_, _05487_);
  nor (_15164_, _15163_, _15160_);
  nor (_15165_, _15164_, _01963_);
  or (_15166_, _15165_, _04950_);
  nor (_15167_, _15166_, _15151_);
  and (_15168_, _15162_, _04950_);
  or (_15169_, _15168_, _04951_);
  nor (_15170_, _15169_, _15167_);
  or (_15171_, _15170_, _15148_);
  and (_15172_, _15171_, _01923_);
  nor (_15173_, _09096_, _06128_);
  nor (_15174_, _15173_, _15136_);
  nor (_15175_, _15174_, _01923_);
  or (_15176_, _15175_, _06278_);
  or (_15177_, _15176_, _15172_);
  and (_15178_, _09112_, _04125_);
  or (_15179_, _15136_, _05049_);
  or (_15180_, _15179_, _15178_);
  and (_15181_, _15140_, _02019_);
  nor (_15182_, _15181_, _02135_);
  and (_15183_, _15182_, _15180_);
  and (_15184_, _15183_, _15177_);
  nor (_15185_, _15184_, _15145_);
  nor (_15186_, _15185_, _02039_);
  nor (_15187_, _15186_, _15142_);
  nor (_15188_, _15187_, _02130_);
  or (_15189_, _15137_, _02131_);
  nor (_15190_, _15189_, _15150_);
  or (_15191_, _15190_, _02016_);
  nor (_15192_, _15191_, _15188_);
  nor (_15193_, _09111_, _06128_);
  nor (_15194_, _15193_, _15136_);
  and (_15195_, _15194_, _02016_);
  nor (_15196_, _15195_, _15192_);
  and (_15197_, _15196_, _05474_);
  nor (_15198_, _08974_, _06128_);
  nor (_15199_, _15198_, _15136_);
  nor (_15200_, _15199_, _05474_);
  or (_15201_, _15200_, _15197_);
  and (_15202_, _15201_, _02168_);
  nor (_15203_, _15157_, _02168_);
  or (_15204_, _15203_, _01594_);
  nor (_15205_, _15204_, _15202_);
  and (_15206_, _08965_, _04125_);
  nor (_15207_, _15206_, _15136_);
  and (_15208_, _15207_, _01594_);
  nor (_15209_, _15208_, _15205_);
  or (_15210_, _15209_, _26506_);
  or (_15211_, _26505_, \oc8051_golden_model_1.TH0 [6]);
  and (_15212_, _15211_, _25964_);
  and (_27875_, _15212_, _15210_);
  not (_15213_, \oc8051_golden_model_1.TH1 [0]);
  nor (_15214_, _04138_, _15213_);
  nor (_15215_, _04405_, _06046_);
  nor (_15216_, _15215_, _15214_);
  and (_15217_, _15216_, _02266_);
  and (_15218_, _04138_, \oc8051_golden_model_1.ACC [0]);
  nor (_15219_, _15218_, _15214_);
  nor (_15220_, _15219_, _01964_);
  nor (_15221_, _15220_, _04950_);
  nor (_15222_, _15216_, _02438_);
  nor (_15223_, _04571_, _15213_);
  nor (_15224_, _15219_, _05488_);
  nor (_15225_, _15224_, _15223_);
  nor (_15226_, _15225_, _01969_);
  or (_15227_, _15226_, _01967_);
  nor (_15228_, _15227_, _15222_);
  or (_15229_, _15228_, _01963_);
  and (_15230_, _15229_, _15221_);
  and (_15231_, _04138_, _03334_);
  or (_15232_, _15214_, _11952_);
  nor (_15233_, _15232_, _15231_);
  nor (_15234_, _15233_, _15230_);
  nor (_15235_, _15234_, _04951_);
  and (_15236_, _04138_, _03677_);
  nor (_15237_, _15214_, _05513_);
  not (_15238_, _15237_);
  nor (_15239_, _15238_, _15236_);
  nor (_15240_, _15239_, _15235_);
  nor (_15241_, _15240_, _01602_);
  nor (_15242_, _07815_, _06046_);
  or (_15243_, _15214_, _01923_);
  nor (_15244_, _15243_, _15242_);
  or (_15245_, _15244_, _02019_);
  nor (_15246_, _15245_, _15241_);
  and (_15247_, _04138_, _05531_);
  nor (_15248_, _15247_, _15214_);
  nand (_15249_, _15248_, _05049_);
  and (_15250_, _15249_, _06278_);
  nor (_15251_, _15250_, _15246_);
  and (_15252_, _07829_, _04138_);
  nor (_15253_, _15252_, _15214_);
  and (_15254_, _15253_, _02018_);
  nor (_15255_, _15254_, _15251_);
  and (_15256_, _15255_, _02136_);
  and (_15257_, _07834_, _04138_);
  nor (_15258_, _15257_, _15214_);
  nor (_15259_, _15258_, _02136_);
  or (_15260_, _15259_, _15256_);
  and (_15261_, _15260_, _05076_);
  or (_15262_, _15248_, _05076_);
  nor (_15263_, _15262_, _15215_);
  nor (_15264_, _15263_, _15261_);
  nor (_15265_, _15264_, _02130_);
  and (_15266_, _07833_, _04138_);
  or (_15267_, _15266_, _15214_);
  and (_15268_, _15267_, _02130_);
  or (_15269_, _15268_, _15265_);
  and (_15270_, _15269_, _05104_);
  nor (_15271_, _07828_, _06046_);
  nor (_15272_, _15271_, _15214_);
  nor (_15273_, _15272_, _05104_);
  or (_15274_, _15273_, _15270_);
  and (_15275_, _15274_, _05474_);
  nor (_15276_, _07696_, _06046_);
  nor (_15277_, _15276_, _15214_);
  nor (_15278_, _15277_, _05474_);
  nor (_15279_, _15278_, _02266_);
  not (_15280_, _15279_);
  nor (_15281_, _15280_, _15275_);
  nor (_15282_, _15281_, _15217_);
  or (_15283_, _15282_, _26506_);
  or (_15284_, _26505_, \oc8051_golden_model_1.TH1 [0]);
  and (_15285_, _15284_, _25964_);
  and (_27878_, _15285_, _15283_);
  nor (_15286_, _04138_, \oc8051_golden_model_1.TH1 [1]);
  and (_15287_, _07909_, _04138_);
  nor (_15288_, _15287_, _15286_);
  nor (_15289_, _15288_, _02168_);
  not (_15290_, _15286_);
  nor (_15291_, _07893_, _06046_);
  nor (_15292_, _15291_, _05076_);
  and (_15293_, _15292_, _15290_);
  nor (_15294_, _08029_, _06046_);
  nor (_15295_, _15294_, _02136_);
  and (_15296_, _15295_, _15290_);
  and (_15297_, _04138_, _03613_);
  not (_15298_, \oc8051_golden_model_1.TH1 [1]);
  nor (_15299_, _04138_, _15298_);
  nor (_15300_, _15299_, _05513_);
  not (_15301_, _15300_);
  nor (_15302_, _15301_, _15297_);
  not (_15303_, _15302_);
  nor (_15304_, _06046_, _03393_);
  nor (_15305_, _15304_, _15299_);
  and (_15306_, _15305_, _04950_);
  and (_15307_, _04138_, _01705_);
  nor (_15308_, _15307_, _15286_);
  and (_15309_, _15308_, _04571_);
  nor (_15310_, _04571_, _15298_);
  or (_15311_, _15310_, _15309_);
  and (_15312_, _15311_, _02438_);
  and (_15313_, _15288_, _01969_);
  or (_15314_, _15313_, _15312_);
  and (_15315_, _15314_, _05487_);
  nor (_15316_, _15305_, _05487_);
  nor (_15317_, _15316_, _15315_);
  nor (_15318_, _15317_, _01963_);
  and (_15319_, _15308_, _01963_);
  nor (_15320_, _15319_, _04950_);
  not (_15321_, _15320_);
  nor (_15322_, _15321_, _15318_);
  nor (_15323_, _15322_, _15306_);
  nor (_15324_, _15323_, _04951_);
  nor (_15325_, _15324_, _01602_);
  and (_15326_, _15325_, _15303_);
  and (_15327_, _08009_, _04138_);
  nor (_15328_, _15327_, _01923_);
  and (_15329_, _15328_, _15290_);
  nor (_15330_, _15329_, _15326_);
  nor (_15331_, _15330_, _06278_);
  nor (_15332_, _08023_, _06046_);
  nor (_15333_, _15332_, _05049_);
  and (_15334_, _04138_, _02676_);
  nor (_15335_, _15334_, _04979_);
  nor (_15336_, _15335_, _15333_);
  nor (_15337_, _15336_, _15286_);
  nor (_15338_, _15337_, _15331_);
  nor (_15339_, _15338_, _02135_);
  nor (_15340_, _15339_, _15296_);
  nor (_15341_, _15340_, _02039_);
  nor (_15342_, _15341_, _15293_);
  nor (_15343_, _15342_, _02130_);
  nor (_15344_, _15299_, _05741_);
  nor (_15345_, _15344_, _02131_);
  and (_15346_, _15345_, _15308_);
  nor (_15347_, _15346_, _15343_);
  nor (_15348_, _15347_, _02128_);
  and (_15349_, _15334_, _04452_);
  nor (_15350_, _15349_, _05104_);
  nand (_15351_, _15307_, _04452_);
  and (_15352_, _15351_, _02126_);
  or (_15353_, _15352_, _15350_);
  and (_15354_, _15353_, _15290_);
  or (_15355_, _15354_, _02164_);
  nor (_15356_, _15355_, _15348_);
  nor (_15357_, _15356_, _15289_);
  nor (_15358_, _15357_, _01594_);
  nor (_15359_, _15299_, _15287_);
  and (_15360_, _15359_, _01594_);
  nor (_15361_, _15360_, _15358_);
  or (_15362_, _15361_, _26506_);
  or (_15363_, _26505_, \oc8051_golden_model_1.TH1 [1]);
  and (_15364_, _15363_, _25964_);
  and (_27879_, _15364_, _15362_);
  not (_15365_, \oc8051_golden_model_1.TH1 [2]);
  nor (_15366_, _04138_, _15365_);
  and (_15367_, _04138_, _03564_);
  nor (_15368_, _15367_, _15366_);
  or (_15369_, _15368_, _05513_);
  and (_15370_, _04138_, \oc8051_golden_model_1.ACC [2]);
  nor (_15371_, _15370_, _15366_);
  nor (_15372_, _15371_, _01964_);
  nor (_15373_, _15371_, _05488_);
  nor (_15374_, _04571_, _15365_);
  or (_15375_, _15374_, _15373_);
  and (_15376_, _15375_, _02438_);
  nor (_15377_, _08095_, _06046_);
  nor (_15378_, _15377_, _15366_);
  nor (_15379_, _15378_, _02438_);
  or (_15380_, _15379_, _15376_);
  and (_15381_, _15380_, _05487_);
  nor (_15382_, _06046_, _03272_);
  nor (_15383_, _15382_, _15366_);
  nor (_15384_, _15383_, _05487_);
  nor (_15385_, _15384_, _15381_);
  nor (_15386_, _15385_, _01963_);
  or (_15387_, _15386_, _04950_);
  nor (_15388_, _15387_, _15372_);
  and (_15389_, _15383_, _04950_);
  or (_15390_, _15389_, _04951_);
  or (_15391_, _15390_, _15388_);
  and (_15392_, _15391_, _01923_);
  and (_15393_, _15392_, _15369_);
  nor (_15394_, _08216_, _06046_);
  or (_15395_, _15366_, _01923_);
  nor (_15396_, _15395_, _15394_);
  or (_15397_, _15396_, _02019_);
  nor (_15398_, _15397_, _15393_);
  and (_15399_, _04138_, _05563_);
  nor (_15400_, _15399_, _15366_);
  nand (_15401_, _15400_, _05049_);
  and (_15402_, _15401_, _06278_);
  nor (_15403_, _15402_, _15398_);
  and (_15404_, _08230_, _04138_);
  nor (_15405_, _15404_, _15366_);
  and (_15406_, _15405_, _02018_);
  nor (_15407_, _15406_, _15403_);
  and (_15408_, _15407_, _02136_);
  and (_15409_, _08237_, _04138_);
  nor (_15410_, _15409_, _15366_);
  nor (_15411_, _15410_, _02136_);
  or (_15412_, _15411_, _15408_);
  and (_15413_, _15412_, _05076_);
  nor (_15414_, _15366_, _05739_);
  not (_15415_, _15414_);
  nor (_15416_, _15400_, _05076_);
  and (_15417_, _15416_, _15415_);
  nor (_15418_, _15417_, _15413_);
  nor (_15419_, _15418_, _02130_);
  or (_15420_, _15414_, _02131_);
  nor (_15421_, _15420_, _15371_);
  or (_15422_, _15421_, _02016_);
  nor (_15423_, _15422_, _15419_);
  nor (_15424_, _08229_, _06046_);
  nor (_15425_, _15424_, _15366_);
  and (_15426_, _15425_, _02016_);
  nor (_15427_, _15426_, _15423_);
  and (_15428_, _15427_, _05474_);
  nor (_15429_, _08236_, _06046_);
  nor (_15430_, _15429_, _15366_);
  nor (_15431_, _15430_, _05474_);
  or (_15432_, _15431_, _15428_);
  and (_15433_, _15432_, _02168_);
  nor (_15434_, _15378_, _02168_);
  or (_15435_, _15434_, _01594_);
  nor (_15436_, _15435_, _15433_);
  and (_15437_, _08285_, _04138_);
  nor (_15438_, _15437_, _15366_);
  and (_15439_, _15438_, _01594_);
  nor (_15440_, _15439_, _15436_);
  or (_15441_, _15440_, _26506_);
  or (_15442_, _26505_, \oc8051_golden_model_1.TH1 [2]);
  and (_15443_, _15442_, _25964_);
  and (_27880_, _15443_, _15441_);
  not (_15444_, \oc8051_golden_model_1.TH1 [3]);
  nor (_15445_, _04138_, _15444_);
  and (_15446_, _04138_, \oc8051_golden_model_1.ACC [3]);
  nor (_15447_, _15446_, _15445_);
  nor (_15448_, _15447_, _05488_);
  nor (_15449_, _04571_, _15444_);
  or (_15450_, _15449_, _15448_);
  and (_15451_, _15450_, _02438_);
  nor (_15452_, _08337_, _06046_);
  nor (_15453_, _15452_, _15445_);
  nor (_15454_, _15453_, _02438_);
  or (_15455_, _15454_, _15451_);
  and (_15456_, _15455_, _05487_);
  nor (_15457_, _06046_, _03473_);
  nor (_15458_, _15457_, _15445_);
  nor (_15459_, _15458_, _05487_);
  nor (_15460_, _15459_, _15456_);
  nor (_15461_, _15460_, _01963_);
  nor (_15462_, _15447_, _01964_);
  nor (_15463_, _15462_, _04950_);
  not (_15464_, _15463_);
  nor (_15465_, _15464_, _15461_);
  and (_15466_, _15458_, _04950_);
  or (_15467_, _15466_, _04951_);
  or (_15468_, _15467_, _15465_);
  and (_15469_, _04138_, _03516_);
  nor (_15470_, _15469_, _15445_);
  or (_15471_, _15470_, _05513_);
  and (_15472_, _15471_, _01923_);
  and (_15473_, _15472_, _15468_);
  nor (_15474_, _08425_, _06046_);
  or (_15475_, _15445_, _01923_);
  nor (_15476_, _15475_, _15474_);
  or (_15477_, _15476_, _02019_);
  nor (_15478_, _15477_, _15473_);
  and (_15479_, _04138_, _05529_);
  nor (_15480_, _15479_, _15445_);
  nand (_15481_, _15480_, _05049_);
  and (_15482_, _15481_, _06278_);
  nor (_15483_, _15482_, _15478_);
  and (_15484_, _08441_, _04138_);
  nor (_15485_, _15484_, _15445_);
  and (_15486_, _15485_, _02018_);
  nor (_15487_, _15486_, _15483_);
  and (_15488_, _15487_, _02136_);
  and (_15489_, _08304_, _04138_);
  nor (_15490_, _15489_, _15445_);
  nor (_15491_, _15490_, _02136_);
  or (_15492_, _15491_, _15488_);
  and (_15493_, _15492_, _05076_);
  nor (_15494_, _15445_, _05737_);
  not (_15495_, _15494_);
  nor (_15496_, _15480_, _05076_);
  and (_15497_, _15496_, _15495_);
  nor (_15498_, _15497_, _15493_);
  nor (_15499_, _15498_, _02130_);
  or (_15500_, _15494_, _02131_);
  nor (_15501_, _15500_, _15447_);
  or (_15502_, _15501_, _02016_);
  nor (_15503_, _15502_, _15499_);
  nor (_15504_, _08440_, _06046_);
  nor (_15505_, _15504_, _15445_);
  and (_15506_, _15505_, _02016_);
  nor (_15507_, _15506_, _15503_);
  and (_15508_, _15507_, _05474_);
  nor (_15510_, _08303_, _06046_);
  nor (_15511_, _15510_, _15445_);
  nor (_15512_, _15511_, _05474_);
  or (_15513_, _15512_, _15508_);
  and (_15514_, _15513_, _02168_);
  nor (_15515_, _15453_, _02168_);
  or (_15516_, _15515_, _01594_);
  nor (_15517_, _15516_, _15514_);
  and (_15518_, _08507_, _04138_);
  nor (_15519_, _15518_, _15445_);
  and (_15521_, _15519_, _01594_);
  nor (_15522_, _15521_, _15517_);
  or (_15523_, _15522_, _26506_);
  or (_15524_, _26505_, \oc8051_golden_model_1.TH1 [3]);
  and (_15525_, _15524_, _25964_);
  and (_27881_, _15525_, _15523_);
  not (_15526_, \oc8051_golden_model_1.TH1 [4]);
  nor (_15527_, _04138_, _15526_);
  and (_15528_, _08527_, _04138_);
  nor (_15529_, _15528_, _15527_);
  nor (_15530_, _15529_, _02136_);
  and (_15531_, _04138_, _05524_);
  nor (_15532_, _15531_, _15527_);
  and (_15533_, _15532_, _02019_);
  nor (_15534_, _06046_, _04024_);
  nor (_15535_, _15534_, _15527_);
  and (_15536_, _15535_, _04950_);
  and (_15537_, _04138_, \oc8051_golden_model_1.ACC [4]);
  nor (_15538_, _15537_, _15527_);
  nor (_15539_, _15538_, _01964_);
  nor (_15542_, _15538_, _05488_);
  nor (_15543_, _04571_, _15526_);
  or (_15544_, _15543_, _15542_);
  and (_15545_, _15544_, _02438_);
  nor (_15546_, _08548_, _06046_);
  nor (_15547_, _15546_, _15527_);
  nor (_15548_, _15547_, _02438_);
  or (_15549_, _15548_, _15545_);
  and (_15550_, _15549_, _05487_);
  nor (_15551_, _15535_, _05487_);
  nor (_15553_, _15551_, _15550_);
  nor (_15554_, _15553_, _01963_);
  or (_15555_, _15554_, _04950_);
  nor (_15556_, _15555_, _15539_);
  nor (_15557_, _15556_, _15536_);
  nor (_15558_, _15557_, _04951_);
  and (_15559_, _04138_, _03903_);
  nor (_15560_, _15527_, _05513_);
  not (_15561_, _15560_);
  nor (_15562_, _15561_, _15559_);
  or (_15564_, _15562_, _01602_);
  nor (_15565_, _15564_, _15558_);
  nor (_15566_, _08663_, _06046_);
  nor (_15567_, _15566_, _15527_);
  nor (_15568_, _15567_, _01923_);
  or (_15569_, _15568_, _02019_);
  nor (_15570_, _15569_, _15565_);
  nor (_15571_, _15570_, _15533_);
  or (_15572_, _15571_, _02018_);
  and (_15573_, _08531_, _04138_);
  or (_15575_, _15573_, _15527_);
  or (_15576_, _15575_, _05049_);
  and (_15577_, _15576_, _02136_);
  and (_15578_, _15577_, _15572_);
  nor (_15579_, _15578_, _15530_);
  nor (_15580_, _15579_, _02039_);
  nor (_15581_, _15527_, _08729_);
  not (_15582_, _15581_);
  nor (_15583_, _15532_, _05076_);
  and (_15584_, _15583_, _15582_);
  nor (_15586_, _15584_, _15580_);
  nor (_15587_, _15586_, _02130_);
  or (_15588_, _15581_, _02131_);
  nor (_15589_, _15588_, _15538_);
  or (_15590_, _15589_, _02016_);
  nor (_15591_, _15590_, _15587_);
  nor (_15592_, _08530_, _06046_);
  nor (_15593_, _15592_, _15527_);
  and (_15594_, _15593_, _02016_);
  nor (_15595_, _15594_, _15591_);
  and (_15597_, _15595_, _05474_);
  nor (_15598_, _08526_, _06046_);
  nor (_15599_, _15598_, _15527_);
  nor (_15600_, _15599_, _05474_);
  or (_15601_, _15600_, _15597_);
  and (_15602_, _15601_, _02168_);
  nor (_15603_, _15547_, _02168_);
  or (_15604_, _15603_, _01594_);
  nor (_15605_, _15604_, _15602_);
  and (_15606_, _08732_, _04138_);
  nor (_15608_, _15606_, _15527_);
  and (_15609_, _15608_, _01594_);
  nor (_15610_, _15609_, _15605_);
  or (_15611_, _15610_, _26506_);
  or (_15612_, _26505_, \oc8051_golden_model_1.TH1 [4]);
  and (_15613_, _15612_, _25964_);
  and (_27882_, _15613_, _15611_);
  not (_15614_, \oc8051_golden_model_1.TH1 [5]);
  nor (_15615_, _04138_, _15614_);
  and (_15616_, _08750_, _04138_);
  nor (_15618_, _15616_, _15615_);
  nor (_15619_, _15618_, _02136_);
  and (_15620_, _04138_, _05548_);
  nor (_15621_, _15620_, _15615_);
  and (_15622_, _15621_, _02019_);
  and (_15623_, _04138_, \oc8051_golden_model_1.ACC [5]);
  nor (_15624_, _15623_, _15615_);
  nor (_15625_, _15624_, _01964_);
  nor (_15626_, _15624_, _05488_);
  nor (_15627_, _04571_, _15614_);
  or (_15629_, _15627_, _15626_);
  and (_15630_, _15629_, _02438_);
  nor (_15631_, _08771_, _06046_);
  nor (_15632_, _15631_, _15615_);
  nor (_15633_, _15632_, _02438_);
  or (_15634_, _15633_, _15630_);
  and (_15635_, _15634_, _05487_);
  nor (_15636_, _06046_, _03976_);
  nor (_15637_, _15636_, _15615_);
  nor (_15638_, _15637_, _05487_);
  nor (_15640_, _15638_, _15635_);
  nor (_15641_, _15640_, _01963_);
  or (_15642_, _15641_, _04950_);
  nor (_15643_, _15642_, _15625_);
  and (_15644_, _15637_, _04950_);
  nor (_15645_, _15644_, _15643_);
  nor (_15646_, _15645_, _04951_);
  and (_15647_, _04138_, _03850_);
  nor (_15648_, _15615_, _05513_);
  not (_15649_, _15648_);
  nor (_15651_, _15649_, _15647_);
  or (_15652_, _15651_, _01602_);
  nor (_15653_, _15652_, _15646_);
  nor (_15654_, _08874_, _06046_);
  nor (_15655_, _15654_, _15615_);
  nor (_15656_, _15655_, _01923_);
  or (_15657_, _15656_, _02019_);
  nor (_15658_, _15657_, _15653_);
  nor (_15659_, _15658_, _15622_);
  or (_15660_, _15659_, _02018_);
  and (_15662_, _08890_, _04138_);
  or (_15663_, _15662_, _15615_);
  or (_15664_, _15663_, _05049_);
  and (_15665_, _15664_, _02136_);
  and (_15666_, _15665_, _15660_);
  nor (_15667_, _15666_, _15619_);
  nor (_15668_, _15667_, _02039_);
  nor (_15669_, _15615_, _08946_);
  not (_15670_, _15669_);
  nor (_15671_, _15621_, _05076_);
  and (_15673_, _15671_, _15670_);
  nor (_15674_, _15673_, _15668_);
  nor (_15675_, _15674_, _02130_);
  or (_15676_, _15669_, _02131_);
  nor (_15677_, _15676_, _15624_);
  or (_15678_, _15677_, _02016_);
  nor (_15679_, _15678_, _15675_);
  nor (_15680_, _08889_, _06046_);
  nor (_15681_, _15680_, _15615_);
  and (_15682_, _15681_, _02016_);
  nor (_15684_, _15682_, _15679_);
  and (_15685_, _15684_, _05474_);
  nor (_15686_, _08749_, _06046_);
  nor (_15687_, _15686_, _15615_);
  nor (_15688_, _15687_, _05474_);
  or (_15689_, _15688_, _15685_);
  and (_15690_, _15689_, _02168_);
  nor (_15691_, _15632_, _02168_);
  or (_15692_, _15691_, _01594_);
  nor (_15693_, _15692_, _15690_);
  and (_15695_, _08949_, _04138_);
  nor (_15696_, _15695_, _15615_);
  and (_15697_, _15696_, _01594_);
  nor (_15698_, _15697_, _15693_);
  or (_15699_, _15698_, _26506_);
  or (_15700_, _26505_, \oc8051_golden_model_1.TH1 [5]);
  and (_15701_, _15700_, _25964_);
  and (_27883_, _15701_, _15699_);
  not (_15702_, \oc8051_golden_model_1.TH1 [6]);
  nor (_15703_, _04138_, _15702_);
  and (_15705_, _08975_, _04138_);
  nor (_15706_, _15705_, _15703_);
  nor (_15707_, _15706_, _02136_);
  and (_15708_, _04138_, _03748_);
  or (_15709_, _15708_, _15703_);
  and (_15710_, _15709_, _04951_);
  and (_15711_, _04138_, \oc8051_golden_model_1.ACC [6]);
  nor (_15712_, _15711_, _15703_);
  nor (_15713_, _15712_, _01964_);
  nor (_15714_, _15712_, _05488_);
  nor (_15716_, _04571_, _15702_);
  or (_15717_, _15716_, _15714_);
  and (_15718_, _15717_, _02438_);
  nor (_15719_, _08995_, _06046_);
  nor (_15720_, _15719_, _15703_);
  nor (_15721_, _15720_, _02438_);
  or (_15722_, _15721_, _15718_);
  and (_15723_, _15722_, _05487_);
  nor (_15724_, _06046_, _04074_);
  nor (_15725_, _15724_, _15703_);
  nor (_15727_, _15725_, _05487_);
  nor (_15728_, _15727_, _15723_);
  nor (_15729_, _15728_, _01963_);
  or (_15730_, _15729_, _04950_);
  nor (_15731_, _15730_, _15713_);
  and (_15732_, _15725_, _04950_);
  or (_15733_, _15732_, _04951_);
  nor (_15734_, _15733_, _15731_);
  or (_15735_, _15734_, _15710_);
  and (_15736_, _15735_, _01923_);
  nor (_15738_, _09096_, _06046_);
  nor (_15739_, _15738_, _15703_);
  nor (_15740_, _15739_, _01923_);
  or (_15741_, _15740_, _06278_);
  or (_15742_, _15741_, _15736_);
  and (_15743_, _09112_, _04138_);
  or (_15744_, _15703_, _05049_);
  or (_15745_, _15744_, _15743_);
  and (_15746_, _04138_, _09103_);
  nor (_15747_, _15746_, _15703_);
  and (_15749_, _15747_, _02019_);
  nor (_15750_, _15749_, _02135_);
  and (_15751_, _15750_, _15745_);
  and (_15752_, _15751_, _15742_);
  nor (_15753_, _15752_, _15707_);
  nor (_15754_, _15753_, _02039_);
  nor (_15755_, _15703_, _05735_);
  not (_15756_, _15755_);
  nor (_15757_, _15747_, _05076_);
  and (_15758_, _15757_, _15756_);
  nor (_15760_, _15758_, _15754_);
  nor (_15761_, _15760_, _02130_);
  or (_15762_, _15755_, _02131_);
  nor (_15763_, _15762_, _15712_);
  or (_15764_, _15763_, _02016_);
  nor (_15765_, _15764_, _15761_);
  nor (_15766_, _09111_, _06046_);
  nor (_15767_, _15766_, _15703_);
  and (_15768_, _15767_, _02016_);
  nor (_15769_, _15768_, _15765_);
  and (_15771_, _15769_, _05474_);
  nor (_15772_, _08974_, _06046_);
  nor (_15773_, _15772_, _15703_);
  nor (_15774_, _15773_, _05474_);
  or (_15775_, _15774_, _15771_);
  and (_15776_, _15775_, _02168_);
  nor (_15777_, _15720_, _02168_);
  or (_15778_, _15777_, _01594_);
  nor (_15779_, _15778_, _15776_);
  and (_15780_, _08965_, _04138_);
  nor (_15782_, _15780_, _15703_);
  and (_15783_, _15782_, _01594_);
  nor (_15784_, _15783_, _15779_);
  or (_15785_, _15784_, _26506_);
  or (_15786_, _26505_, \oc8051_golden_model_1.TH1 [6]);
  and (_15787_, _15786_, _25964_);
  and (_27884_, _15787_, _15785_);
  not (_15788_, \oc8051_golden_model_1.TL0 [0]);
  nor (_15789_, _04143_, _15788_);
  nor (_15790_, _04405_, _05963_);
  nor (_15792_, _15790_, _15789_);
  and (_15793_, _15792_, _02266_);
  and (_15794_, _04143_, _03334_);
  nor (_15795_, _15794_, _15789_);
  and (_15796_, _15795_, _04950_);
  and (_15797_, _04143_, \oc8051_golden_model_1.ACC [0]);
  nor (_15798_, _15797_, _15789_);
  nor (_15799_, _15798_, _05488_);
  nor (_15800_, _04571_, _15788_);
  or (_15801_, _15800_, _15799_);
  and (_15803_, _15801_, _02438_);
  nor (_15804_, _15792_, _02438_);
  or (_15805_, _15804_, _15803_);
  and (_15806_, _15805_, _05487_);
  nor (_15807_, _15795_, _05487_);
  nor (_15808_, _15807_, _15806_);
  nor (_15809_, _15808_, _01963_);
  nor (_15810_, _15798_, _01964_);
  nor (_15811_, _15810_, _04950_);
  not (_15812_, _15811_);
  nor (_15814_, _15812_, _15809_);
  nor (_15815_, _15814_, _15796_);
  nor (_15816_, _15815_, _04951_);
  and (_15817_, _04143_, _03677_);
  nor (_15818_, _15789_, _05513_);
  not (_15819_, _15818_);
  nor (_15820_, _15819_, _15817_);
  nor (_15821_, _15820_, _15816_);
  nor (_15822_, _15821_, _01602_);
  nor (_15823_, _07815_, _05963_);
  or (_15825_, _15789_, _01923_);
  nor (_15826_, _15825_, _15823_);
  or (_15827_, _15826_, _02019_);
  nor (_15828_, _15827_, _15822_);
  and (_15829_, _04143_, _05531_);
  nor (_15830_, _15829_, _15789_);
  nand (_15831_, _15830_, _05049_);
  and (_15832_, _15831_, _06278_);
  nor (_15833_, _15832_, _15828_);
  and (_15834_, _07829_, _04143_);
  nor (_15836_, _15834_, _15789_);
  and (_15837_, _15836_, _02018_);
  nor (_15838_, _15837_, _15833_);
  and (_15839_, _15838_, _02136_);
  and (_15840_, _07834_, _04143_);
  nor (_15841_, _15840_, _15789_);
  nor (_15842_, _15841_, _02136_);
  or (_15843_, _15842_, _15839_);
  and (_15844_, _15843_, _05076_);
  or (_15845_, _15830_, _05076_);
  nor (_15847_, _15845_, _15790_);
  nor (_15848_, _15847_, _15844_);
  nor (_15849_, _15848_, _02130_);
  and (_15850_, _07833_, _04143_);
  or (_15851_, _15850_, _15789_);
  and (_15852_, _15851_, _02130_);
  or (_15853_, _15852_, _15849_);
  and (_15854_, _15853_, _05104_);
  nor (_15855_, _07828_, _05963_);
  nor (_15856_, _15855_, _15789_);
  nor (_15858_, _15856_, _05104_);
  or (_15859_, _15858_, _15854_);
  and (_15860_, _15859_, _05474_);
  nor (_15861_, _07696_, _05963_);
  nor (_15862_, _15861_, _15789_);
  nor (_15863_, _15862_, _05474_);
  nor (_15864_, _15863_, _02266_);
  not (_15865_, _15864_);
  nor (_15866_, _15865_, _15860_);
  nor (_15867_, _15866_, _15793_);
  or (_15869_, _15867_, _26506_);
  or (_15870_, _26505_, \oc8051_golden_model_1.TL0 [0]);
  and (_15871_, _15870_, _25964_);
  and (_27887_, _15871_, _15869_);
  nor (_15872_, _04143_, \oc8051_golden_model_1.TL0 [1]);
  and (_15873_, _07909_, _04143_);
  nor (_15874_, _15873_, _15872_);
  nor (_15875_, _15874_, _02168_);
  not (_15876_, _15872_);
  nor (_15877_, _08029_, _05963_);
  nor (_15879_, _15877_, _02136_);
  and (_15880_, _15879_, _15876_);
  and (_15881_, _04143_, _03613_);
  not (_15882_, \oc8051_golden_model_1.TL0 [1]);
  nor (_15883_, _04143_, _15882_);
  nor (_15884_, _15883_, _05513_);
  not (_15885_, _15884_);
  nor (_15886_, _15885_, _15881_);
  not (_15887_, _15886_);
  nor (_15888_, _05963_, _03393_);
  nor (_15890_, _15888_, _15883_);
  and (_15891_, _15890_, _04950_);
  and (_15892_, _04143_, _01705_);
  nor (_15893_, _15892_, _15872_);
  and (_15894_, _15893_, _04571_);
  nor (_15895_, _04571_, _15882_);
  or (_15896_, _15895_, _15894_);
  and (_15897_, _15896_, _02438_);
  and (_15898_, _15874_, _01969_);
  or (_15899_, _15898_, _15897_);
  and (_15901_, _15899_, _05487_);
  nor (_15902_, _15890_, _05487_);
  nor (_15903_, _15902_, _15901_);
  nor (_15904_, _15903_, _01963_);
  and (_15905_, _15893_, _01963_);
  nor (_15906_, _15905_, _04950_);
  not (_15907_, _15906_);
  nor (_15908_, _15907_, _15904_);
  nor (_15909_, _15908_, _15891_);
  nor (_15910_, _15909_, _04951_);
  nor (_15912_, _15910_, _01602_);
  and (_15913_, _15912_, _15887_);
  and (_15914_, _08009_, _04143_);
  nor (_15915_, _15914_, _01923_);
  and (_15916_, _15915_, _15876_);
  nor (_15917_, _15916_, _15913_);
  nor (_15918_, _15917_, _06278_);
  nor (_15919_, _08023_, _05963_);
  nor (_15920_, _15919_, _05049_);
  and (_15921_, _04143_, _02676_);
  nor (_15923_, _15921_, _04979_);
  or (_15924_, _15923_, _15920_);
  and (_15925_, _15924_, _15876_);
  nor (_15926_, _15925_, _15918_);
  nor (_15927_, _15926_, _02135_);
  nor (_15928_, _15927_, _15880_);
  nor (_15929_, _15928_, _02039_);
  nor (_15930_, _07893_, _05963_);
  nor (_15931_, _15930_, _05076_);
  and (_15932_, _15931_, _15876_);
  nor (_15934_, _15932_, _15929_);
  nor (_15935_, _15934_, _02130_);
  nor (_15936_, _15883_, _05741_);
  nor (_15937_, _15936_, _02131_);
  and (_15938_, _15937_, _15893_);
  nor (_15939_, _15938_, _15935_);
  nor (_15940_, _15939_, _02128_);
  and (_15941_, _15921_, _04452_);
  nor (_15942_, _15941_, _05104_);
  and (_15943_, _15892_, _04452_);
  nor (_15945_, _15943_, _05474_);
  or (_15946_, _15945_, _15942_);
  and (_15947_, _15946_, _15876_);
  or (_15948_, _15947_, _02164_);
  nor (_15949_, _15948_, _15940_);
  nor (_15950_, _15949_, _15875_);
  nor (_15951_, _15950_, _01594_);
  nor (_15952_, _15883_, _15873_);
  and (_15953_, _15952_, _01594_);
  nor (_15954_, _15953_, _15951_);
  or (_15956_, _15954_, _26506_);
  or (_15957_, _26505_, \oc8051_golden_model_1.TL0 [1]);
  and (_15958_, _15957_, _25964_);
  and (_27888_, _15958_, _15956_);
  not (_15959_, \oc8051_golden_model_1.TL0 [2]);
  nor (_15960_, _04143_, _15959_);
  and (_15961_, _04143_, _03564_);
  nor (_15962_, _15961_, _15960_);
  or (_15963_, _15962_, _05513_);
  and (_15964_, _04143_, \oc8051_golden_model_1.ACC [2]);
  nor (_15966_, _15964_, _15960_);
  nor (_15967_, _15966_, _01964_);
  nor (_15968_, _15966_, _05488_);
  nor (_15969_, _04571_, _15959_);
  or (_15970_, _15969_, _15968_);
  and (_15971_, _15970_, _02438_);
  nor (_15972_, _08095_, _05963_);
  nor (_15973_, _15972_, _15960_);
  nor (_15974_, _15973_, _02438_);
  or (_15975_, _15974_, _15971_);
  and (_15977_, _15975_, _05487_);
  nor (_15978_, _05963_, _03272_);
  nor (_15979_, _15978_, _15960_);
  nor (_15980_, _15979_, _05487_);
  nor (_15981_, _15980_, _15977_);
  nor (_15982_, _15981_, _01963_);
  or (_15983_, _15982_, _04950_);
  nor (_15984_, _15983_, _15967_);
  and (_15985_, _15979_, _04950_);
  or (_15986_, _15985_, _04951_);
  or (_15988_, _15986_, _15984_);
  and (_15989_, _15988_, _01923_);
  and (_15990_, _15989_, _15963_);
  nor (_15991_, _08216_, _05963_);
  or (_15992_, _15960_, _01923_);
  nor (_15993_, _15992_, _15991_);
  or (_15994_, _15993_, _02019_);
  nor (_15995_, _15994_, _15990_);
  and (_15996_, _04143_, _05563_);
  nor (_15997_, _15996_, _15960_);
  nand (_15999_, _15997_, _05049_);
  and (_16000_, _15999_, _06278_);
  nor (_16001_, _16000_, _15995_);
  and (_16002_, _08230_, _04143_);
  nor (_16003_, _16002_, _15960_);
  and (_16004_, _16003_, _02018_);
  nor (_16005_, _16004_, _16001_);
  and (_16006_, _16005_, _02136_);
  and (_16007_, _08237_, _04143_);
  nor (_16008_, _16007_, _15960_);
  nor (_16010_, _16008_, _02136_);
  or (_16011_, _16010_, _16006_);
  and (_16012_, _16011_, _05076_);
  nor (_16013_, _15960_, _05739_);
  not (_16014_, _16013_);
  nor (_16015_, _15997_, _05076_);
  and (_16016_, _16015_, _16014_);
  nor (_16017_, _16016_, _16012_);
  nor (_16018_, _16017_, _02130_);
  or (_16019_, _16013_, _02131_);
  nor (_16021_, _16019_, _15966_);
  or (_16022_, _16021_, _02016_);
  nor (_16023_, _16022_, _16018_);
  nor (_16024_, _08229_, _05963_);
  nor (_16025_, _16024_, _15960_);
  and (_16026_, _16025_, _02016_);
  nor (_16027_, _16026_, _16023_);
  and (_16028_, _16027_, _05474_);
  nor (_16029_, _08236_, _05963_);
  nor (_16030_, _16029_, _15960_);
  nor (_16032_, _16030_, _05474_);
  or (_16033_, _16032_, _16028_);
  and (_16034_, _16033_, _02168_);
  nand (_16035_, _15973_, _01595_);
  and (_16036_, _16035_, _02266_);
  nor (_16037_, _16036_, _16034_);
  and (_16038_, _08285_, _04143_);
  nor (_16039_, _16038_, _15960_);
  and (_16040_, _16039_, _01594_);
  nor (_16041_, _16040_, _16037_);
  or (_16043_, _16041_, _26506_);
  or (_16044_, _26505_, \oc8051_golden_model_1.TL0 [2]);
  and (_16045_, _16044_, _25964_);
  and (_27889_, _16045_, _16043_);
  not (_16046_, \oc8051_golden_model_1.TL0 [3]);
  nor (_16047_, _04143_, _16046_);
  and (_16048_, _04143_, \oc8051_golden_model_1.ACC [3]);
  nor (_16049_, _16048_, _16047_);
  nor (_16050_, _16049_, _05488_);
  nor (_16051_, _04571_, _16046_);
  or (_16053_, _16051_, _16050_);
  and (_16054_, _16053_, _02438_);
  nor (_16055_, _08337_, _05963_);
  nor (_16056_, _16055_, _16047_);
  nor (_16057_, _16056_, _02438_);
  or (_16058_, _16057_, _16054_);
  and (_16059_, _16058_, _05487_);
  nor (_16060_, _05963_, _03473_);
  nor (_16061_, _16060_, _16047_);
  nor (_16062_, _16061_, _05487_);
  nor (_16064_, _16062_, _16059_);
  nor (_16065_, _16064_, _01963_);
  nor (_16066_, _16049_, _01964_);
  nor (_16067_, _16066_, _04950_);
  not (_16068_, _16067_);
  nor (_16069_, _16068_, _16065_);
  and (_16070_, _16061_, _04950_);
  or (_16071_, _16070_, _04951_);
  or (_16072_, _16071_, _16069_);
  and (_16073_, _04143_, _03516_);
  nor (_16075_, _16073_, _16047_);
  or (_16076_, _16075_, _05513_);
  and (_16077_, _16076_, _01923_);
  and (_16078_, _16077_, _16072_);
  nor (_16079_, _08425_, _05963_);
  or (_16080_, _16047_, _01923_);
  nor (_16081_, _16080_, _16079_);
  or (_16082_, _16081_, _02019_);
  nor (_16083_, _16082_, _16078_);
  and (_16084_, _04143_, _05529_);
  nor (_16086_, _16084_, _16047_);
  nand (_16087_, _16086_, _05049_);
  and (_16088_, _16087_, _06278_);
  nor (_16089_, _16088_, _16083_);
  and (_16090_, _08441_, _04143_);
  nor (_16091_, _16090_, _16047_);
  and (_16092_, _16091_, _02018_);
  nor (_16093_, _16092_, _16089_);
  and (_16094_, _16093_, _02136_);
  and (_16095_, _08304_, _04143_);
  nor (_16097_, _16095_, _16047_);
  nor (_16098_, _16097_, _02136_);
  or (_16099_, _16098_, _16094_);
  and (_16100_, _16099_, _05076_);
  nor (_16101_, _16047_, _05737_);
  not (_16102_, _16101_);
  nor (_16103_, _16086_, _05076_);
  and (_16104_, _16103_, _16102_);
  nor (_16105_, _16104_, _16100_);
  nor (_16106_, _16105_, _02130_);
  or (_16108_, _16101_, _02131_);
  nor (_16109_, _16108_, _16049_);
  or (_16110_, _16109_, _02016_);
  nor (_16111_, _16110_, _16106_);
  nor (_16112_, _08440_, _05963_);
  nor (_16113_, _16112_, _16047_);
  and (_16114_, _16113_, _02016_);
  nor (_16115_, _16114_, _16111_);
  and (_16116_, _16115_, _05474_);
  nor (_16117_, _08303_, _05963_);
  nor (_16119_, _16117_, _16047_);
  nor (_16120_, _16119_, _05474_);
  or (_16121_, _16120_, _16116_);
  and (_16122_, _16121_, _02168_);
  nand (_16123_, _16056_, _01595_);
  and (_16124_, _16123_, _02266_);
  nor (_16125_, _16124_, _16122_);
  and (_16126_, _08507_, _04143_);
  nor (_16127_, _16126_, _16047_);
  and (_16128_, _16127_, _01594_);
  nor (_16130_, _16128_, _16125_);
  or (_16131_, _16130_, _26506_);
  or (_16132_, _26505_, \oc8051_golden_model_1.TL0 [3]);
  and (_16133_, _16132_, _25964_);
  and (_27890_, _16133_, _16131_);
  not (_16134_, \oc8051_golden_model_1.TL0 [4]);
  nor (_16135_, _04143_, _16134_);
  and (_16136_, _08527_, _04143_);
  nor (_16137_, _16136_, _16135_);
  nor (_16138_, _16137_, _02136_);
  and (_16140_, _04143_, _05524_);
  nor (_16141_, _16140_, _16135_);
  and (_16142_, _16141_, _02019_);
  nor (_16143_, _05963_, _04024_);
  nor (_16144_, _16143_, _16135_);
  and (_16145_, _16144_, _04950_);
  and (_16146_, _04143_, \oc8051_golden_model_1.ACC [4]);
  nor (_16147_, _16146_, _16135_);
  nor (_16148_, _16147_, _05488_);
  nor (_16149_, _04571_, _16134_);
  or (_16151_, _16149_, _16148_);
  and (_16152_, _16151_, _02438_);
  nor (_16153_, _08548_, _05963_);
  nor (_16154_, _16153_, _16135_);
  nor (_16155_, _16154_, _02438_);
  or (_16156_, _16155_, _16152_);
  and (_16157_, _16156_, _05487_);
  nor (_16158_, _16144_, _05487_);
  nor (_16159_, _16158_, _16157_);
  nor (_16160_, _16159_, _01963_);
  nor (_16161_, _16147_, _01964_);
  nor (_16162_, _16161_, _04950_);
  not (_16163_, _16162_);
  nor (_16164_, _16163_, _16160_);
  nor (_16165_, _16164_, _16145_);
  nor (_16166_, _16165_, _04951_);
  and (_16167_, _04143_, _03903_);
  nor (_16168_, _16135_, _05513_);
  not (_16169_, _16168_);
  nor (_16170_, _16169_, _16167_);
  or (_16173_, _16170_, _01602_);
  nor (_16174_, _16173_, _16166_);
  nor (_16175_, _08663_, _05963_);
  nor (_16176_, _16175_, _16135_);
  nor (_16177_, _16176_, _01923_);
  or (_16178_, _16177_, _02019_);
  nor (_16179_, _16178_, _16174_);
  nor (_16180_, _16179_, _16142_);
  or (_16181_, _16180_, _02018_);
  and (_16182_, _08531_, _04143_);
  or (_16184_, _16182_, _16135_);
  or (_16185_, _16184_, _05049_);
  and (_16186_, _16185_, _02136_);
  and (_16187_, _16186_, _16181_);
  nor (_16188_, _16187_, _16138_);
  nor (_16189_, _16188_, _02039_);
  nor (_16190_, _16135_, _08729_);
  not (_16191_, _16190_);
  nor (_16192_, _16141_, _05076_);
  and (_16193_, _16192_, _16191_);
  nor (_16195_, _16193_, _16189_);
  nor (_16196_, _16195_, _02130_);
  or (_16197_, _16190_, _02131_);
  nor (_16198_, _16197_, _16147_);
  or (_16199_, _16198_, _02016_);
  nor (_16200_, _16199_, _16196_);
  nor (_16201_, _08530_, _05963_);
  nor (_16202_, _16201_, _16135_);
  and (_16203_, _16202_, _02016_);
  nor (_16204_, _16203_, _16200_);
  and (_16206_, _16204_, _05474_);
  nor (_16207_, _08526_, _05963_);
  nor (_16208_, _16207_, _16135_);
  nor (_16209_, _16208_, _05474_);
  or (_16210_, _16209_, _16206_);
  and (_16211_, _16210_, _02168_);
  nor (_16212_, _16154_, _02168_);
  or (_16213_, _16212_, _01594_);
  nor (_16214_, _16213_, _16211_);
  and (_16215_, _08732_, _04143_);
  nor (_16217_, _16215_, _16135_);
  and (_16218_, _16217_, _01594_);
  nor (_16219_, _16218_, _16214_);
  or (_16220_, _16219_, _26506_);
  or (_16221_, _26505_, \oc8051_golden_model_1.TL0 [4]);
  and (_16222_, _16221_, _25964_);
  and (_27891_, _16222_, _16220_);
  not (_16223_, \oc8051_golden_model_1.TL0 [5]);
  nor (_16224_, _04143_, _16223_);
  and (_16225_, _08750_, _04143_);
  nor (_16227_, _16225_, _16224_);
  nor (_16228_, _16227_, _02136_);
  and (_16229_, _04143_, _05548_);
  nor (_16230_, _16229_, _16224_);
  and (_16231_, _16230_, _02019_);
  nor (_16232_, _05963_, _03976_);
  nor (_16233_, _16232_, _16224_);
  and (_16234_, _16233_, _04950_);
  and (_16235_, _04143_, \oc8051_golden_model_1.ACC [5]);
  nor (_16236_, _16235_, _16224_);
  nor (_16238_, _16236_, _01964_);
  nor (_16239_, _16236_, _05488_);
  nor (_16240_, _04571_, _16223_);
  or (_16241_, _16240_, _16239_);
  and (_16242_, _16241_, _02438_);
  nor (_16243_, _08771_, _05963_);
  nor (_16244_, _16243_, _16224_);
  nor (_16245_, _16244_, _02438_);
  or (_16246_, _16245_, _16242_);
  and (_16247_, _16246_, _05487_);
  nor (_16249_, _16233_, _05487_);
  nor (_16250_, _16249_, _16247_);
  nor (_16251_, _16250_, _01963_);
  or (_16252_, _16251_, _04950_);
  nor (_16253_, _16252_, _16238_);
  nor (_16254_, _16253_, _16234_);
  nor (_16255_, _16254_, _04951_);
  and (_16256_, _04143_, _03850_);
  nor (_16257_, _16224_, _05513_);
  not (_16258_, _16257_);
  nor (_16260_, _16258_, _16256_);
  or (_16261_, _16260_, _01602_);
  nor (_16262_, _16261_, _16255_);
  nor (_16263_, _08874_, _05963_);
  nor (_16264_, _16263_, _16224_);
  nor (_16265_, _16264_, _01923_);
  or (_16266_, _16265_, _02019_);
  nor (_16267_, _16266_, _16262_);
  nor (_16268_, _16267_, _16231_);
  or (_16269_, _16268_, _02018_);
  and (_16271_, _08890_, _04143_);
  or (_16272_, _16271_, _16224_);
  or (_16273_, _16272_, _05049_);
  and (_16274_, _16273_, _02136_);
  and (_16275_, _16274_, _16269_);
  nor (_16276_, _16275_, _16228_);
  nor (_16277_, _16276_, _02039_);
  nor (_16278_, _16224_, _08946_);
  not (_16279_, _16278_);
  nor (_16280_, _16230_, _05076_);
  and (_16282_, _16280_, _16279_);
  nor (_16283_, _16282_, _16277_);
  nor (_16284_, _16283_, _02130_);
  or (_16285_, _16278_, _02131_);
  nor (_16286_, _16285_, _16236_);
  or (_16287_, _16286_, _02016_);
  nor (_16288_, _16287_, _16284_);
  nor (_16289_, _08889_, _05963_);
  nor (_16290_, _16289_, _16224_);
  and (_16291_, _16290_, _02016_);
  nor (_16293_, _16291_, _16288_);
  and (_16294_, _16293_, _05474_);
  nor (_16295_, _08749_, _05963_);
  nor (_16296_, _16295_, _16224_);
  nor (_16297_, _16296_, _05474_);
  or (_16298_, _16297_, _16294_);
  and (_16299_, _16298_, _02168_);
  nor (_16300_, _16244_, _02168_);
  or (_16301_, _16300_, _01594_);
  nor (_16302_, _16301_, _16299_);
  and (_16304_, _08949_, _04143_);
  nor (_16305_, _16304_, _16224_);
  and (_16306_, _16305_, _01594_);
  nor (_16307_, _16306_, _16302_);
  or (_16308_, _16307_, _26506_);
  or (_16309_, _26505_, \oc8051_golden_model_1.TL0 [5]);
  and (_16310_, _16309_, _25964_);
  and (_27892_, _16310_, _16308_);
  not (_16311_, \oc8051_golden_model_1.TL0 [6]);
  nor (_16312_, _04143_, _16311_);
  nor (_16314_, _16312_, _05735_);
  not (_16315_, _16314_);
  and (_16316_, _04143_, _09103_);
  nor (_16317_, _16316_, _16312_);
  nor (_16318_, _16317_, _05076_);
  and (_16319_, _16318_, _16315_);
  and (_16320_, _08975_, _04143_);
  nor (_16321_, _16320_, _16312_);
  nor (_16322_, _16321_, _02136_);
  and (_16323_, _04143_, _03748_);
  or (_16325_, _16323_, _16312_);
  and (_16326_, _16325_, _04951_);
  and (_16327_, _04143_, \oc8051_golden_model_1.ACC [6]);
  nor (_16328_, _16327_, _16312_);
  nor (_16329_, _16328_, _05488_);
  nor (_16330_, _04571_, _16311_);
  or (_16331_, _16330_, _16329_);
  and (_16332_, _16331_, _02438_);
  nor (_16333_, _08995_, _05963_);
  nor (_16334_, _16333_, _16312_);
  nor (_16336_, _16334_, _02438_);
  or (_16337_, _16336_, _16332_);
  and (_16338_, _16337_, _05487_);
  nor (_16339_, _05963_, _04074_);
  nor (_16340_, _16339_, _16312_);
  nor (_16341_, _16340_, _05487_);
  nor (_16342_, _16341_, _16338_);
  nor (_16343_, _16342_, _01963_);
  nor (_16344_, _16328_, _01964_);
  nor (_16345_, _16344_, _04950_);
  not (_16347_, _16345_);
  nor (_16348_, _16347_, _16343_);
  and (_16349_, _16340_, _04950_);
  or (_16350_, _16349_, _04951_);
  nor (_16351_, _16350_, _16348_);
  or (_16352_, _16351_, _16326_);
  and (_16353_, _16352_, _01923_);
  nor (_16354_, _09096_, _05963_);
  nor (_16355_, _16354_, _16312_);
  nor (_16356_, _16355_, _01923_);
  or (_16358_, _16356_, _06278_);
  or (_16359_, _16358_, _16353_);
  and (_16360_, _09112_, _04143_);
  or (_16361_, _16312_, _05049_);
  or (_16362_, _16361_, _16360_);
  and (_16363_, _16317_, _02019_);
  nor (_16364_, _16363_, _02135_);
  and (_16365_, _16364_, _16362_);
  and (_16366_, _16365_, _16359_);
  nor (_16367_, _16366_, _16322_);
  nor (_16369_, _16367_, _02039_);
  nor (_16370_, _16369_, _16319_);
  nor (_16371_, _16370_, _02130_);
  or (_16372_, _16314_, _02131_);
  nor (_16373_, _16372_, _16328_);
  or (_16374_, _16373_, _02016_);
  nor (_16375_, _16374_, _16371_);
  nor (_16376_, _09111_, _05963_);
  nor (_16377_, _16376_, _16312_);
  and (_16378_, _16377_, _02016_);
  nor (_16380_, _16378_, _16375_);
  and (_16381_, _16380_, _05474_);
  nor (_16382_, _08974_, _05963_);
  nor (_16383_, _16382_, _16312_);
  nor (_16384_, _16383_, _05474_);
  or (_16385_, _16384_, _16381_);
  and (_16386_, _16385_, _02168_);
  nor (_16387_, _16334_, _02168_);
  or (_16388_, _16387_, _01594_);
  nor (_16389_, _16388_, _16386_);
  and (_16391_, _08965_, _04143_);
  nor (_16392_, _16391_, _16312_);
  and (_16393_, _16392_, _01594_);
  nor (_16394_, _16393_, _16389_);
  or (_16395_, _16394_, _26506_);
  or (_16396_, _26505_, \oc8051_golden_model_1.TL0 [6]);
  and (_16397_, _16396_, _25964_);
  and (_27893_, _16397_, _16395_);
  not (_16398_, \oc8051_golden_model_1.TL1 [0]);
  nor (_16399_, _04147_, _16398_);
  nor (_16401_, _04405_, _05800_);
  nor (_16402_, _16401_, _16399_);
  and (_16403_, _16402_, _02266_);
  and (_16404_, _04147_, \oc8051_golden_model_1.ACC [0]);
  nor (_16405_, _16404_, _16399_);
  nor (_16406_, _16405_, _01964_);
  nor (_16407_, _16406_, _04950_);
  nor (_16408_, _16402_, _02438_);
  nor (_16409_, _04571_, _16398_);
  nor (_16410_, _16405_, _05488_);
  nor (_16412_, _16410_, _16409_);
  nor (_16413_, _16412_, _01969_);
  or (_16414_, _16413_, _01967_);
  nor (_16415_, _16414_, _16408_);
  or (_16416_, _16415_, _01963_);
  and (_16417_, _16416_, _16407_);
  and (_16418_, _04147_, _03334_);
  or (_16419_, _16399_, _11952_);
  nor (_16420_, _16419_, _16418_);
  nor (_16421_, _16420_, _16417_);
  nor (_16423_, _16421_, _04951_);
  and (_16424_, _04147_, _03677_);
  nor (_16425_, _16399_, _05513_);
  not (_16426_, _16425_);
  nor (_16427_, _16426_, _16424_);
  nor (_16428_, _16427_, _16423_);
  nor (_16429_, _16428_, _01602_);
  nor (_16430_, _07815_, _05800_);
  or (_16431_, _16399_, _01923_);
  nor (_16432_, _16431_, _16430_);
  or (_16434_, _16432_, _02019_);
  nor (_16435_, _16434_, _16429_);
  and (_16436_, _04147_, _05531_);
  nor (_16437_, _16436_, _16399_);
  nand (_16438_, _16437_, _05049_);
  and (_16439_, _16438_, _06278_);
  nor (_16440_, _16439_, _16435_);
  and (_16441_, _07829_, _04147_);
  nor (_16442_, _16441_, _16399_);
  and (_16443_, _16442_, _02018_);
  nor (_16445_, _16443_, _16440_);
  and (_16446_, _16445_, _02136_);
  and (_16447_, _07834_, _04147_);
  nor (_16448_, _16447_, _16399_);
  nor (_16449_, _16448_, _02136_);
  or (_16450_, _16449_, _16446_);
  and (_16451_, _16450_, _05076_);
  or (_16452_, _16437_, _05076_);
  nor (_16453_, _16452_, _16401_);
  nor (_16454_, _16453_, _16451_);
  nor (_16456_, _16454_, _02130_);
  and (_16457_, _07833_, _04147_);
  or (_16458_, _16457_, _16399_);
  and (_16459_, _16458_, _02130_);
  or (_16460_, _16459_, _16456_);
  and (_16461_, _16460_, _05104_);
  nor (_16462_, _07828_, _05800_);
  nor (_16463_, _16462_, _16399_);
  nor (_16464_, _16463_, _05104_);
  or (_16465_, _16464_, _16461_);
  and (_16467_, _16465_, _05474_);
  nor (_16468_, _07696_, _05800_);
  nor (_16469_, _16468_, _16399_);
  nor (_16470_, _16469_, _05474_);
  nor (_16471_, _16470_, _02266_);
  not (_16472_, _16471_);
  nor (_16473_, _16472_, _16467_);
  nor (_16474_, _16473_, _16403_);
  or (_16475_, _16474_, _26506_);
  or (_16476_, _26505_, \oc8051_golden_model_1.TL1 [0]);
  and (_16478_, _16476_, _25964_);
  and (_27896_, _16478_, _16475_);
  nor (_16479_, _04147_, \oc8051_golden_model_1.TL1 [1]);
  and (_16480_, _07909_, _04147_);
  nor (_16481_, _16480_, _16479_);
  nor (_16482_, _16481_, _02168_);
  not (_16483_, _16479_);
  nor (_16484_, _08029_, _05800_);
  nor (_16485_, _16484_, _02136_);
  and (_16486_, _16485_, _16483_);
  and (_16487_, _04147_, _03613_);
  not (_16488_, \oc8051_golden_model_1.TL1 [1]);
  nor (_16489_, _04147_, _16488_);
  nor (_16490_, _16489_, _05513_);
  not (_16491_, _16490_);
  nor (_16492_, _16491_, _16487_);
  not (_16493_, _16492_);
  and (_16494_, _04147_, _01705_);
  nor (_16495_, _16494_, _16479_);
  and (_16496_, _16495_, _01963_);
  and (_16499_, _16495_, _04571_);
  nor (_16500_, _04571_, _16488_);
  or (_16501_, _16500_, _16499_);
  and (_16502_, _16501_, _02438_);
  and (_16503_, _16481_, _01969_);
  or (_16504_, _16503_, _16502_);
  and (_16505_, _16504_, _05487_);
  nor (_16506_, _05800_, _03393_);
  nor (_16507_, _16506_, _16489_);
  nor (_16508_, _16507_, _05487_);
  nor (_16510_, _16508_, _16505_);
  nor (_16511_, _16510_, _01963_);
  or (_16512_, _16511_, _04950_);
  nor (_16513_, _16512_, _16496_);
  and (_16514_, _16507_, _04950_);
  nor (_16515_, _16514_, _16513_);
  nor (_16516_, _16515_, _04951_);
  nor (_16517_, _16516_, _01602_);
  and (_16518_, _16517_, _16493_);
  and (_16519_, _08009_, _04147_);
  nor (_16521_, _16519_, _01923_);
  and (_16522_, _16521_, _16483_);
  nor (_16523_, _16522_, _16518_);
  nor (_16524_, _16523_, _06278_);
  nor (_16525_, _08023_, _05800_);
  nor (_16526_, _16525_, _05049_);
  and (_16527_, _04147_, _02676_);
  nor (_16528_, _16527_, _04979_);
  or (_16529_, _16528_, _16526_);
  and (_16530_, _16529_, _16483_);
  nor (_16532_, _16530_, _16524_);
  nor (_16533_, _16532_, _02135_);
  nor (_16534_, _16533_, _16486_);
  nor (_16535_, _16534_, _02039_);
  nor (_16536_, _07893_, _05800_);
  nor (_16537_, _16536_, _05076_);
  and (_16538_, _16537_, _16483_);
  nor (_16539_, _16538_, _16535_);
  nor (_16540_, _16539_, _02130_);
  nor (_16541_, _16489_, _05741_);
  nor (_16543_, _16541_, _02131_);
  and (_16544_, _16543_, _16495_);
  nor (_16545_, _16544_, _16540_);
  nor (_16546_, _16545_, _02128_);
  and (_16547_, _16527_, _04452_);
  nor (_16548_, _16547_, _05104_);
  nand (_16549_, _16494_, _04452_);
  and (_16550_, _16549_, _02126_);
  or (_16551_, _16550_, _16548_);
  and (_16552_, _16551_, _16483_);
  or (_16554_, _16552_, _02164_);
  nor (_16555_, _16554_, _16546_);
  nor (_16556_, _16555_, _16482_);
  nor (_16557_, _16556_, _01594_);
  nor (_16558_, _16489_, _16480_);
  and (_16559_, _16558_, _01594_);
  nor (_16560_, _16559_, _16557_);
  or (_16561_, _16560_, _26506_);
  or (_16562_, _26505_, \oc8051_golden_model_1.TL1 [1]);
  and (_16563_, _16562_, _25964_);
  and (_27897_, _16563_, _16561_);
  not (_16565_, \oc8051_golden_model_1.TL1 [2]);
  nor (_16566_, _04147_, _16565_);
  nor (_16567_, _16566_, _05739_);
  not (_16568_, _16567_);
  and (_16569_, _04147_, _05563_);
  nor (_16570_, _16569_, _16566_);
  nor (_16571_, _16570_, _05076_);
  and (_16572_, _16571_, _16568_);
  and (_16573_, _04147_, _03564_);
  nor (_16575_, _16573_, _16566_);
  or (_16576_, _16575_, _05513_);
  and (_16577_, _04147_, \oc8051_golden_model_1.ACC [2]);
  nor (_16578_, _16577_, _16566_);
  nor (_16579_, _16578_, _01964_);
  nor (_16580_, _16578_, _05488_);
  nor (_16581_, _04571_, _16565_);
  or (_16582_, _16581_, _16580_);
  and (_16583_, _16582_, _02438_);
  nor (_16584_, _08095_, _05800_);
  nor (_16586_, _16584_, _16566_);
  nor (_16587_, _16586_, _02438_);
  or (_16588_, _16587_, _16583_);
  and (_16589_, _16588_, _05487_);
  nor (_16590_, _05800_, _03272_);
  nor (_16591_, _16590_, _16566_);
  nor (_16592_, _16591_, _05487_);
  nor (_16593_, _16592_, _16589_);
  nor (_16594_, _16593_, _01963_);
  or (_16595_, _16594_, _04950_);
  nor (_16597_, _16595_, _16579_);
  and (_16598_, _16591_, _04950_);
  or (_16599_, _16598_, _04951_);
  or (_16600_, _16599_, _16597_);
  and (_16601_, _16600_, _01923_);
  and (_16602_, _16601_, _16576_);
  nor (_16603_, _08216_, _05800_);
  or (_16604_, _16566_, _01923_);
  nor (_16605_, _16604_, _16603_);
  or (_16606_, _16605_, _02019_);
  nor (_16608_, _16606_, _16602_);
  nand (_16609_, _16570_, _05049_);
  and (_16610_, _16609_, _06278_);
  nor (_16611_, _16610_, _16608_);
  and (_16612_, _08230_, _04147_);
  nor (_16613_, _16612_, _16566_);
  and (_16614_, _16613_, _02018_);
  nor (_16615_, _16614_, _16611_);
  and (_16616_, _16615_, _02136_);
  and (_16617_, _08237_, _04147_);
  nor (_16619_, _16617_, _16566_);
  nor (_16620_, _16619_, _02136_);
  or (_16621_, _16620_, _16616_);
  and (_16622_, _16621_, _05076_);
  nor (_16623_, _16622_, _16572_);
  nor (_16624_, _16623_, _02130_);
  or (_16625_, _16567_, _02131_);
  nor (_16626_, _16625_, _16578_);
  or (_16627_, _16626_, _02016_);
  nor (_16628_, _16627_, _16624_);
  nor (_16630_, _08229_, _05800_);
  nor (_16631_, _16630_, _16566_);
  and (_16632_, _16631_, _02016_);
  nor (_16633_, _16632_, _16628_);
  and (_16634_, _16633_, _05474_);
  nor (_16635_, _08236_, _05800_);
  nor (_16636_, _16635_, _16566_);
  nor (_16637_, _16636_, _05474_);
  or (_16638_, _16637_, _16634_);
  and (_16639_, _16638_, _02168_);
  nor (_16641_, _16586_, _02168_);
  or (_16642_, _16641_, _01594_);
  nor (_16643_, _16642_, _16639_);
  and (_16644_, _08285_, _04147_);
  nor (_16645_, _16644_, _16566_);
  and (_16646_, _16645_, _01594_);
  nor (_16647_, _16646_, _16643_);
  or (_16648_, _16647_, _26506_);
  or (_16649_, _26505_, \oc8051_golden_model_1.TL1 [2]);
  and (_16650_, _16649_, _25964_);
  and (_27898_, _16650_, _16648_);
  not (_16652_, \oc8051_golden_model_1.TL1 [3]);
  nor (_16653_, _04147_, _16652_);
  nor (_16654_, _16653_, _05737_);
  not (_16655_, _16654_);
  and (_16656_, _04147_, _05529_);
  nor (_16657_, _16656_, _16653_);
  nor (_16658_, _16657_, _05076_);
  and (_16659_, _16658_, _16655_);
  and (_16660_, _04147_, \oc8051_golden_model_1.ACC [3]);
  nor (_16662_, _16660_, _16653_);
  nor (_16663_, _16662_, _05488_);
  nor (_16664_, _04571_, _16652_);
  or (_16665_, _16664_, _16663_);
  and (_16666_, _16665_, _02438_);
  nor (_16667_, _08337_, _05800_);
  nor (_16668_, _16667_, _16653_);
  nor (_16669_, _16668_, _02438_);
  or (_16670_, _16669_, _16666_);
  and (_16671_, _16670_, _05487_);
  nor (_16673_, _05800_, _03473_);
  nor (_16674_, _16673_, _16653_);
  nor (_16675_, _16674_, _05487_);
  nor (_16676_, _16675_, _16671_);
  nor (_16677_, _16676_, _01963_);
  nor (_16678_, _16662_, _01964_);
  nor (_16679_, _16678_, _04950_);
  not (_16680_, _16679_);
  nor (_16681_, _16680_, _16677_);
  and (_16682_, _16674_, _04950_);
  or (_16684_, _16682_, _04951_);
  or (_16685_, _16684_, _16681_);
  and (_16686_, _04147_, _03516_);
  nor (_16687_, _16686_, _16653_);
  or (_16688_, _16687_, _05513_);
  and (_16689_, _16688_, _01923_);
  and (_16690_, _16689_, _16685_);
  nor (_16691_, _08425_, _05800_);
  or (_16692_, _16653_, _01923_);
  nor (_16693_, _16692_, _16691_);
  or (_16695_, _16693_, _02019_);
  nor (_16696_, _16695_, _16690_);
  nand (_16697_, _16657_, _05049_);
  and (_16698_, _16697_, _06278_);
  nor (_16699_, _16698_, _16696_);
  and (_16700_, _08441_, _04147_);
  nor (_16701_, _16700_, _16653_);
  and (_16702_, _16701_, _02018_);
  nor (_16703_, _16702_, _16699_);
  and (_16704_, _16703_, _02136_);
  and (_16706_, _08304_, _04147_);
  nor (_16707_, _16706_, _16653_);
  nor (_16708_, _16707_, _02136_);
  or (_16709_, _16708_, _16704_);
  and (_16710_, _16709_, _05076_);
  nor (_16711_, _16710_, _16659_);
  nor (_16712_, _16711_, _02130_);
  or (_16713_, _16654_, _02131_);
  nor (_16714_, _16713_, _16662_);
  or (_16715_, _16714_, _02016_);
  nor (_16717_, _16715_, _16712_);
  nor (_16718_, _08440_, _05800_);
  nor (_16719_, _16718_, _16653_);
  and (_16720_, _16719_, _02016_);
  nor (_16721_, _16720_, _16717_);
  and (_16722_, _16721_, _05474_);
  nor (_16723_, _08303_, _05800_);
  nor (_16724_, _16723_, _16653_);
  nor (_16725_, _16724_, _05474_);
  or (_16726_, _16725_, _16722_);
  and (_16728_, _16726_, _02168_);
  nor (_16729_, _16668_, _02168_);
  or (_16730_, _16729_, _01594_);
  nor (_16731_, _16730_, _16728_);
  and (_16732_, _08507_, _04147_);
  nor (_16733_, _16732_, _16653_);
  and (_16734_, _16733_, _01594_);
  nor (_16735_, _16734_, _16731_);
  or (_16736_, _16735_, _26506_);
  or (_16737_, _26505_, \oc8051_golden_model_1.TL1 [3]);
  and (_16739_, _16737_, _25964_);
  and (_27899_, _16739_, _16736_);
  not (_16740_, \oc8051_golden_model_1.TL1 [4]);
  nor (_16741_, _04147_, _16740_);
  and (_16742_, _08527_, _04147_);
  nor (_16743_, _16742_, _16741_);
  nor (_16744_, _16743_, _02136_);
  and (_16745_, _04147_, _05524_);
  nor (_16746_, _16745_, _16741_);
  and (_16747_, _16746_, _02019_);
  nor (_16749_, _05800_, _04024_);
  nor (_16750_, _16749_, _16741_);
  and (_16751_, _16750_, _04950_);
  and (_16752_, _04147_, \oc8051_golden_model_1.ACC [4]);
  nor (_16753_, _16752_, _16741_);
  nor (_16754_, _16753_, _05488_);
  nor (_16755_, _04571_, _16740_);
  or (_16756_, _16755_, _16754_);
  and (_16757_, _16756_, _02438_);
  nor (_16758_, _08548_, _05800_);
  nor (_16760_, _16758_, _16741_);
  nor (_16761_, _16760_, _02438_);
  or (_16762_, _16761_, _16757_);
  and (_16763_, _16762_, _05487_);
  nor (_16764_, _16750_, _05487_);
  nor (_16765_, _16764_, _16763_);
  nor (_16766_, _16765_, _01963_);
  nor (_16767_, _16753_, _01964_);
  nor (_16768_, _16767_, _04950_);
  not (_16769_, _16768_);
  nor (_16771_, _16769_, _16766_);
  nor (_16772_, _16771_, _16751_);
  nor (_16773_, _16772_, _04951_);
  and (_16774_, _04147_, _03903_);
  nor (_16775_, _16741_, _05513_);
  not (_16776_, _16775_);
  nor (_16777_, _16776_, _16774_);
  or (_16778_, _16777_, _01602_);
  nor (_16779_, _16778_, _16773_);
  nor (_16780_, _08663_, _05800_);
  nor (_16782_, _16780_, _16741_);
  nor (_16783_, _16782_, _01923_);
  or (_16784_, _16783_, _02019_);
  nor (_16785_, _16784_, _16779_);
  nor (_16786_, _16785_, _16747_);
  or (_16787_, _16786_, _02018_);
  and (_16788_, _08531_, _04147_);
  or (_16789_, _16788_, _16741_);
  or (_16790_, _16789_, _05049_);
  and (_16791_, _16790_, _02136_);
  and (_16793_, _16791_, _16787_);
  nor (_16794_, _16793_, _16744_);
  nor (_16795_, _16794_, _02039_);
  nor (_16796_, _16741_, _08729_);
  not (_16797_, _16796_);
  nor (_16798_, _16746_, _05076_);
  and (_16799_, _16798_, _16797_);
  nor (_16800_, _16799_, _16795_);
  nor (_16801_, _16800_, _02130_);
  or (_16802_, _16796_, _02131_);
  nor (_16804_, _16802_, _16753_);
  or (_16805_, _16804_, _02016_);
  nor (_16806_, _16805_, _16801_);
  nor (_16807_, _08530_, _05800_);
  nor (_16808_, _16807_, _16741_);
  and (_16809_, _16808_, _02016_);
  nor (_16810_, _16809_, _16806_);
  and (_16811_, _16810_, _05474_);
  nor (_16812_, _08526_, _05800_);
  nor (_16813_, _16812_, _16741_);
  nor (_16815_, _16813_, _05474_);
  or (_16816_, _16815_, _16811_);
  and (_16817_, _16816_, _02168_);
  nor (_16818_, _16760_, _02168_);
  or (_16819_, _16818_, _01594_);
  nor (_16820_, _16819_, _16817_);
  and (_16821_, _08732_, _04147_);
  nor (_16822_, _16821_, _16741_);
  and (_16823_, _16822_, _01594_);
  nor (_16824_, _16823_, _16820_);
  or (_16826_, _16824_, _26506_);
  or (_16827_, _26505_, \oc8051_golden_model_1.TL1 [4]);
  and (_16828_, _16827_, _25964_);
  and (_27900_, _16828_, _16826_);
  not (_16829_, \oc8051_golden_model_1.TL1 [5]);
  nor (_16830_, _04147_, _16829_);
  and (_16831_, _08750_, _04147_);
  nor (_16832_, _16831_, _16830_);
  nor (_16833_, _16832_, _02136_);
  and (_16834_, _04147_, _05548_);
  nor (_16836_, _16834_, _16830_);
  and (_16837_, _16836_, _02019_);
  and (_16838_, _04147_, \oc8051_golden_model_1.ACC [5]);
  nor (_16839_, _16838_, _16830_);
  nor (_16840_, _16839_, _01964_);
  nor (_16841_, _16839_, _05488_);
  nor (_16842_, _04571_, _16829_);
  or (_16843_, _16842_, _16841_);
  and (_16844_, _16843_, _02438_);
  nor (_16845_, _08771_, _05800_);
  nor (_16847_, _16845_, _16830_);
  nor (_16848_, _16847_, _02438_);
  or (_16849_, _16848_, _16844_);
  and (_16850_, _16849_, _05487_);
  nor (_16851_, _05800_, _03976_);
  nor (_16852_, _16851_, _16830_);
  nor (_16853_, _16852_, _05487_);
  nor (_16854_, _16853_, _16850_);
  nor (_16855_, _16854_, _01963_);
  or (_16856_, _16855_, _04950_);
  nor (_16857_, _16856_, _16840_);
  and (_16858_, _16852_, _04950_);
  nor (_16859_, _16858_, _16857_);
  nor (_16860_, _16859_, _04951_);
  and (_16861_, _04147_, _03850_);
  nor (_16862_, _16830_, _05513_);
  not (_16863_, _16862_);
  nor (_16864_, _16863_, _16861_);
  or (_16865_, _16864_, _01602_);
  nor (_16866_, _16865_, _16860_);
  nor (_16869_, _08874_, _05800_);
  nor (_16870_, _16869_, _16830_);
  nor (_16871_, _16870_, _01923_);
  or (_16872_, _16871_, _02019_);
  nor (_16873_, _16872_, _16866_);
  nor (_16874_, _16873_, _16837_);
  or (_16875_, _16874_, _02018_);
  and (_16876_, _08890_, _04147_);
  or (_16877_, _16876_, _16830_);
  or (_16878_, _16877_, _05049_);
  and (_16880_, _16878_, _02136_);
  and (_16881_, _16880_, _16875_);
  nor (_16882_, _16881_, _16833_);
  nor (_16883_, _16882_, _02039_);
  nor (_16884_, _16830_, _08946_);
  not (_16885_, _16884_);
  nor (_16886_, _16836_, _05076_);
  and (_16887_, _16886_, _16885_);
  nor (_16888_, _16887_, _16883_);
  nor (_16889_, _16888_, _02130_);
  or (_16891_, _16884_, _02131_);
  nor (_16892_, _16891_, _16839_);
  or (_16893_, _16892_, _02016_);
  nor (_16894_, _16893_, _16889_);
  nor (_16895_, _08889_, _05800_);
  nor (_16896_, _16895_, _16830_);
  and (_16897_, _16896_, _02016_);
  nor (_16898_, _16897_, _16894_);
  and (_16899_, _16898_, _05474_);
  nor (_16900_, _08749_, _05800_);
  nor (_16902_, _16900_, _16830_);
  nor (_16903_, _16902_, _05474_);
  or (_16904_, _16903_, _16899_);
  and (_16905_, _16904_, _02168_);
  nor (_16906_, _16847_, _02168_);
  or (_16907_, _16906_, _01594_);
  nor (_16908_, _16907_, _16905_);
  and (_16909_, _08949_, _04147_);
  nor (_16910_, _16909_, _16830_);
  and (_16911_, _16910_, _01594_);
  nor (_16913_, _16911_, _16908_);
  or (_16914_, _16913_, _26506_);
  or (_16915_, _26505_, \oc8051_golden_model_1.TL1 [5]);
  and (_16916_, _16915_, _25964_);
  and (_27901_, _16916_, _16914_);
  not (_16917_, \oc8051_golden_model_1.TL1 [6]);
  nor (_16918_, _04147_, _16917_);
  and (_16919_, _08975_, _04147_);
  nor (_16920_, _16919_, _16918_);
  nor (_16921_, _16920_, _02136_);
  and (_16923_, _04147_, _03748_);
  or (_16924_, _16923_, _16918_);
  and (_16925_, _16924_, _04951_);
  and (_16926_, _04147_, \oc8051_golden_model_1.ACC [6]);
  nor (_16927_, _16926_, _16918_);
  nor (_16928_, _16927_, _01964_);
  nor (_16929_, _16927_, _05488_);
  nor (_16930_, _04571_, _16917_);
  or (_16931_, _16930_, _16929_);
  and (_16932_, _16931_, _02438_);
  nor (_16934_, _08995_, _05800_);
  nor (_16935_, _16934_, _16918_);
  nor (_16936_, _16935_, _02438_);
  or (_16937_, _16936_, _16932_);
  and (_16938_, _16937_, _05487_);
  nor (_16939_, _05800_, _04074_);
  nor (_16940_, _16939_, _16918_);
  nor (_16941_, _16940_, _05487_);
  nor (_16942_, _16941_, _16938_);
  nor (_16943_, _16942_, _01963_);
  or (_16945_, _16943_, _04950_);
  nor (_16946_, _16945_, _16928_);
  and (_16947_, _16940_, _04950_);
  or (_16948_, _16947_, _04951_);
  nor (_16949_, _16948_, _16946_);
  or (_16950_, _16949_, _16925_);
  and (_16951_, _16950_, _01923_);
  nor (_16952_, _09096_, _05800_);
  nor (_16953_, _16952_, _16918_);
  nor (_16954_, _16953_, _01923_);
  or (_16956_, _16954_, _06278_);
  or (_16957_, _16956_, _16951_);
  and (_16958_, _09112_, _04147_);
  or (_16959_, _16918_, _05049_);
  or (_16960_, _16959_, _16958_);
  and (_16961_, _04147_, _09103_);
  nor (_16962_, _16961_, _16918_);
  and (_16963_, _16962_, _02019_);
  nor (_16964_, _16963_, _02135_);
  and (_16965_, _16964_, _16960_);
  and (_16967_, _16965_, _16957_);
  nor (_16968_, _16967_, _16921_);
  nor (_16969_, _16968_, _02039_);
  nor (_16970_, _16918_, _05735_);
  not (_16971_, _16970_);
  nor (_16972_, _16962_, _05076_);
  and (_16973_, _16972_, _16971_);
  nor (_16974_, _16973_, _16969_);
  nor (_16975_, _16974_, _02130_);
  or (_16976_, _16970_, _02131_);
  nor (_16978_, _16976_, _16927_);
  or (_16979_, _16978_, _02016_);
  nor (_16980_, _16979_, _16975_);
  nor (_16981_, _09111_, _05800_);
  nor (_16982_, _16981_, _16918_);
  and (_16983_, _16982_, _02016_);
  nor (_16984_, _16983_, _16980_);
  and (_16985_, _16984_, _05474_);
  nor (_16986_, _08974_, _05800_);
  nor (_16987_, _16986_, _16918_);
  nor (_16989_, _16987_, _05474_);
  or (_16990_, _16989_, _16985_);
  and (_16991_, _16990_, _02168_);
  nor (_16992_, _16935_, _02168_);
  or (_16993_, _16992_, _01594_);
  nor (_16994_, _16993_, _16991_);
  and (_16995_, _08965_, _04147_);
  nor (_16996_, _16995_, _16918_);
  and (_16997_, _16996_, _01594_);
  nor (_16998_, _16997_, _16994_);
  or (_17000_, _16998_, _26506_);
  or (_17001_, _26505_, \oc8051_golden_model_1.TL1 [6]);
  and (_17002_, _17001_, _25964_);
  and (_27902_, _17002_, _17000_);
  not (_17003_, \oc8051_golden_model_1.TMOD [0]);
  nor (_17004_, _04134_, _17003_);
  nor (_17005_, _04405_, _05480_);
  nor (_17006_, _17005_, _17004_);
  and (_17007_, _17006_, _02266_);
  and (_17008_, _04134_, _05531_);
  nor (_17010_, _17008_, _17004_);
  nor (_17011_, _17010_, _05076_);
  not (_17012_, _17011_);
  nor (_17013_, _17012_, _17005_);
  and (_17014_, _04134_, _03334_);
  nor (_17015_, _17014_, _17004_);
  and (_17016_, _17015_, _04950_);
  and (_17017_, _04134_, \oc8051_golden_model_1.ACC [0]);
  nor (_17018_, _17017_, _17004_);
  nor (_17019_, _17018_, _01964_);
  nor (_17021_, _17018_, _05488_);
  nor (_17022_, _04571_, _17003_);
  or (_17023_, _17022_, _17021_);
  and (_17024_, _17023_, _02438_);
  nor (_17025_, _17006_, _02438_);
  or (_17026_, _17025_, _17024_);
  and (_17027_, _17026_, _05487_);
  nor (_17028_, _17015_, _05487_);
  nor (_17029_, _17028_, _17027_);
  nor (_17030_, _17029_, _01963_);
  or (_17032_, _17030_, _04950_);
  nor (_17033_, _17032_, _17019_);
  nor (_17034_, _17033_, _17016_);
  nor (_17035_, _17034_, _04951_);
  and (_17036_, _04134_, _03677_);
  nor (_17037_, _17004_, _05513_);
  not (_17038_, _17037_);
  nor (_17039_, _17038_, _17036_);
  nor (_17040_, _17039_, _17035_);
  nor (_17041_, _17040_, _01602_);
  nor (_17043_, _07815_, _05480_);
  or (_17044_, _17004_, _01923_);
  nor (_17045_, _17044_, _17043_);
  or (_17046_, _17045_, _02019_);
  nor (_17047_, _17046_, _17041_);
  nor (_17048_, _17010_, _04979_);
  or (_17049_, _17048_, _17047_);
  and (_17050_, _17049_, _05049_);
  and (_17051_, _07829_, _04134_);
  nor (_17052_, _17051_, _17004_);
  nor (_17054_, _17052_, _05049_);
  or (_17055_, _17054_, _17050_);
  and (_17056_, _17055_, _02136_);
  and (_17057_, _07834_, _04134_);
  nor (_17058_, _17057_, _17004_);
  nor (_17059_, _17058_, _02136_);
  or (_17060_, _17059_, _17056_);
  and (_17061_, _17060_, _05076_);
  nor (_17062_, _17061_, _17013_);
  nor (_17063_, _17062_, _02130_);
  and (_17065_, _07833_, _04134_);
  or (_17066_, _17065_, _17004_);
  and (_17067_, _17066_, _02130_);
  or (_17068_, _17067_, _17063_);
  and (_17069_, _17068_, _05104_);
  nor (_17070_, _07828_, _05480_);
  nor (_17071_, _17070_, _17004_);
  nor (_17072_, _17071_, _05104_);
  or (_17073_, _17072_, _17069_);
  and (_17074_, _17073_, _05474_);
  nor (_17076_, _07696_, _05480_);
  nor (_17077_, _17076_, _17004_);
  nor (_17078_, _17077_, _05474_);
  nor (_17079_, _17078_, _02266_);
  not (_17080_, _17079_);
  nor (_17081_, _17080_, _17074_);
  nor (_17082_, _17081_, _17007_);
  or (_17083_, _17082_, _26506_);
  or (_17084_, _26505_, \oc8051_golden_model_1.TMOD [0]);
  and (_17085_, _17084_, _25964_);
  and (_27905_, _17085_, _17083_);
  nor (_17087_, _04134_, \oc8051_golden_model_1.TMOD [1]);
  and (_17088_, _07909_, _04134_);
  nor (_17089_, _17088_, _17087_);
  nor (_17090_, _17089_, _02168_);
  not (_17091_, _17087_);
  nor (_17092_, _08029_, _05480_);
  nor (_17093_, _17092_, _02136_);
  and (_17094_, _17093_, _17091_);
  and (_17095_, _04134_, _03613_);
  not (_17097_, \oc8051_golden_model_1.TMOD [1]);
  nor (_17098_, _04134_, _17097_);
  nor (_17099_, _17098_, _05513_);
  not (_17100_, _17099_);
  nor (_17101_, _17100_, _17095_);
  not (_17102_, _17101_);
  nor (_17103_, _05480_, _03393_);
  nor (_17104_, _17103_, _17098_);
  and (_17105_, _17104_, _04950_);
  and (_17106_, _04134_, _01705_);
  nor (_17108_, _17106_, _17087_);
  and (_17109_, _17108_, _01963_);
  and (_17110_, _17108_, _04571_);
  nor (_17111_, _04571_, _17097_);
  or (_17112_, _17111_, _17110_);
  and (_17113_, _17112_, _02438_);
  and (_17114_, _17089_, _01969_);
  or (_17115_, _17114_, _17113_);
  and (_17116_, _17115_, _05487_);
  nor (_17117_, _17104_, _05487_);
  nor (_17119_, _17117_, _17116_);
  nor (_17120_, _17119_, _01963_);
  or (_17121_, _17120_, _04950_);
  nor (_17122_, _17121_, _17109_);
  nor (_17123_, _17122_, _17105_);
  nor (_17124_, _17123_, _04951_);
  nor (_17125_, _17124_, _01602_);
  and (_17126_, _17125_, _17102_);
  and (_17127_, _08009_, _04134_);
  nor (_17128_, _17127_, _01923_);
  and (_17130_, _17128_, _17091_);
  nor (_17131_, _17130_, _17126_);
  nor (_17132_, _17131_, _06278_);
  nor (_17133_, _08023_, _05480_);
  nor (_17134_, _17133_, _05049_);
  and (_17135_, _04134_, _02676_);
  nor (_17136_, _17135_, _04979_);
  or (_17137_, _17136_, _17134_);
  and (_17138_, _17137_, _17091_);
  nor (_17139_, _17138_, _17132_);
  nor (_17141_, _17139_, _02135_);
  nor (_17142_, _17141_, _17094_);
  nor (_17143_, _17142_, _02039_);
  nor (_17144_, _07893_, _05480_);
  nor (_17145_, _17144_, _05076_);
  and (_17146_, _17145_, _17091_);
  nor (_17147_, _17146_, _17143_);
  nor (_17148_, _17147_, _02130_);
  nor (_17149_, _17098_, _05741_);
  nor (_17150_, _17149_, _02131_);
  and (_17152_, _17150_, _17108_);
  nor (_17153_, _17152_, _17148_);
  nor (_17154_, _17153_, _02128_);
  and (_17155_, _17135_, _04452_);
  nor (_17156_, _17155_, _05104_);
  nand (_17157_, _17106_, _04452_);
  and (_17158_, _17157_, _02126_);
  or (_17159_, _17158_, _17156_);
  and (_17160_, _17159_, _17091_);
  or (_17161_, _17160_, _02164_);
  nor (_17163_, _17161_, _17154_);
  nor (_17164_, _17163_, _17090_);
  nor (_17165_, _17164_, _01594_);
  nor (_17166_, _17098_, _17088_);
  and (_17167_, _17166_, _01594_);
  nor (_17168_, _17167_, _17165_);
  or (_17169_, _17168_, _26506_);
  or (_17170_, _26505_, \oc8051_golden_model_1.TMOD [1]);
  and (_17171_, _17170_, _25964_);
  and (_27906_, _17171_, _17169_);
  not (_17173_, \oc8051_golden_model_1.TMOD [2]);
  nor (_17174_, _04134_, _17173_);
  and (_17175_, _04134_, _03564_);
  nor (_17176_, _17175_, _17174_);
  or (_17177_, _17176_, _05513_);
  and (_17178_, _04134_, \oc8051_golden_model_1.ACC [2]);
  nor (_17179_, _17178_, _17174_);
  nor (_17180_, _17179_, _01964_);
  nor (_17181_, _17179_, _05488_);
  nor (_17182_, _04571_, _17173_);
  or (_17184_, _17182_, _17181_);
  and (_17185_, _17184_, _02438_);
  nor (_17186_, _08095_, _05480_);
  nor (_17187_, _17186_, _17174_);
  nor (_17188_, _17187_, _02438_);
  or (_17189_, _17188_, _17185_);
  and (_17190_, _17189_, _05487_);
  nor (_17191_, _05480_, _03272_);
  nor (_17192_, _17191_, _17174_);
  nor (_17193_, _17192_, _05487_);
  nor (_17195_, _17193_, _17190_);
  nor (_17196_, _17195_, _01963_);
  or (_17197_, _17196_, _04950_);
  nor (_17198_, _17197_, _17180_);
  and (_17199_, _17192_, _04950_);
  or (_17200_, _17199_, _04951_);
  or (_17201_, _17200_, _17198_);
  and (_17202_, _17201_, _01923_);
  and (_17203_, _17202_, _17177_);
  nor (_17204_, _08216_, _05480_);
  or (_17206_, _17174_, _01923_);
  nor (_17207_, _17206_, _17204_);
  or (_17208_, _17207_, _02019_);
  nor (_17209_, _17208_, _17203_);
  and (_17210_, _04134_, _05563_);
  nor (_17211_, _17210_, _17174_);
  nor (_17212_, _17211_, _04979_);
  or (_17213_, _17212_, _17209_);
  and (_17214_, _17213_, _05049_);
  and (_17215_, _08230_, _04134_);
  nor (_17216_, _17215_, _17174_);
  nor (_17217_, _17216_, _05049_);
  or (_17218_, _17217_, _17214_);
  and (_17219_, _17218_, _02136_);
  and (_17220_, _08237_, _04134_);
  nor (_17221_, _17220_, _17174_);
  nor (_17222_, _17221_, _02136_);
  or (_17223_, _17222_, _17219_);
  and (_17224_, _17223_, _05076_);
  nor (_17225_, _17174_, _05739_);
  or (_17227_, _17211_, _05076_);
  nor (_17228_, _17227_, _17225_);
  nor (_17229_, _17228_, _17224_);
  nor (_17230_, _17229_, _02130_);
  or (_17231_, _17225_, _02131_);
  nor (_17232_, _17231_, _17179_);
  or (_17233_, _17232_, _02016_);
  nor (_17234_, _17233_, _17230_);
  nor (_17235_, _08229_, _05480_);
  nor (_17236_, _17235_, _17174_);
  and (_17238_, _17236_, _02016_);
  nor (_17239_, _17238_, _17234_);
  and (_17240_, _17239_, _05474_);
  nor (_17241_, _08236_, _05480_);
  nor (_17242_, _17241_, _17174_);
  nor (_17243_, _17242_, _05474_);
  or (_17244_, _17243_, _17240_);
  and (_17245_, _17244_, _02168_);
  nor (_17246_, _17187_, _02168_);
  or (_17247_, _17246_, _01594_);
  nor (_17249_, _17247_, _17245_);
  and (_17250_, _08285_, _04134_);
  nor (_17251_, _17250_, _17174_);
  and (_17252_, _17251_, _01594_);
  nor (_17253_, _17252_, _17249_);
  or (_17254_, _17253_, _26506_);
  or (_17255_, _26505_, \oc8051_golden_model_1.TMOD [2]);
  and (_17256_, _17255_, _25964_);
  and (_27907_, _17256_, _17254_);
  not (_17257_, \oc8051_golden_model_1.TMOD [3]);
  nor (_17259_, _04134_, _17257_);
  and (_17260_, _08304_, _04134_);
  nor (_17261_, _17260_, _17259_);
  nor (_17262_, _17261_, _02136_);
  and (_17263_, _04134_, _03516_);
  or (_17264_, _17263_, _17259_);
  and (_17265_, _17264_, _04951_);
  and (_17266_, _04134_, \oc8051_golden_model_1.ACC [3]);
  nor (_17267_, _17266_, _17259_);
  nor (_17268_, _17267_, _01964_);
  nor (_17270_, _17267_, _05488_);
  nor (_17271_, _04571_, _17257_);
  or (_17272_, _17271_, _17270_);
  and (_17273_, _17272_, _02438_);
  nor (_17274_, _08337_, _05480_);
  nor (_17275_, _17274_, _17259_);
  nor (_17276_, _17275_, _02438_);
  or (_17277_, _17276_, _17273_);
  and (_17278_, _17277_, _05487_);
  nor (_17279_, _05480_, _03473_);
  nor (_17281_, _17279_, _17259_);
  nor (_17282_, _17281_, _05487_);
  nor (_17283_, _17282_, _17278_);
  nor (_17284_, _17283_, _01963_);
  or (_17285_, _17284_, _04950_);
  nor (_17286_, _17285_, _17268_);
  and (_17287_, _17281_, _04950_);
  or (_17288_, _17287_, _04951_);
  nor (_17289_, _17288_, _17286_);
  or (_17290_, _17289_, _17265_);
  and (_17292_, _17290_, _01923_);
  nor (_17293_, _08425_, _05480_);
  nor (_17294_, _17293_, _17259_);
  nor (_17295_, _17294_, _01923_);
  or (_17296_, _17295_, _06278_);
  or (_17297_, _17296_, _17292_);
  and (_17298_, _08441_, _04134_);
  or (_17299_, _17259_, _05049_);
  or (_17300_, _17299_, _17298_);
  and (_17301_, _04134_, _05529_);
  nor (_17303_, _17301_, _17259_);
  and (_17304_, _17303_, _02019_);
  nor (_17305_, _17304_, _02135_);
  and (_17306_, _17305_, _17300_);
  and (_17307_, _17306_, _17297_);
  nor (_17308_, _17307_, _17262_);
  nor (_17309_, _17308_, _02039_);
  nor (_17310_, _17259_, _05737_);
  not (_17311_, _17310_);
  nor (_17312_, _17303_, _05076_);
  and (_17314_, _17312_, _17311_);
  nor (_17315_, _17314_, _17309_);
  nor (_17316_, _17315_, _02130_);
  or (_17317_, _17310_, _02131_);
  nor (_17318_, _17317_, _17267_);
  or (_17319_, _17318_, _02016_);
  nor (_17320_, _17319_, _17316_);
  nor (_17321_, _08440_, _05480_);
  nor (_17322_, _17321_, _17259_);
  and (_17323_, _17322_, _02016_);
  nor (_17325_, _17323_, _17320_);
  and (_17326_, _17325_, _05474_);
  nor (_17327_, _08303_, _05480_);
  nor (_17328_, _17327_, _17259_);
  nor (_17329_, _17328_, _05474_);
  or (_17330_, _17329_, _17326_);
  and (_17331_, _17330_, _02168_);
  nor (_17332_, _17275_, _02168_);
  or (_17333_, _17332_, _01594_);
  nor (_17334_, _17333_, _17331_);
  and (_17336_, _08507_, _04134_);
  nor (_17337_, _17336_, _17259_);
  and (_17338_, _17337_, _01594_);
  nor (_17339_, _17338_, _17334_);
  or (_17340_, _17339_, _26506_);
  or (_17341_, _26505_, \oc8051_golden_model_1.TMOD [3]);
  and (_17342_, _17341_, _25964_);
  and (_27908_, _17342_, _17340_);
  not (_17343_, \oc8051_golden_model_1.TMOD [4]);
  nor (_17344_, _04134_, _17343_);
  and (_17346_, _08527_, _04134_);
  nor (_17347_, _17346_, _17344_);
  nor (_17348_, _17347_, _02136_);
  and (_17349_, _04134_, _05524_);
  nor (_17350_, _17349_, _17344_);
  and (_17351_, _17350_, _02019_);
  nor (_17352_, _05480_, _04024_);
  nor (_17353_, _17352_, _17344_);
  and (_17354_, _17353_, _04950_);
  and (_17355_, _04134_, \oc8051_golden_model_1.ACC [4]);
  nor (_17356_, _17355_, _17344_);
  nor (_17357_, _17356_, _01964_);
  nor (_17358_, _17356_, _05488_);
  nor (_17359_, _04571_, _17343_);
  or (_17360_, _17359_, _17358_);
  and (_17361_, _17360_, _02438_);
  nor (_17362_, _08548_, _05480_);
  nor (_17363_, _17362_, _17344_);
  nor (_17364_, _17363_, _02438_);
  or (_17365_, _17364_, _17361_);
  and (_17367_, _17365_, _05487_);
  nor (_17368_, _17353_, _05487_);
  nor (_17369_, _17368_, _17367_);
  nor (_17370_, _17369_, _01963_);
  or (_17371_, _17370_, _04950_);
  nor (_17372_, _17371_, _17357_);
  nor (_17373_, _17372_, _17354_);
  nor (_17374_, _17373_, _04951_);
  and (_17375_, _04134_, _03903_);
  nor (_17376_, _17344_, _05513_);
  not (_17378_, _17376_);
  nor (_17379_, _17378_, _17375_);
  or (_17380_, _17379_, _01602_);
  nor (_17381_, _17380_, _17374_);
  nor (_17382_, _08663_, _05480_);
  nor (_17383_, _17382_, _17344_);
  nor (_17384_, _17383_, _01923_);
  or (_17385_, _17384_, _02019_);
  nor (_17386_, _17385_, _17381_);
  nor (_17387_, _17386_, _17351_);
  or (_17389_, _17387_, _02018_);
  and (_17390_, _08531_, _04134_);
  or (_17391_, _17390_, _17344_);
  or (_17392_, _17391_, _05049_);
  and (_17393_, _17392_, _02136_);
  and (_17394_, _17393_, _17389_);
  nor (_17395_, _17394_, _17348_);
  nor (_17396_, _17395_, _02039_);
  nor (_17397_, _17344_, _08729_);
  not (_17398_, _17397_);
  nor (_17400_, _17350_, _05076_);
  and (_17401_, _17400_, _17398_);
  nor (_17402_, _17401_, _17396_);
  nor (_17403_, _17402_, _02130_);
  or (_17404_, _17397_, _02131_);
  nor (_17405_, _17404_, _17356_);
  or (_17406_, _17405_, _02016_);
  nor (_17407_, _17406_, _17403_);
  nor (_17408_, _08530_, _05480_);
  nor (_17409_, _17408_, _17344_);
  and (_17411_, _17409_, _02016_);
  nor (_17412_, _17411_, _17407_);
  and (_17413_, _17412_, _05474_);
  nor (_17414_, _08526_, _05480_);
  nor (_17415_, _17414_, _17344_);
  nor (_17416_, _17415_, _05474_);
  or (_17417_, _17416_, _17413_);
  and (_17418_, _17417_, _02168_);
  nor (_17419_, _17363_, _02168_);
  or (_17420_, _17419_, _01594_);
  nor (_17422_, _17420_, _17418_);
  and (_17423_, _08732_, _04134_);
  nor (_17424_, _17423_, _17344_);
  and (_17425_, _17424_, _01594_);
  nor (_17426_, _17425_, _17422_);
  or (_17427_, _17426_, _26506_);
  or (_17428_, _26505_, \oc8051_golden_model_1.TMOD [4]);
  and (_17429_, _17428_, _25964_);
  and (_27909_, _17429_, _17427_);
  not (_17430_, \oc8051_golden_model_1.TMOD [5]);
  nor (_17432_, _04134_, _17430_);
  and (_17433_, _08750_, _04134_);
  nor (_17434_, _17433_, _17432_);
  nor (_17435_, _17434_, _02136_);
  nor (_17436_, _08874_, _05480_);
  or (_17437_, _17432_, _01923_);
  or (_17438_, _17437_, _17436_);
  nor (_17439_, _08771_, _05480_);
  nor (_17440_, _17439_, _17432_);
  nor (_17441_, _17440_, _02438_);
  nor (_17443_, _04571_, _17430_);
  and (_17444_, _04134_, \oc8051_golden_model_1.ACC [5]);
  nor (_17445_, _17444_, _17432_);
  nor (_17446_, _17445_, _05488_);
  nor (_17447_, _17446_, _17443_);
  nor (_17448_, _17447_, _01969_);
  or (_17449_, _17448_, _17441_);
  and (_17450_, _17449_, _05487_);
  nor (_17451_, _05480_, _03976_);
  nor (_17452_, _17451_, _17432_);
  nor (_17454_, _17452_, _05487_);
  or (_17455_, _17454_, _17450_);
  and (_17456_, _17455_, _01964_);
  nor (_17457_, _17445_, _01964_);
  nor (_17458_, _17457_, _04950_);
  not (_17459_, _17458_);
  nor (_17460_, _17459_, _17456_);
  and (_17461_, _17452_, _04950_);
  or (_17462_, _17461_, _04951_);
  nor (_17463_, _17462_, _17460_);
  and (_17465_, _04134_, _03850_);
  or (_17466_, _17465_, _17432_);
  and (_17467_, _17466_, _04951_);
  or (_17468_, _17467_, _01602_);
  or (_17469_, _17468_, _17463_);
  and (_17470_, _17469_, _17438_);
  and (_17471_, _17470_, _04979_);
  and (_17472_, _04134_, _05548_);
  nor (_17473_, _17472_, _17432_);
  nor (_17474_, _17473_, _04979_);
  or (_17476_, _17474_, _17471_);
  or (_17477_, _17476_, _02018_);
  and (_17478_, _08890_, _04134_);
  or (_17479_, _17478_, _17432_);
  or (_17480_, _17479_, _05049_);
  and (_17481_, _17480_, _02136_);
  and (_17482_, _17481_, _17477_);
  nor (_17483_, _17482_, _17435_);
  nor (_17484_, _17483_, _02039_);
  nor (_17485_, _17432_, _08946_);
  not (_17487_, _17485_);
  nor (_17488_, _17473_, _05076_);
  and (_17489_, _17488_, _17487_);
  nor (_17490_, _17489_, _17484_);
  nor (_17491_, _17490_, _02130_);
  or (_17492_, _17485_, _02131_);
  nor (_17493_, _17492_, _17445_);
  or (_17494_, _17493_, _02016_);
  nor (_17495_, _17494_, _17491_);
  nor (_17496_, _08889_, _05480_);
  nor (_17498_, _17496_, _17432_);
  and (_17499_, _17498_, _02016_);
  nor (_17500_, _17499_, _17495_);
  and (_17501_, _17500_, _05474_);
  nor (_17502_, _08749_, _05480_);
  nor (_17503_, _17502_, _17432_);
  nor (_17504_, _17503_, _05474_);
  or (_17505_, _17504_, _17501_);
  and (_17506_, _17505_, _02168_);
  nor (_17507_, _17440_, _02168_);
  or (_17509_, _17507_, _01594_);
  nor (_17510_, _17509_, _17506_);
  and (_17511_, _08949_, _04134_);
  nor (_17512_, _17511_, _17432_);
  and (_17513_, _17512_, _01594_);
  nor (_17514_, _17513_, _17510_);
  or (_17515_, _17514_, _26506_);
  or (_17516_, _26505_, \oc8051_golden_model_1.TMOD [5]);
  and (_17517_, _17516_, _25964_);
  and (_27910_, _17517_, _17515_);
  not (_17519_, \oc8051_golden_model_1.TMOD [6]);
  nor (_17520_, _04134_, _17519_);
  and (_17521_, _08975_, _04134_);
  nor (_17522_, _17521_, _17520_);
  nor (_17523_, _17522_, _02136_);
  and (_17524_, _04134_, _03748_);
  or (_17525_, _17524_, _17520_);
  and (_17526_, _17525_, _04951_);
  and (_17527_, _04134_, \oc8051_golden_model_1.ACC [6]);
  nor (_17528_, _17527_, _17520_);
  nor (_17530_, _17528_, _01964_);
  nor (_17531_, _17528_, _05488_);
  nor (_17532_, _04571_, _17519_);
  or (_17533_, _17532_, _17531_);
  and (_17534_, _17533_, _02438_);
  nor (_17535_, _08995_, _05480_);
  nor (_17536_, _17535_, _17520_);
  nor (_17537_, _17536_, _02438_);
  or (_17538_, _17537_, _17534_);
  and (_17539_, _17538_, _05487_);
  nor (_17541_, _05480_, _04074_);
  nor (_17542_, _17541_, _17520_);
  nor (_17543_, _17542_, _05487_);
  nor (_17544_, _17543_, _17539_);
  nor (_17545_, _17544_, _01963_);
  or (_17546_, _17545_, _04950_);
  nor (_17547_, _17546_, _17530_);
  and (_17548_, _17542_, _04950_);
  or (_17549_, _17548_, _04951_);
  nor (_17550_, _17549_, _17547_);
  or (_17551_, _17550_, _17526_);
  and (_17552_, _17551_, _01923_);
  nor (_17553_, _09096_, _05480_);
  nor (_17554_, _17553_, _17520_);
  nor (_17555_, _17554_, _01923_);
  or (_17556_, _17555_, _06278_);
  or (_17557_, _17556_, _17552_);
  and (_17558_, _09112_, _04134_);
  or (_17559_, _17520_, _05049_);
  or (_17560_, _17559_, _17558_);
  and (_17562_, _04134_, _09103_);
  nor (_17563_, _17562_, _17520_);
  and (_17564_, _17563_, _02019_);
  nor (_17565_, _17564_, _02135_);
  and (_17566_, _17565_, _17560_);
  and (_17567_, _17566_, _17557_);
  nor (_17568_, _17567_, _17523_);
  nor (_17569_, _17568_, _02039_);
  nor (_17570_, _17520_, _05735_);
  not (_17571_, _17570_);
  nor (_17573_, _17563_, _05076_);
  and (_17574_, _17573_, _17571_);
  nor (_17575_, _17574_, _17569_);
  nor (_17576_, _17575_, _02130_);
  or (_17577_, _17570_, _02131_);
  nor (_17578_, _17577_, _17528_);
  or (_17579_, _17578_, _02016_);
  nor (_17580_, _17579_, _17576_);
  nor (_17581_, _09111_, _05480_);
  nor (_17582_, _17581_, _17520_);
  and (_17584_, _17582_, _02016_);
  nor (_17585_, _17584_, _17580_);
  and (_17586_, _17585_, _05474_);
  nor (_17587_, _08974_, _05480_);
  nor (_17588_, _17587_, _17520_);
  nor (_17589_, _17588_, _05474_);
  or (_17590_, _17589_, _17586_);
  and (_17591_, _17590_, _02168_);
  nor (_17592_, _17536_, _02168_);
  or (_17593_, _17592_, _01594_);
  nor (_17595_, _17593_, _17591_);
  and (_17596_, _08965_, _04134_);
  nor (_17597_, _17596_, _17520_);
  and (_17598_, _17597_, _01594_);
  nor (_17599_, _17598_, _17595_);
  or (_17600_, _17599_, _26506_);
  or (_17601_, _26505_, \oc8051_golden_model_1.TMOD [6]);
  and (_17602_, _17601_, _25964_);
  and (_27911_, _17602_, _17600_);
  nor (_17603_, _02026_, _01657_);
  not (_17605_, _17603_);
  and (_17606_, _17605_, _02516_);
  and (_17607_, _05457_, _05445_);
  nor (_17608_, _17607_, _01325_);
  and (_17609_, _05397_, _02818_);
  nor (_17610_, _17609_, _01325_);
  not (_17611_, _01663_);
  nor (_17612_, _05097_, _02016_);
  nor (_17613_, _17612_, _01325_);
  not (_17614_, _01666_);
  nor (_17615_, _05069_, _02039_);
  nor (_17616_, _17615_, _01325_);
  not (_17617_, _01653_);
  and (_17618_, _02830_, _05049_);
  nor (_17619_, _17618_, _01325_);
  and (_17620_, _02019_, _01325_);
  nor (_17621_, _02516_, _01632_);
  and (_17622_, _03909_, _01325_);
  and (_17623_, _02516_, \oc8051_golden_model_1.PC [0]);
  nor (_17624_, _17623_, _03117_);
  not (_17627_, _17624_);
  nor (_17628_, _17627_, _03909_);
  or (_17629_, _17628_, _17622_);
  nor (_17630_, _17629_, _03187_);
  and (_17631_, _04085_, _01325_);
  nor (_17632_, _17627_, _04085_);
  or (_17633_, _17632_, _17631_);
  nor (_17634_, _17633_, _04090_);
  nor (_17635_, _04734_, _04725_);
  nor (_17636_, _17635_, _01325_);
  not (_17638_, _01630_);
  and (_17639_, _04715_, _01325_);
  and (_17640_, _04710_, \oc8051_golden_model_1.PC [0]);
  and (_17641_, _02409_, _01325_);
  nor (_17642_, _17641_, _04648_);
  and (_17643_, _17642_, _04707_);
  or (_17644_, _17643_, _04709_);
  nor (_17645_, _17644_, _17640_);
  nor (_17646_, _02516_, _01628_);
  nor (_17647_, _04564_, _01325_);
  nor (_17649_, _17647_, _04558_);
  and (_17650_, _04561_, _01325_);
  nor (_17651_, _04561_, _01325_);
  nor (_17652_, _17651_, _17650_);
  and (_17653_, _17652_, _01625_);
  or (_17654_, _17653_, _04567_);
  and (_17655_, _17654_, _17649_);
  or (_17656_, _17655_, _04557_);
  nor (_17657_, _17656_, _17646_);
  or (_17658_, _17657_, _04715_);
  nor (_17660_, _17658_, _17645_);
  or (_17661_, _17660_, _17639_);
  and (_17662_, _17661_, _02438_);
  not (_17663_, _17662_);
  and (_17664_, _04553_, _01325_);
  and (_17665_, _17624_, _04551_);
  nor (_17666_, _17665_, _17664_);
  nor (_17667_, _17666_, _02438_);
  nor (_17668_, _17667_, _04094_);
  and (_17669_, _17668_, _17663_);
  and (_17671_, _04094_, \oc8051_golden_model_1.PC [0]);
  nor (_17672_, _17671_, _06363_);
  not (_17673_, _17672_);
  nor (_17674_, _17673_, _17669_);
  nor (_17675_, _02516_, _01621_);
  not (_17676_, _17635_);
  nor (_17677_, _17676_, _17675_);
  not (_17678_, _17677_);
  nor (_17679_, _17678_, _17674_);
  or (_17680_, _17679_, _17638_);
  nor (_17682_, _17680_, _17636_);
  nor (_17683_, _02516_, _01630_);
  nor (_17684_, _17683_, _04089_);
  not (_17685_, _17684_);
  nor (_17686_, _17685_, _17682_);
  nor (_17687_, _17686_, _17634_);
  nor (_17688_, _17687_, _03185_);
  or (_17689_, _17688_, _01951_);
  nor (_17690_, _17689_, _17630_);
  and (_17691_, _04874_, _01325_);
  nor (_17693_, _17627_, _04874_);
  nor (_17694_, _17693_, _17691_);
  nor (_17695_, _17694_, _02378_);
  nor (_17696_, _17695_, _17690_);
  nor (_17697_, _17696_, _03179_);
  and (_17698_, _02912_, \oc8051_golden_model_1.PC [0]);
  nor (_17699_, _17624_, _02912_);
  or (_17700_, _17699_, _04749_);
  nor (_17701_, _17700_, _17698_);
  or (_17702_, _17701_, _17697_);
  and (_17704_, _17702_, _02881_);
  and (_17705_, _02880_, _01325_);
  or (_17706_, _17705_, _17704_);
  and (_17707_, _17706_, _01632_);
  or (_17708_, _17707_, _04908_);
  nor (_17709_, _17708_, _17621_);
  not (_17710_, _01618_);
  nor (_17711_, _04905_, _01325_);
  nor (_17712_, _17711_, _17710_);
  not (_17713_, _17712_);
  nor (_17715_, _17713_, _17709_);
  nor (_17716_, _02516_, _01618_);
  and (_17717_, _04928_, _01616_);
  not (_17718_, _17717_);
  nor (_17719_, _17718_, _17716_);
  not (_17720_, _17719_);
  nor (_17721_, _17720_, _17715_);
  nor (_17722_, _17717_, _01325_);
  nor (_17723_, _17722_, _01606_);
  not (_17724_, _17723_);
  nor (_17726_, _17724_, _17721_);
  nor (_17727_, _02516_, _07270_);
  nor (_17728_, _04960_, _01602_);
  and (_17729_, _17728_, _02002_);
  not (_17730_, _17729_);
  nor (_17731_, _17730_, _17727_);
  not (_17732_, _17731_);
  nor (_17733_, _17732_, _17726_);
  nor (_17734_, _17729_, _01325_);
  nor (_17735_, _17734_, _01654_);
  not (_17737_, _17735_);
  nor (_17738_, _17737_, _17733_);
  not (_17739_, _01654_);
  nor (_17740_, _02516_, _17739_);
  or (_17741_, _17740_, _04968_);
  nor (_17742_, _17741_, _17738_);
  nor (_17743_, _17642_, _04969_);
  nor (_17744_, _17743_, _17742_);
  and (_17745_, _17744_, _04979_);
  or (_17746_, _17745_, _17620_);
  and (_17747_, _17746_, _04985_);
  and (_17748_, _04984_, _01614_);
  or (_17749_, _17748_, _17747_);
  and (_17750_, _17749_, _01651_);
  nor (_17751_, _02516_, _01651_);
  or (_17752_, _17751_, _17750_);
  and (_17753_, _17752_, _05027_);
  not (_17754_, _17618_);
  nor (_17755_, _17642_, _05038_);
  and (_17756_, _05038_, _01325_);
  nor (_17758_, _17756_, _05027_);
  not (_17759_, _17758_);
  nor (_17760_, _17759_, _17755_);
  nor (_17761_, _17760_, _17754_);
  not (_17762_, _17761_);
  nor (_17763_, _17762_, _17753_);
  nor (_17764_, _17763_, _17619_);
  and (_17765_, _17764_, _17617_);
  nor (_17766_, _02516_, _17617_);
  or (_17767_, _17766_, _17765_);
  and (_17769_, _17767_, _05060_);
  not (_17770_, _17615_);
  nor (_17771_, _05038_, _01325_);
  and (_17772_, _17642_, _05038_);
  or (_17773_, _17772_, _17771_);
  and (_17774_, _17773_, _05059_);
  nor (_17775_, _17774_, _17770_);
  not (_17776_, _17775_);
  nor (_17777_, _17776_, _17769_);
  nor (_17778_, _17777_, _17616_);
  and (_17780_, _17778_, _17614_);
  nor (_17781_, _02516_, _17614_);
  or (_17782_, _17781_, _17780_);
  and (_17783_, _17782_, _05087_);
  not (_17784_, _17612_);
  nor (_17785_, _17642_, \oc8051_golden_model_1.PSW [7]);
  and (_17786_, \oc8051_golden_model_1.PSW [7], _01325_);
  nor (_17787_, _17786_, _05087_);
  not (_17788_, _17787_);
  nor (_17789_, _17788_, _17785_);
  nor (_17791_, _17789_, _17784_);
  not (_17792_, _17791_);
  nor (_17793_, _17792_, _17783_);
  nor (_17794_, _17793_, _17613_);
  and (_17795_, _17794_, _17611_);
  nor (_17796_, _02516_, _17611_);
  or (_17797_, _17796_, _17795_);
  and (_17798_, _17797_, _05115_);
  and (_17799_, _05092_, \oc8051_golden_model_1.PC [0]);
  and (_17800_, _17642_, \oc8051_golden_model_1.PSW [7]);
  or (_17802_, _17800_, _17799_);
  and (_17803_, _17802_, _05114_);
  and (_17804_, _05139_, _05146_);
  not (_17805_, _17804_);
  nor (_17806_, _17805_, _17803_);
  not (_17807_, _17806_);
  nor (_17808_, _17807_, _17798_);
  nor (_17809_, _17804_, _01325_);
  or (_17810_, _17809_, _02146_);
  nor (_17811_, _17810_, _17808_);
  and (_17813_, _03677_, _02146_);
  or (_17814_, _17813_, _17811_);
  and (_17815_, _17814_, _05157_);
  nor (_17816_, _02516_, _05157_);
  or (_17817_, _17816_, _17815_);
  and (_17818_, _17817_, _02153_);
  not (_17819_, _17609_);
  and (_17820_, _17627_, _05386_);
  nor (_17821_, _05386_, _01325_);
  or (_17822_, _17821_, _02153_);
  nor (_17824_, _17822_, _17820_);
  nor (_17825_, _17824_, _17819_);
  not (_17826_, _17825_);
  nor (_17827_, _17826_, _17818_);
  nor (_17828_, _17827_, _17610_);
  and (_17829_, _17828_, _01596_);
  and (_17830_, _03677_, _01585_);
  or (_17831_, _17830_, _17829_);
  and (_17832_, _17831_, _05407_);
  nor (_17833_, _02516_, _05407_);
  or (_17835_, _17833_, _02022_);
  or (_17836_, _17835_, _17832_);
  and (_17837_, _05430_, _05418_);
  and (_17838_, _05386_, \oc8051_golden_model_1.PC [0]);
  nor (_17839_, _17624_, _05386_);
  nor (_17840_, _17839_, _17838_);
  or (_17841_, _17840_, _02558_);
  and (_17842_, _17841_, _17837_);
  and (_17843_, _17842_, _17836_);
  nor (_17844_, _17837_, \oc8051_golden_model_1.PC [0]);
  nor (_17846_, _17844_, _06467_);
  not (_17847_, _17846_);
  nor (_17848_, _17847_, _17843_);
  and (_17849_, _06467_, _02516_);
  nor (_17850_, _17849_, _02025_);
  not (_17851_, _17850_);
  nor (_17852_, _17851_, _17848_);
  not (_17853_, _17607_);
  and (_17854_, _17840_, _02025_);
  nor (_17855_, _17854_, _17853_);
  not (_17857_, _17855_);
  nor (_17858_, _17857_, _17852_);
  nor (_17859_, _17858_, _17608_);
  nor (_17860_, _17605_, _17859_);
  or (_17861_, _17860_, _05464_);
  nor (_17862_, _17861_, _17606_);
  and (_17863_, _05464_, _01325_);
  nor (_17864_, _17863_, _17862_);
  nand (_17865_, _17864_, _26505_);
  or (_17866_, _26505_, \oc8051_golden_model_1.PC [0]);
  and (_17868_, _17866_, _25964_);
  and (_27914_, _17868_, _17865_);
  and (_17869_, _03115_, _05464_);
  not (_17870_, _17869_);
  and (_17871_, _01594_, _01298_);
  and (_17872_, _05386_, _03115_);
  nor (_17873_, _03119_, _03117_);
  nor (_17874_, _17873_, _03120_);
  nor (_17875_, _17874_, _05386_);
  nor (_17876_, _17875_, _17872_);
  and (_17878_, _17876_, _02025_);
  and (_17879_, _02164_, _01298_);
  and (_17880_, _02032_, _01580_);
  and (_17881_, _02032_, _01659_);
  and (_17882_, _05097_, _01690_);
  and (_17883_, _02032_, _01665_);
  and (_17884_, _04960_, _01690_);
  and (_17885_, _02880_, _01690_);
  and (_17886_, _04085_, _01690_);
  not (_17887_, _17874_);
  nor (_17889_, _17887_, _04085_);
  or (_17890_, _17889_, _17886_);
  nor (_17891_, _17890_, _04090_);
  and (_17892_, _04734_, _01690_);
  nor (_17893_, _02676_, _01627_);
  not (_17894_, _04562_);
  and (_17895_, _02857_, _01970_);
  and (_17896_, _17895_, _01690_);
  or (_17897_, _01626_, _01591_);
  not (_17898_, _17897_);
  and (_17900_, _04559_, _03115_);
  not (_17901_, _04559_);
  and (_17902_, _04560_, \oc8051_golden_model_1.PC [0]);
  nor (_17903_, _17902_, _04571_);
  and (_17904_, _17903_, _01298_);
  nor (_17905_, _17903_, _01298_);
  nor (_17906_, _17905_, _17904_);
  and (_17907_, _17906_, _17901_);
  or (_17908_, _17907_, _17900_);
  and (_17909_, _17908_, _01625_);
  nor (_17911_, _02676_, _01625_);
  nor (_17912_, _17911_, _17909_);
  nor (_17913_, _17912_, _17898_);
  nor (_17914_, _17897_, _01690_);
  nor (_17915_, _17914_, _17895_);
  not (_17916_, _17915_);
  nor (_17917_, _17916_, _17913_);
  or (_17918_, _17917_, _01971_);
  nor (_17919_, _17918_, _17896_);
  and (_17920_, _01971_, _01298_);
  or (_17921_, _17920_, _17919_);
  and (_17922_, _17921_, _17894_);
  and (_17923_, _04562_, _03115_);
  or (_17924_, _17923_, _17922_);
  and (_17925_, _17924_, _01627_);
  or (_17926_, _17925_, _04557_);
  nor (_17927_, _17926_, _17893_);
  or (_17928_, _04707_, \oc8051_golden_model_1.PC [1]);
  nor (_17929_, _04650_, _04648_);
  nor (_17930_, _17929_, _04651_);
  nand (_17932_, _17930_, _04707_);
  and (_17933_, _17932_, _17928_);
  and (_17934_, _17933_, _04557_);
  or (_17935_, _17934_, _17927_);
  nand (_17936_, _17935_, _07515_);
  and (_17937_, _04715_, _01690_);
  nor (_17938_, _17937_, _01969_);
  nand (_17939_, _17938_, _17936_);
  not (_17940_, _04094_);
  or (_17941_, _17874_, _04553_);
  or (_17943_, _04551_, _01690_);
  and (_17944_, _17943_, _01969_);
  nand (_17945_, _17944_, _17941_);
  and (_17946_, _17945_, _17940_);
  nand (_17947_, _17946_, _17939_);
  and (_17948_, _04094_, _01690_);
  nor (_17949_, _17948_, _01959_);
  nand (_17950_, _17949_, _17947_);
  and (_17951_, _01959_, _01298_);
  nor (_17952_, _17951_, _06363_);
  nand (_17954_, _17952_, _17950_);
  and (_17955_, _02676_, _06363_);
  nor (_17956_, _17955_, _01967_);
  nand (_17957_, _17956_, _17954_);
  and (_17958_, _01967_, _01298_);
  nor (_17959_, _17958_, _04725_);
  nand (_17960_, _17959_, _17957_);
  and (_17961_, _04725_, _01690_);
  nor (_17962_, _17961_, _01963_);
  nand (_17963_, _17962_, _17960_);
  and (_17965_, _01963_, _01298_);
  nor (_17966_, _17965_, _04734_);
  and (_17967_, _17966_, _17963_);
  or (_17968_, _17967_, _17892_);
  nand (_17969_, _17968_, _06229_);
  and (_17970_, _01957_, \oc8051_golden_model_1.PC [1]);
  nor (_17971_, _17970_, _17638_);
  and (_17972_, _17971_, _17969_);
  nor (_17973_, _02676_, _01630_);
  or (_17974_, _17973_, _17972_);
  nand (_17976_, _17974_, _02457_);
  and (_17977_, _01953_, _01298_);
  nor (_17978_, _17977_, _04089_);
  and (_17979_, _17978_, _17976_);
  or (_17980_, _17979_, _17891_);
  nand (_17981_, _17980_, _03187_);
  or (_17982_, _17887_, _03909_);
  nand (_17983_, _03909_, _01690_);
  and (_17984_, _17983_, _03185_);
  nand (_17985_, _17984_, _17982_);
  nand (_17987_, _17985_, _17981_);
  nand (_17988_, _17987_, _02378_);
  and (_17989_, _04874_, _01690_);
  not (_17990_, _17989_);
  nor (_17991_, _17887_, _04874_);
  nor (_17992_, _17991_, _02378_);
  and (_17993_, _17992_, _17990_);
  nor (_17994_, _17993_, _03179_);
  nand (_17995_, _17994_, _17988_);
  and (_17996_, _02912_, _03115_);
  nor (_17998_, _17874_, _02912_);
  or (_17999_, _17998_, _04749_);
  or (_18000_, _17999_, _17996_);
  and (_18001_, _18000_, _02881_);
  and (_18002_, _18001_, _17995_);
  or (_18003_, _18002_, _17885_);
  nand (_18004_, _18003_, _04885_);
  and (_18005_, _01946_, \oc8051_golden_model_1.PC [1]);
  nor (_18006_, _18005_, _06393_);
  nand (_18007_, _18006_, _18004_);
  not (_18009_, _04897_);
  nor (_18010_, _02676_, _01632_);
  nor (_18011_, _18010_, _18009_);
  nand (_18012_, _18011_, _18007_);
  nor (_18013_, _04897_, _01298_);
  nor (_18014_, _18013_, _04903_);
  and (_18015_, _18014_, _18012_);
  nor (_18016_, _04904_, _03115_);
  nor (_18017_, _18016_, _04905_);
  or (_18018_, _18017_, _18015_);
  and (_18020_, _04904_, _01690_);
  nor (_18021_, _18020_, _01931_);
  nand (_18022_, _18021_, _18018_);
  and (_18023_, _01931_, _01298_);
  nor (_18024_, _18023_, _17710_);
  nand (_18025_, _18024_, _18022_);
  and (_18026_, _02676_, _17710_);
  nor (_18027_, _18026_, _01930_);
  nand (_18028_, _18027_, _18025_);
  and (_18029_, _01930_, _01298_);
  nor (_18031_, _18029_, _04925_);
  and (_18032_, _18031_, _18028_);
  and (_18033_, _04925_, _01690_);
  or (_18034_, _18033_, _18032_);
  nor (_18035_, _04920_, _04915_);
  nand (_18036_, _18035_, _18034_);
  nor (_18037_, _18035_, _03115_);
  nor (_18038_, _18037_, _04923_);
  nand (_18039_, _18038_, _18036_);
  and (_18040_, _04923_, _03115_);
  nor (_18041_, _18040_, _04932_);
  nand (_18042_, _18041_, _18039_);
  and (_18043_, _04932_, \oc8051_golden_model_1.PC [1]);
  nor (_18044_, _18043_, _01611_);
  nand (_18045_, _18044_, _18042_);
  and (_18046_, _03115_, _01611_);
  nor (_18047_, _18046_, _01924_);
  and (_18048_, _18047_, _18045_);
  and (_18049_, _01924_, \oc8051_golden_model_1.PC [1]);
  or (_18050_, _18049_, _18048_);
  nand (_18053_, _18050_, _07270_);
  and (_18054_, _02676_, _01606_);
  nor (_18055_, _18054_, _02001_);
  nand (_18056_, _18055_, _18053_);
  and (_18057_, _02001_, _01690_);
  nor (_18058_, _18057_, _04953_);
  nand (_18059_, _18058_, _18056_);
  nor (_18060_, _04952_, _01298_);
  nor (_18061_, _18060_, _01602_);
  and (_18062_, _18061_, _18059_);
  nor (_18064_, _04960_, _01690_);
  nor (_18065_, _18064_, _17728_);
  nor (_18066_, _18065_, _18062_);
  or (_18067_, _18066_, _17884_);
  nand (_18068_, _18067_, _02519_);
  and (_18069_, _01920_, \oc8051_golden_model_1.PC [1]);
  nor (_18070_, _18069_, _01654_);
  and (_18071_, _18070_, _18068_);
  nor (_18072_, _02676_, _17739_);
  or (_18073_, _18072_, _18071_);
  nand (_18075_, _18073_, _04969_);
  and (_18076_, _17930_, _04968_);
  nor (_18077_, _18076_, _02859_);
  and (_18078_, _18077_, _18075_);
  nor (_18079_, _02019_, \oc8051_golden_model_1.PC [1]);
  nor (_18080_, _18079_, _07508_);
  or (_18081_, _18080_, _18078_);
  and (_18082_, _02019_, _01690_);
  nor (_18083_, _18082_, _02853_);
  and (_18084_, _18083_, _18081_);
  and (_18085_, _02853_, \oc8051_golden_model_1.PC [1]);
  or (_18086_, _18085_, _18084_);
  nand (_18087_, _18086_, _04985_);
  and (_18088_, _04984_, _01700_);
  nor (_18089_, _18088_, _01919_);
  nand (_18090_, _18089_, _18087_);
  and (_18091_, _01919_, _01298_);
  nor (_18092_, _18091_, _01650_);
  nand (_18093_, _18092_, _18090_);
  and (_18094_, _02676_, _01650_);
  nor (_18096_, _18094_, _05026_);
  nand (_18097_, _18096_, _18093_);
  nand (_18098_, _05038_, _01298_);
  nand (_18099_, _17930_, _05040_);
  and (_18100_, _18099_, _18098_);
  or (_18101_, _18100_, _05027_);
  and (_18102_, _18101_, _18097_);
  or (_18103_, _18102_, _02311_);
  and (_18104_, _02311_, _03115_);
  or (_18105_, _02804_, _02010_);
  or (_18107_, _08712_, _18105_);
  and (_18108_, _18107_, _01652_);
  nor (_18109_, _18108_, _18104_);
  nand (_18110_, _18109_, _18103_);
  and (_18111_, _18108_, _01690_);
  nor (_18112_, _18111_, _02823_);
  nand (_18113_, _18112_, _18110_);
  and (_18114_, _02823_, _03115_);
  nor (_18115_, _18114_, _05047_);
  nand (_18116_, _18115_, _18113_);
  and (_18118_, _05047_, \oc8051_golden_model_1.PC [1]);
  nor (_18119_, _18118_, _02018_);
  nand (_18120_, _18119_, _18116_);
  and (_18121_, _02018_, _01690_);
  nor (_18122_, _18121_, _02135_);
  and (_18123_, _18122_, _18120_);
  and (_18124_, _02135_, \oc8051_golden_model_1.PC [1]);
  or (_18125_, _18124_, _18123_);
  nand (_18126_, _18125_, _17617_);
  and (_18127_, _02676_, _01653_);
  nor (_18129_, _18127_, _05059_);
  and (_18130_, _18129_, _18126_);
  nor (_18131_, _05038_, \oc8051_golden_model_1.PC [1]);
  and (_18132_, _17930_, _05038_);
  or (_18133_, _18132_, _18131_);
  and (_18134_, _18133_, _05059_);
  nor (_18135_, _18134_, _18130_);
  or (_18136_, _18135_, _17883_);
  and (_18137_, _17883_, _03115_);
  nor (_18138_, _02009_, _02531_);
  nor (_18140_, _18138_, _18137_);
  nand (_18141_, _18140_, _18136_);
  and (_18142_, _18138_, _01690_);
  nor (_18143_, _02857_, _04886_);
  nand (_18144_, _18143_, _02695_);
  and (_18145_, _18144_, _01665_);
  nor (_18146_, _18145_, _18142_);
  nand (_18147_, _18146_, _18141_);
  and (_18148_, _18145_, _03115_);
  nor (_18149_, _18148_, _05072_);
  nand (_18151_, _18149_, _18147_);
  and (_18152_, _05072_, \oc8051_golden_model_1.PC [1]);
  nor (_18153_, _18152_, _02039_);
  nand (_18154_, _18153_, _18151_);
  and (_18155_, _02039_, _01690_);
  nor (_18156_, _18155_, _02130_);
  and (_18157_, _18156_, _18154_);
  and (_18158_, _02130_, \oc8051_golden_model_1.PC [1]);
  or (_18159_, _18158_, _18157_);
  nand (_18160_, _18159_, _17614_);
  and (_18162_, _02676_, _01666_);
  nor (_18163_, _18162_, _05086_);
  nand (_18164_, _18163_, _18160_);
  nor (_18165_, _17930_, \oc8051_golden_model_1.PSW [7]);
  and (_18166_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  nor (_18167_, _18166_, _05087_);
  not (_18168_, _18167_);
  nor (_18169_, _18168_, _18165_);
  nor (_18170_, _18169_, _05097_);
  and (_18171_, _18170_, _18164_);
  or (_18173_, _18171_, _17882_);
  nand (_18174_, _18173_, _05105_);
  and (_18175_, _05101_, \oc8051_golden_model_1.PC [1]);
  nor (_18176_, _18175_, _02016_);
  nand (_18177_, _18176_, _18174_);
  and (_18178_, _02016_, _01690_);
  nor (_18179_, _18178_, _02126_);
  and (_18180_, _18179_, _18177_);
  and (_18181_, _02126_, \oc8051_golden_model_1.PC [1]);
  or (_18182_, _18181_, _18180_);
  nand (_18184_, _18182_, _17611_);
  and (_18185_, _02676_, _01663_);
  nor (_18186_, _18185_, _05114_);
  and (_18187_, _18186_, _18184_);
  nor (_18188_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and (_18189_, _17930_, \oc8051_golden_model_1.PSW [7]);
  or (_18190_, _18189_, _18188_);
  and (_18191_, _18190_, _05114_);
  nor (_18192_, _18191_, _18187_);
  or (_18193_, _18192_, _17881_);
  and (_18195_, _17881_, _03115_);
  not (_18196_, _18195_);
  nor (_18197_, _01935_, _01609_);
  and (_18198_, _18197_, _01659_);
  or (_18199_, _18198_, _05131_);
  or (_18200_, _18199_, _02681_);
  or (_18201_, _18200_, _05132_);
  or (_18202_, _18201_, _05136_);
  nor (_18203_, _18202_, _05129_);
  and (_18204_, _18203_, _18196_);
  nand (_18206_, _18204_, _18193_);
  nor (_18207_, _18203_, _03115_);
  nor (_18208_, _18207_, _05124_);
  nand (_18209_, _18208_, _18206_);
  and (_18210_, _05124_, _03115_);
  nor (_18211_, _18210_, _02273_);
  nand (_18212_, _18211_, _18209_);
  and (_18213_, _02273_, \oc8051_golden_model_1.PC [1]);
  nor (_18214_, _18213_, _05145_);
  nand (_18215_, _18214_, _18212_);
  and (_18217_, _05145_, _03115_);
  nor (_18218_, _18217_, _02146_);
  and (_18219_, _18218_, _18215_);
  nor (_18220_, _03613_, _02718_);
  or (_18221_, _18220_, _18219_);
  nand (_18222_, _18221_, _05157_);
  and (_18223_, _02676_, _01660_);
  nor (_18224_, _18223_, _02015_);
  and (_18225_, _18224_, _18222_);
  and (_18226_, _17874_, _05386_);
  nor (_18228_, _05386_, _03115_);
  nor (_18229_, _18228_, _18226_);
  nor (_18230_, _18229_, _02153_);
  nor (_18231_, _18230_, _18225_);
  or (_18232_, _18231_, _17880_);
  and (_18233_, _17880_, _03115_);
  not (_18234_, _18233_);
  or (_18235_, _02446_, _02550_);
  and (_18236_, _18235_, _02809_);
  and (_18237_, _18236_, _18234_);
  nand (_18239_, _18237_, _18232_);
  nor (_18240_, _18236_, _03115_);
  nor (_18241_, _18240_, _02813_);
  nand (_18242_, _18241_, _18239_);
  and (_18243_, _02813_, _03115_);
  nor (_18244_, _18243_, _02788_);
  nand (_18245_, _18244_, _18242_);
  and (_18246_, _02788_, \oc8051_golden_model_1.PC [1]);
  nor (_18247_, _18246_, _05396_);
  nand (_18248_, _18247_, _18245_);
  and (_18250_, _05396_, _03115_);
  nor (_18251_, _18250_, _01585_);
  and (_18252_, _18251_, _18248_);
  nor (_18253_, _03613_, _01596_);
  or (_18254_, _18253_, _18252_);
  nand (_18255_, _18254_, _05407_);
  and (_18256_, _02676_, _01581_);
  nor (_18257_, _18256_, _02022_);
  nand (_18258_, _18257_, _18255_);
  and (_18259_, _17876_, _02022_);
  nor (_18261_, _18259_, _05416_);
  and (_18262_, _18261_, _18258_);
  nor (_18263_, _05415_, _03115_);
  or (_18264_, _18263_, _18262_);
  nand (_18265_, _18264_, _07623_);
  and (_18266_, _05417_, _01690_);
  nor (_18267_, _18266_, _02164_);
  and (_18268_, _18267_, _18265_);
  or (_18269_, _18268_, _17879_);
  nand (_18270_, _18269_, _05430_);
  and (_18271_, _05426_, _03115_);
  nor (_18272_, _18271_, _06467_);
  nand (_18273_, _18272_, _18270_);
  and (_18274_, _06467_, _02676_);
  nor (_18275_, _18274_, _02025_);
  and (_18276_, _18275_, _18273_);
  or (_18277_, _18276_, _17878_);
  nand (_18278_, _18277_, _08714_);
  nor (_18279_, _05441_, _08517_);
  not (_18280_, _18279_);
  nor (_18282_, _08714_, _01690_);
  nor (_18283_, _18282_, _18280_);
  nand (_18284_, _18283_, _18278_);
  nor (_18285_, _18279_, _03115_);
  nor (_18286_, _18285_, _01594_);
  and (_18287_, _18286_, _18284_);
  or (_18288_, _18287_, _17871_);
  nand (_18289_, _18288_, _05457_);
  and (_18290_, _05453_, _03115_);
  nor (_18291_, _18290_, _17605_);
  nand (_18293_, _18291_, _18289_);
  and (_18294_, _17605_, _02676_);
  nor (_18295_, _18294_, _05464_);
  nand (_18296_, _18295_, _18293_);
  nand (_18297_, _18296_, _17870_);
  or (_18298_, _18297_, _26506_);
  or (_18299_, _26505_, \oc8051_golden_model_1.PC [1]);
  and (_18300_, _18299_, _25964_);
  and (_27915_, _18300_, _18298_);
  and (_18301_, _01770_, _01594_);
  and (_18303_, _02164_, _01770_);
  nor (_18304_, _02818_, _01724_);
  nor (_18305_, _03564_, _02718_);
  nor (_18306_, _05139_, _01724_);
  and (_18307_, _05097_, _02057_);
  nor (_18308_, _02830_, _01724_);
  and (_18309_, _01924_, _01792_);
  nor (_18310_, _04928_, _01724_);
  nor (_18311_, _04897_, _01770_);
  and (_18312_, _02880_, _02057_);
  and (_18314_, _04874_, _03112_);
  and (_18315_, _03124_, _03121_);
  nor (_18316_, _18315_, _03125_);
  not (_18317_, _18316_);
  nor (_18318_, _18317_, _04874_);
  nor (_18319_, _18318_, _18314_);
  or (_18320_, _18319_, _02378_);
  and (_18321_, _04085_, _03112_);
  nor (_18322_, _18317_, _04085_);
  or (_18323_, _18322_, _18321_);
  nor (_18325_, _18323_, _04090_);
  and (_18326_, _01967_, _01770_);
  and (_18327_, _04710_, _01770_);
  and (_18328_, _04655_, _04652_);
  nor (_18329_, _18328_, _04656_);
  and (_18330_, _18329_, _04707_);
  or (_18331_, _18330_, _18327_);
  nor (_18332_, _18331_, _04709_);
  and (_18333_, _02309_, _04568_);
  not (_18334_, _04563_);
  and (_18336_, _04561_, _18334_);
  nor (_18337_, _18336_, _01724_);
  not (_18338_, _18337_);
  and (_18339_, _04571_, _01792_);
  not (_18340_, _04560_);
  nor (_18341_, _04571_, \oc8051_golden_model_1.PC [2]);
  and (_18342_, _18341_, _18340_);
  nor (_18343_, _18342_, _18339_);
  nor (_18344_, _04563_, _04568_);
  and (_18345_, _18344_, _17901_);
  not (_18347_, _18345_);
  nor (_18348_, _18347_, _18343_);
  nor (_18349_, _18348_, _01971_);
  and (_18350_, _18349_, _18338_);
  not (_18351_, _18350_);
  nor (_18352_, _18351_, _18333_);
  and (_18353_, _01971_, _01770_);
  or (_18354_, _18353_, _18352_);
  and (_18355_, _18354_, _17894_);
  and (_18356_, _04562_, _01724_);
  or (_18358_, _18356_, _18355_);
  and (_18359_, _18358_, _01627_);
  nor (_18360_, _02309_, _01627_);
  nor (_18361_, _18360_, _04557_);
  not (_18362_, _18361_);
  nor (_18363_, _18362_, _18359_);
  or (_18364_, _18363_, _04715_);
  nor (_18365_, _18364_, _18332_);
  and (_18366_, _04715_, _01724_);
  or (_18367_, _18366_, _01969_);
  or (_18369_, _18367_, _18365_);
  and (_18370_, _04553_, _03112_);
  and (_18371_, _18316_, _04551_);
  or (_18372_, _18371_, _02438_);
  or (_18373_, _18372_, _18370_);
  and (_18374_, _18373_, _18369_);
  nor (_18375_, _18374_, _04094_);
  and (_18376_, _04094_, _02057_);
  nor (_18377_, _18376_, _01959_);
  not (_18378_, _18377_);
  nor (_18380_, _18378_, _18375_);
  and (_18381_, _01959_, _01770_);
  or (_18382_, _18381_, _18380_);
  and (_18383_, _18382_, _01621_);
  nor (_18384_, _02309_, _01621_);
  or (_18385_, _18384_, _18383_);
  and (_18386_, _18385_, _05487_);
  or (_18387_, _18386_, _04725_);
  or (_18388_, _18387_, _18326_);
  and (_18389_, _04725_, _02057_);
  nor (_18391_, _18389_, _01963_);
  nand (_18392_, _18391_, _18388_);
  and (_18393_, _01963_, _01770_);
  nor (_18394_, _18393_, _04734_);
  nand (_18395_, _18394_, _18392_);
  and (_18396_, _04734_, _02057_);
  nor (_18397_, _18396_, _01957_);
  nand (_18398_, _18397_, _18395_);
  and (_18399_, _01957_, _01770_);
  nor (_18400_, _18399_, _17638_);
  nand (_18402_, _18400_, _18398_);
  and (_18403_, _02309_, _17638_);
  nor (_18404_, _18403_, _01953_);
  nand (_18405_, _18404_, _18402_);
  and (_18406_, _01953_, _01770_);
  nor (_18407_, _18406_, _04089_);
  and (_18408_, _18407_, _18405_);
  or (_18409_, _18408_, _18325_);
  and (_18410_, _18409_, _03187_);
  and (_18411_, _03909_, _03112_);
  nor (_18413_, _18317_, _03909_);
  or (_18414_, _18413_, _03187_);
  nor (_18415_, _18414_, _18411_);
  or (_18416_, _18415_, _18410_);
  or (_18417_, _18416_, _01951_);
  and (_18418_, _18417_, _18320_);
  or (_18419_, _18418_, _03179_);
  and (_18420_, _03113_, _02912_);
  nor (_18421_, _18316_, _02912_);
  or (_18422_, _18421_, _04749_);
  nor (_18424_, _18422_, _18420_);
  nor (_18425_, _18424_, _02880_);
  and (_18426_, _18425_, _18419_);
  or (_18427_, _18426_, _18312_);
  nand (_18428_, _18427_, _04885_);
  and (_18429_, _01946_, _01792_);
  nor (_18430_, _18429_, _06393_);
  nand (_18431_, _18430_, _18428_);
  nor (_18432_, _02309_, _01632_);
  nor (_18433_, _18432_, _18009_);
  and (_18435_, _18433_, _18431_);
  or (_18436_, _18435_, _18311_);
  nand (_18437_, _18436_, _04905_);
  nor (_18438_, _04905_, _01724_);
  nor (_18439_, _18438_, _01931_);
  nand (_18440_, _18439_, _18437_);
  and (_18441_, _01931_, _01770_);
  nor (_18442_, _18441_, _17710_);
  nand (_18443_, _18442_, _18440_);
  and (_18444_, _02309_, _17710_);
  nor (_18445_, _18444_, _01930_);
  nand (_18446_, _18445_, _18443_);
  and (_18447_, _01930_, _01770_);
  nor (_18448_, _18447_, _04933_);
  and (_18449_, _18448_, _18446_);
  or (_18450_, _18449_, _18310_);
  nand (_18451_, _18450_, _04937_);
  and (_18452_, _04932_, _01792_);
  nor (_18453_, _18452_, _01611_);
  nand (_18454_, _18453_, _18451_);
  and (_18456_, _01724_, _01611_);
  nor (_18457_, _18456_, _01924_);
  and (_18458_, _18457_, _18454_);
  or (_18459_, _18458_, _18309_);
  nand (_18460_, _18459_, _07270_);
  and (_18461_, _02309_, _01606_);
  nor (_18462_, _18461_, _02001_);
  nand (_18463_, _18462_, _18460_);
  and (_18464_, _03112_, _02001_);
  nor (_18465_, _18464_, _04953_);
  nand (_18467_, _18465_, _18463_);
  nor (_18468_, _04952_, _01770_);
  nor (_18469_, _18468_, _01602_);
  and (_18470_, _18469_, _18467_);
  and (_18471_, _03112_, _01602_);
  or (_18472_, _18471_, _04960_);
  or (_18473_, _18472_, _18470_);
  and (_18474_, _04960_, _02057_);
  nor (_18475_, _18474_, _01920_);
  and (_18476_, _18475_, _18473_);
  and (_18478_, _01920_, _01770_);
  or (_18479_, _18478_, _01654_);
  nor (_18480_, _18479_, _18476_);
  and (_18481_, _02309_, _01654_);
  or (_18482_, _18481_, _18480_);
  nand (_18483_, _18482_, _04969_);
  and (_18484_, _02032_, _01649_);
  nor (_18485_, _18329_, _04969_);
  nor (_18486_, _18485_, _18484_);
  nand (_18487_, _18486_, _18483_);
  and (_18489_, _18484_, _01770_);
  nor (_18490_, _02416_, _02035_);
  and (_18491_, _18490_, _02807_);
  nor (_18492_, _18491_, _02856_);
  nor (_18493_, _18492_, _18489_);
  nand (_18494_, _18493_, _18487_);
  and (_18495_, _18492_, _01792_);
  and (_18496_, _07430_, _01927_);
  nor (_18497_, _18496_, _18495_);
  nand (_18498_, _18497_, _18494_);
  not (_18500_, _07049_);
  nand (_18501_, _18496_, _01770_);
  and (_18502_, _18501_, _18500_);
  nand (_18503_, _18502_, _18498_);
  and (_18504_, _07049_, _01792_);
  nor (_18505_, _18504_, _02019_);
  nand (_18506_, _18505_, _18503_);
  and (_18507_, _03112_, _02019_);
  nor (_18508_, _18507_, _02853_);
  and (_18509_, _18508_, _18506_);
  and (_18511_, _02853_, _01792_);
  or (_18512_, _18511_, _18509_);
  nand (_18513_, _18512_, _04985_);
  and (_18514_, _04984_, _01776_);
  nor (_18515_, _18514_, _01919_);
  nand (_18516_, _18515_, _18513_);
  and (_18517_, _01919_, _01770_);
  nor (_18518_, _18517_, _01650_);
  nand (_18519_, _18518_, _18516_);
  and (_18520_, _02309_, _01650_);
  nor (_18522_, _18520_, _05026_);
  nand (_18523_, _18522_, _18519_);
  nor (_18524_, _18329_, _05038_);
  and (_18525_, _05038_, _01792_);
  nor (_18526_, _18525_, _05027_);
  not (_18527_, _18526_);
  nor (_18528_, _18527_, _18524_);
  nor (_18529_, _18528_, _05031_);
  and (_18530_, _18529_, _18523_);
  or (_18531_, _18530_, _18308_);
  nand (_18533_, _18531_, _05050_);
  and (_18534_, _05047_, _01792_);
  nor (_18535_, _18534_, _02018_);
  nand (_18536_, _18535_, _18533_);
  and (_18537_, _03112_, _02018_);
  nor (_18538_, _18537_, _02135_);
  and (_18539_, _18538_, _18536_);
  and (_18540_, _02135_, _01792_);
  or (_18541_, _18540_, _18539_);
  nand (_18542_, _18541_, _17617_);
  and (_18544_, _02309_, _01653_);
  nor (_18545_, _18544_, _05059_);
  nand (_18546_, _18545_, _18542_);
  nor (_18547_, _05038_, _01792_);
  and (_18548_, _18329_, _05038_);
  or (_18549_, _18548_, _18547_);
  and (_18550_, _18549_, _05059_);
  nor (_18551_, _18550_, _05069_);
  nand (_18552_, _18551_, _18546_);
  and (_18553_, _05069_, _02057_);
  nor (_18555_, _18553_, _05072_);
  and (_18556_, _18555_, _18552_);
  and (_18557_, _05072_, _01770_);
  or (_18558_, _18557_, _02039_);
  or (_18559_, _18558_, _18556_);
  and (_18560_, _03113_, _02039_);
  nor (_18561_, _18560_, _02130_);
  nand (_18562_, _18561_, _18559_);
  and (_18563_, _02130_, _01770_);
  nor (_18564_, _18563_, _01666_);
  nand (_18566_, _18564_, _18562_);
  and (_18567_, _02309_, _01666_);
  nor (_18568_, _18567_, _05086_);
  nand (_18569_, _18568_, _18566_);
  nor (_18570_, _18329_, \oc8051_golden_model_1.PSW [7]);
  nor (_18571_, _01770_, _05092_);
  nor (_18572_, _18571_, _05087_);
  not (_18573_, _18572_);
  nor (_18574_, _18573_, _18570_);
  nor (_18575_, _18574_, _05097_);
  and (_18577_, _18575_, _18569_);
  or (_18578_, _18577_, _18307_);
  nand (_18579_, _18578_, _05105_);
  and (_18580_, _05101_, _01792_);
  nor (_18581_, _18580_, _02016_);
  and (_18582_, _18581_, _18579_);
  and (_18583_, _03112_, _02016_);
  or (_18584_, _18583_, _02126_);
  nor (_18585_, _18584_, _18582_);
  and (_18586_, _02126_, _01792_);
  or (_18588_, _18586_, _18585_);
  nand (_18589_, _18588_, _17611_);
  and (_18590_, _02309_, _01663_);
  nor (_18591_, _18590_, _05114_);
  nand (_18592_, _18591_, _18589_);
  nor (_18593_, _18329_, _05092_);
  nor (_18594_, _01770_, \oc8051_golden_model_1.PSW [7]);
  nor (_18595_, _18594_, _05115_);
  not (_18596_, _18595_);
  nor (_18597_, _18596_, _18593_);
  nor (_18599_, _18597_, _05141_);
  and (_18600_, _18599_, _18592_);
  or (_18601_, _18600_, _18306_);
  nand (_18602_, _18601_, _05147_);
  and (_18603_, _02273_, _01792_);
  nor (_18604_, _18603_, _05145_);
  nand (_18605_, _18604_, _18602_);
  and (_18606_, _05145_, _01724_);
  nor (_18607_, _18606_, _02146_);
  and (_18608_, _18607_, _18605_);
  or (_18610_, _18608_, _18305_);
  nand (_18611_, _18610_, _05157_);
  and (_18612_, _02309_, _01660_);
  nor (_18613_, _18612_, _02015_);
  nand (_18614_, _18613_, _18611_);
  nor (_18615_, _05386_, _03112_);
  and (_18616_, _18317_, _05386_);
  or (_18617_, _18616_, _02153_);
  nor (_18618_, _18617_, _18615_);
  nor (_18619_, _18618_, _05161_);
  and (_18621_, _18619_, _18614_);
  or (_18622_, _18621_, _18304_);
  nand (_18623_, _18622_, _05398_);
  and (_18624_, _01792_, _02788_);
  nor (_18625_, _18624_, _05396_);
  nand (_18626_, _18625_, _18623_);
  and (_18627_, _05396_, _01724_);
  nor (_18628_, _18627_, _01585_);
  and (_18629_, _18628_, _18626_);
  nor (_18630_, _03564_, _01596_);
  or (_18632_, _18630_, _18629_);
  nand (_18633_, _18632_, _05407_);
  and (_18634_, _02309_, _01581_);
  nor (_18635_, _18634_, _02022_);
  nand (_18636_, _18635_, _18633_);
  nor (_18637_, _18316_, _05386_);
  and (_18638_, _05386_, _03113_);
  nor (_18639_, _18638_, _18637_);
  and (_18640_, _18639_, _02022_);
  nor (_18641_, _18640_, _05419_);
  nand (_18643_, _18641_, _18636_);
  nor (_18644_, _05418_, _01724_);
  nor (_18645_, _18644_, _02164_);
  and (_18646_, _18645_, _18643_);
  or (_18647_, _18646_, _18303_);
  nand (_18648_, _18647_, _05430_);
  and (_18649_, _05426_, _01724_);
  nor (_18650_, _18649_, _06467_);
  nand (_18651_, _18650_, _18648_);
  and (_18652_, _06467_, _02309_);
  nor (_18654_, _18652_, _02025_);
  nand (_18655_, _18654_, _18651_);
  and (_18656_, _18639_, _02025_);
  nor (_18657_, _18656_, _05446_);
  nand (_18658_, _18657_, _18655_);
  nor (_18659_, _05445_, _01724_);
  nor (_18660_, _18659_, _01594_);
  and (_18661_, _18660_, _18658_);
  or (_18662_, _18661_, _18301_);
  nand (_18663_, _18662_, _05457_);
  and (_18665_, _05453_, _01724_);
  nor (_18666_, _18665_, _17605_);
  nand (_18667_, _18666_, _18663_);
  and (_18668_, _17605_, _02309_);
  nor (_18669_, _18668_, _05464_);
  nand (_18670_, _18669_, _18667_);
  and (_18671_, _01724_, _05464_);
  not (_18672_, _18671_);
  and (_18673_, _18672_, _18670_);
  nand (_18674_, _18673_, _26505_);
  or (_18676_, _26505_, \oc8051_golden_model_1.PC [2]);
  and (_18677_, _18676_, _25964_);
  and (_27916_, _18677_, _18674_);
  and (_18678_, _05464_, _01760_);
  and (_18679_, _01720_, _01594_);
  and (_18680_, _05426_, _01735_);
  nor (_18681_, _02818_, _01760_);
  nor (_18682_, _03516_, _02718_);
  nor (_18683_, _05139_, _01760_);
  and (_18684_, _05097_, _01735_);
  and (_18686_, _05069_, _01735_);
  nor (_18687_, _02830_, _01760_);
  and (_18688_, _01924_, _02060_);
  nor (_18689_, _04928_, _01760_);
  nor (_18690_, _02119_, _01632_);
  and (_18691_, _02880_, _01735_);
  or (_18692_, _03110_, _03109_);
  and (_18693_, _18692_, _03126_);
  nor (_18694_, _18692_, _03126_);
  nor (_18695_, _18694_, _18693_);
  not (_18697_, _18695_);
  nor (_18698_, _18697_, _04874_);
  and (_18699_, _04874_, _03107_);
  nor (_18700_, _18699_, _18698_);
  or (_18701_, _18700_, _02378_);
  and (_18702_, _04085_, _03107_);
  nor (_18703_, _18697_, _04085_);
  or (_18704_, _18703_, _18702_);
  nor (_18705_, _18704_, _04090_);
  and (_18706_, _01967_, _01720_);
  and (_18708_, _04553_, _03107_);
  and (_18709_, _18695_, _04551_);
  or (_18710_, _18709_, _02438_);
  or (_18711_, _18710_, _18708_);
  and (_18712_, _04710_, _01720_);
  or (_18713_, _04645_, _04644_);
  and (_18714_, _18713_, _04657_);
  nor (_18715_, _18713_, _04657_);
  nor (_18716_, _18715_, _18714_);
  and (_18717_, _18716_, _04707_);
  or (_18719_, _18717_, _18712_);
  nor (_18720_, _18719_, _04709_);
  nor (_18721_, _02119_, _01625_);
  and (_18722_, _04571_, _02060_);
  nor (_18723_, _18722_, _04559_);
  nor (_18724_, _04560_, _01294_);
  or (_18725_, _18724_, _04571_);
  and (_18726_, _18725_, _18723_);
  nor (_18727_, _04561_, _01735_);
  or (_18728_, _18727_, _04563_);
  or (_18730_, _18728_, _18726_);
  and (_18731_, _18730_, _01625_);
  nor (_18732_, _18731_, _18721_);
  and (_18733_, _04563_, _01735_);
  nor (_18734_, _18733_, _01971_);
  not (_18735_, _18734_);
  nor (_18736_, _18735_, _18732_);
  and (_18737_, _01971_, _01720_);
  or (_18738_, _18737_, _18736_);
  and (_18739_, _18738_, _17894_);
  and (_18741_, _04562_, _01760_);
  or (_18742_, _18741_, _18739_);
  and (_18743_, _18742_, _01627_);
  nor (_18744_, _02119_, _01627_);
  nor (_18745_, _18744_, _04557_);
  not (_18746_, _18745_);
  nor (_18747_, _18746_, _18743_);
  or (_18748_, _18747_, _04715_);
  nor (_18749_, _18748_, _18720_);
  and (_18750_, _04715_, _01760_);
  or (_18752_, _18750_, _01969_);
  or (_18753_, _18752_, _18749_);
  and (_18754_, _18753_, _18711_);
  nor (_18755_, _18754_, _04094_);
  and (_18756_, _04094_, _01735_);
  nor (_18757_, _18756_, _01959_);
  not (_18758_, _18757_);
  nor (_18759_, _18758_, _18755_);
  and (_18760_, _01959_, _01720_);
  or (_18761_, _18760_, _18759_);
  and (_18763_, _18761_, _01621_);
  nor (_18764_, _02119_, _01621_);
  or (_18765_, _18764_, _18763_);
  and (_18766_, _18765_, _05487_);
  or (_18767_, _18766_, _04725_);
  or (_18768_, _18767_, _18706_);
  and (_18769_, _04725_, _01735_);
  nor (_18770_, _18769_, _01963_);
  nand (_18771_, _18770_, _18768_);
  and (_18772_, _01963_, _01720_);
  nor (_18774_, _18772_, _04734_);
  nand (_18775_, _18774_, _18771_);
  and (_18776_, _04734_, _01735_);
  nor (_18777_, _18776_, _01957_);
  nand (_18778_, _18777_, _18775_);
  and (_18779_, _01957_, _01720_);
  nor (_18780_, _18779_, _17638_);
  nand (_18781_, _18780_, _18778_);
  and (_18782_, _02119_, _17638_);
  nor (_18783_, _18782_, _01953_);
  nand (_18785_, _18783_, _18781_);
  and (_18786_, _01953_, _01720_);
  nor (_18787_, _18786_, _04089_);
  and (_18788_, _18787_, _18785_);
  or (_18789_, _18788_, _18705_);
  and (_18790_, _18789_, _03187_);
  and (_18791_, _03909_, _03107_);
  nor (_18792_, _18697_, _03909_);
  or (_18793_, _18792_, _18791_);
  nor (_18794_, _18793_, _03187_);
  or (_18796_, _18794_, _18790_);
  or (_18797_, _18796_, _01951_);
  and (_18798_, _18797_, _18701_);
  or (_18799_, _18798_, _03179_);
  nor (_18800_, _18695_, _02912_);
  and (_18801_, _03108_, _02912_);
  or (_18802_, _18801_, _04749_);
  or (_18803_, _18802_, _18800_);
  and (_18804_, _18803_, _02881_);
  and (_18805_, _18804_, _18799_);
  or (_18807_, _18805_, _18691_);
  nand (_18808_, _18807_, _04885_);
  and (_18809_, _01946_, _02060_);
  nor (_18810_, _18809_, _06393_);
  nand (_18811_, _18810_, _18808_);
  nand (_18812_, _18811_, _04897_);
  nor (_18813_, _18812_, _18690_);
  nor (_18814_, _04897_, _01720_);
  or (_18815_, _18814_, _18813_);
  nand (_18816_, _18815_, _04905_);
  nor (_18818_, _04905_, _01760_);
  nor (_18819_, _18818_, _01931_);
  nand (_18820_, _18819_, _18816_);
  and (_18821_, _01931_, _01720_);
  nor (_18822_, _18821_, _17710_);
  nand (_18823_, _18822_, _18820_);
  and (_18824_, _02119_, _17710_);
  nor (_18825_, _18824_, _01930_);
  nand (_18826_, _18825_, _18823_);
  and (_18827_, _01930_, _01720_);
  nor (_18829_, _18827_, _04933_);
  and (_18830_, _18829_, _18826_);
  or (_18831_, _18830_, _18689_);
  nand (_18832_, _18831_, _04937_);
  and (_18833_, _04932_, _02060_);
  nor (_18834_, _18833_, _01611_);
  nand (_18835_, _18834_, _18832_);
  and (_18836_, _01611_, _01760_);
  nor (_18837_, _18836_, _01924_);
  and (_18838_, _18837_, _18835_);
  or (_18840_, _18838_, _18688_);
  nand (_18841_, _18840_, _07270_);
  and (_18842_, _02119_, _01606_);
  nor (_18843_, _18842_, _02001_);
  nand (_18844_, _18843_, _18841_);
  and (_18845_, _03107_, _02001_);
  nor (_18846_, _18845_, _04953_);
  nand (_18847_, _18846_, _18844_);
  nor (_18848_, _04952_, _01720_);
  nor (_18849_, _18848_, _01602_);
  and (_18851_, _18849_, _18847_);
  nor (_18852_, _04960_, _03107_);
  nor (_18853_, _18852_, _17728_);
  or (_18854_, _18853_, _18851_);
  and (_18855_, _04960_, _01735_);
  nor (_18856_, _18855_, _01920_);
  nand (_18857_, _18856_, _18854_);
  and (_18858_, _01920_, _01720_);
  nor (_18859_, _18858_, _01654_);
  nand (_18860_, _18859_, _18857_);
  and (_18862_, _02119_, _01654_);
  nor (_18863_, _18862_, _04968_);
  nand (_18864_, _18863_, _18860_);
  and (_18865_, _18716_, _04968_);
  nor (_18866_, _18865_, _02859_);
  nand (_18867_, _18866_, _18864_);
  and (_18868_, _02859_, _02060_);
  nor (_18869_, _18868_, _02019_);
  nand (_18870_, _18869_, _18867_);
  and (_18871_, _03107_, _02019_);
  nor (_18873_, _18871_, _02853_);
  and (_18874_, _18873_, _18870_);
  and (_18875_, _02853_, _02060_);
  or (_18876_, _18875_, _18874_);
  nand (_18877_, _18876_, _04985_);
  nor (_18878_, _04985_, _01757_);
  nor (_18879_, _18878_, _01919_);
  nand (_18880_, _18879_, _18877_);
  and (_18881_, _01919_, _01720_);
  nor (_18882_, _18881_, _01650_);
  nand (_18884_, _18882_, _18880_);
  and (_18885_, _02119_, _01650_);
  nor (_18886_, _18885_, _05026_);
  nand (_18887_, _18886_, _18884_);
  and (_18888_, _05038_, _01720_);
  and (_18889_, _18716_, _05040_);
  or (_18890_, _18889_, _18888_);
  and (_18891_, _18890_, _05026_);
  nor (_18892_, _18891_, _05031_);
  and (_18893_, _18892_, _18887_);
  or (_18895_, _18893_, _18687_);
  nand (_18896_, _18895_, _05050_);
  and (_18897_, _05047_, _02060_);
  nor (_18898_, _18897_, _02018_);
  and (_18899_, _18898_, _18896_);
  and (_18900_, _03107_, _02018_);
  or (_18901_, _18900_, _02135_);
  nor (_18902_, _18901_, _18899_);
  and (_18903_, _02135_, _02060_);
  or (_18904_, _18903_, _18902_);
  nand (_18906_, _18904_, _17617_);
  and (_18907_, _02119_, _01653_);
  nor (_18908_, _18907_, _05059_);
  nand (_18909_, _18908_, _18906_);
  and (_18910_, _05040_, _01720_);
  and (_18911_, _18716_, _05038_);
  or (_18912_, _18911_, _18910_);
  and (_18913_, _18912_, _05059_);
  nor (_18914_, _18913_, _05069_);
  and (_18915_, _18914_, _18909_);
  or (_18917_, _18915_, _18686_);
  nand (_18918_, _18917_, _05077_);
  and (_18919_, _05072_, _02060_);
  nor (_18920_, _18919_, _02039_);
  and (_18921_, _18920_, _18918_);
  and (_18922_, _03107_, _02039_);
  or (_18923_, _18922_, _02130_);
  nor (_18924_, _18923_, _18921_);
  and (_18925_, _02130_, _02060_);
  or (_18926_, _18925_, _18924_);
  nand (_18928_, _18926_, _17614_);
  and (_18929_, _02119_, _01666_);
  nor (_18930_, _18929_, _05086_);
  nand (_18931_, _18930_, _18928_);
  nor (_18932_, _18716_, \oc8051_golden_model_1.PSW [7]);
  nor (_18933_, _01720_, _05092_);
  nor (_18934_, _18933_, _05087_);
  not (_18935_, _18934_);
  nor (_18936_, _18935_, _18932_);
  nor (_18937_, _18936_, _05097_);
  and (_18939_, _18937_, _18931_);
  or (_18940_, _18939_, _18684_);
  nand (_18941_, _18940_, _05105_);
  and (_18942_, _05101_, _02060_);
  nor (_18943_, _18942_, _02016_);
  and (_18944_, _18943_, _18941_);
  and (_18945_, _03107_, _02016_);
  or (_18946_, _18945_, _02126_);
  nor (_18947_, _18946_, _18944_);
  and (_18948_, _02126_, _02060_);
  or (_18950_, _18948_, _18947_);
  nand (_18951_, _18950_, _17611_);
  and (_18952_, _02119_, _01663_);
  nor (_18953_, _18952_, _05114_);
  nand (_18954_, _18953_, _18951_);
  nor (_18955_, _18716_, _05092_);
  nor (_18956_, _01720_, \oc8051_golden_model_1.PSW [7]);
  nor (_18957_, _18956_, _05115_);
  not (_18958_, _18957_);
  nor (_18959_, _18958_, _18955_);
  nor (_18961_, _18959_, _05141_);
  and (_18962_, _18961_, _18954_);
  or (_18963_, _18962_, _18683_);
  nand (_18964_, _18963_, _05147_);
  and (_18965_, _02273_, _02060_);
  nor (_18966_, _18965_, _05145_);
  nand (_18967_, _18966_, _18964_);
  and (_18968_, _05145_, _01760_);
  nor (_18969_, _18968_, _02146_);
  and (_18970_, _18969_, _18967_);
  or (_18972_, _18970_, _18682_);
  nand (_18973_, _18972_, _05157_);
  and (_18974_, _02119_, _01660_);
  nor (_18975_, _18974_, _02015_);
  nand (_18976_, _18975_, _18973_);
  and (_18977_, _18697_, _05386_);
  nor (_18978_, _05386_, _03107_);
  or (_18979_, _18978_, _02153_);
  nor (_18980_, _18979_, _18977_);
  nor (_18981_, _18980_, _05161_);
  and (_18982_, _18981_, _18976_);
  or (_18983_, _18982_, _18681_);
  nand (_18984_, _18983_, _05398_);
  and (_18985_, _02060_, _02788_);
  nor (_18986_, _18985_, _05396_);
  nand (_18987_, _18986_, _18984_);
  and (_18988_, _05396_, _01760_);
  nor (_18989_, _18988_, _01585_);
  and (_18990_, _18989_, _18987_);
  nor (_18991_, _03516_, _01596_);
  or (_18994_, _18991_, _18990_);
  nand (_18995_, _18994_, _05407_);
  and (_18996_, _02119_, _01581_);
  nor (_18997_, _18996_, _02022_);
  nand (_18998_, _18997_, _18995_);
  and (_18999_, _05386_, _03108_);
  nor (_19000_, _18695_, _05386_);
  nor (_19001_, _19000_, _18999_);
  and (_19002_, _19001_, _02022_);
  nor (_19003_, _19002_, _05419_);
  nand (_19005_, _19003_, _18998_);
  nor (_19006_, _05418_, _01760_);
  nor (_19007_, _19006_, _02164_);
  nand (_19008_, _19007_, _19005_);
  and (_19009_, _02164_, _01720_);
  nor (_19010_, _19009_, _05426_);
  and (_19011_, _19010_, _19008_);
  or (_19012_, _19011_, _18680_);
  nand (_19013_, _19012_, _06466_);
  and (_19014_, _06467_, _02119_);
  nor (_19016_, _19014_, _02025_);
  nand (_19017_, _19016_, _19013_);
  and (_19018_, _19001_, _02025_);
  nor (_19019_, _19018_, _05446_);
  nand (_19020_, _19019_, _19017_);
  nor (_19021_, _05445_, _01760_);
  nor (_19022_, _19021_, _01594_);
  and (_19023_, _19022_, _19020_);
  or (_19024_, _19023_, _18679_);
  nand (_19025_, _19024_, _05457_);
  and (_19027_, _05453_, _01760_);
  nor (_19028_, _19027_, _17605_);
  nand (_19029_, _19028_, _19025_);
  and (_19030_, _17605_, _02119_);
  nor (_19031_, _19030_, _05464_);
  and (_19032_, _19031_, _19029_);
  or (_19033_, _19032_, _18678_);
  or (_19034_, _19033_, _26506_);
  or (_19035_, _26505_, \oc8051_golden_model_1.PC [3]);
  and (_19036_, _19035_, _25964_);
  and (_27917_, _19036_, _19034_);
  not (_19038_, \oc8051_golden_model_1.PC [4]);
  nor (_19039_, _01312_, _19038_);
  and (_19040_, _01312_, _19038_);
  nor (_19041_, _19040_, _19039_);
  and (_19042_, _19041_, _05464_);
  not (_19043_, _19042_);
  and (_19044_, _06467_, _03101_);
  and (_19045_, _04641_, _05092_);
  and (_19046_, _04662_, _04659_);
  nor (_19048_, _19046_, _04663_);
  and (_19049_, _19048_, \oc8051_golden_model_1.PSW [7]);
  or (_19050_, _19049_, _19045_);
  and (_19051_, _19050_, _05114_);
  and (_19052_, _05038_, _04641_);
  and (_19053_, _19048_, _05040_);
  or (_19054_, _19053_, _19052_);
  and (_19055_, _19054_, _05026_);
  and (_19056_, _04642_, _01924_);
  and (_19057_, _04874_, _03103_);
  and (_19059_, _03131_, _03128_);
  nor (_19060_, _19059_, _03132_);
  not (_19061_, _19060_);
  nor (_19062_, _19061_, _04874_);
  nor (_19063_, _19062_, _19057_);
  nor (_19064_, _19063_, _02378_);
  and (_19065_, _03909_, _03103_);
  nor (_19066_, _19061_, _03909_);
  or (_19067_, _19066_, _19065_);
  and (_19068_, _19067_, _03185_);
  and (_19070_, _04641_, _01959_);
  or (_19071_, _04551_, _03104_);
  or (_19072_, _19061_, _04553_);
  and (_19073_, _19072_, _01969_);
  and (_19074_, _19073_, _19071_);
  and (_19075_, _04710_, _04641_);
  and (_19076_, _19048_, _04707_);
  nor (_19077_, _19076_, _19075_);
  nand (_19078_, _19077_, _04557_);
  and (_19079_, _04642_, _01971_);
  and (_19081_, _03101_, _04568_);
  nor (_19082_, _04560_, \oc8051_golden_model_1.PC [4]);
  or (_19083_, _19082_, _04571_);
  and (_19084_, _04571_, _04641_);
  nor (_19085_, _19084_, _04559_);
  and (_19086_, _19085_, _19083_);
  nor (_19087_, _19041_, _04561_);
  or (_19088_, _19087_, _04563_);
  or (_19089_, _19088_, _19086_);
  and (_19090_, _19089_, _01625_);
  nor (_19092_, _19090_, _19081_);
  and (_19093_, _19041_, _04563_);
  nor (_19094_, _19093_, _01971_);
  not (_19095_, _19094_);
  nor (_19096_, _19095_, _19092_);
  nor (_19097_, _19096_, _19079_);
  and (_19098_, _19097_, _17894_);
  and (_19099_, _19041_, _04562_);
  or (_19100_, _19099_, _19098_);
  and (_19101_, _19100_, _01627_);
  nor (_19103_, _03101_, _01627_);
  nor (_19104_, _19103_, _04557_);
  not (_19105_, _19104_);
  nor (_19106_, _19105_, _19101_);
  nor (_19107_, _19106_, _04715_);
  nand (_19108_, _19107_, _19078_);
  and (_19109_, _19041_, _04715_);
  nor (_19110_, _19109_, _01969_);
  and (_19111_, _19110_, _19108_);
  or (_19112_, _19111_, _19074_);
  nand (_19114_, _19112_, _17940_);
  not (_19115_, _19041_);
  and (_19116_, _19115_, _04094_);
  nor (_19117_, _19116_, _01959_);
  and (_19118_, _19117_, _19114_);
  or (_19119_, _19118_, _19070_);
  and (_19120_, _19119_, _01621_);
  nor (_19121_, _03101_, _01621_);
  or (_19122_, _19121_, _01967_);
  or (_19123_, _19122_, _19120_);
  and (_19125_, _04642_, _01967_);
  nor (_19126_, _19125_, _04725_);
  nand (_19127_, _19126_, _19123_);
  and (_19128_, _19041_, _04725_);
  nor (_19129_, _19128_, _01963_);
  nand (_19130_, _19129_, _19127_);
  and (_19131_, _04642_, _01963_);
  nor (_19132_, _19131_, _04734_);
  and (_19133_, _19132_, _19130_);
  and (_19134_, _19041_, _04734_);
  or (_19136_, _19134_, _01957_);
  or (_19137_, _19136_, _19133_);
  and (_19138_, _04642_, _01957_);
  nor (_19139_, _19138_, _17638_);
  and (_19140_, _19139_, _19137_);
  nor (_19141_, _03101_, _01630_);
  or (_19142_, _19141_, _19140_);
  nand (_19143_, _19142_, _02457_);
  and (_19144_, _04641_, _01953_);
  nor (_19145_, _19144_, _04089_);
  nand (_19147_, _19145_, _19143_);
  and (_19148_, _04085_, _03103_);
  nor (_19149_, _19061_, _04085_);
  or (_19150_, _19149_, _19148_);
  nor (_19151_, _19150_, _04090_);
  nor (_19152_, _19151_, _03185_);
  and (_19153_, _19152_, _19147_);
  nor (_19154_, _19153_, _19068_);
  nor (_19155_, _19154_, _01951_);
  or (_19156_, _19155_, _19064_);
  nand (_19158_, _19156_, _04749_);
  nand (_19159_, _03103_, _02912_);
  not (_19160_, _02912_);
  nand (_19161_, _19060_, _19160_);
  and (_19162_, _19161_, _19159_);
  or (_19163_, _19162_, _04749_);
  and (_19164_, _19163_, _19158_);
  or (_19165_, _19164_, _02880_);
  nand (_19166_, _19041_, _02880_);
  and (_19167_, _19166_, _19165_);
  nand (_19169_, _19167_, _04885_);
  and (_19170_, _04642_, _01946_);
  nor (_19171_, _19170_, _06393_);
  nand (_19172_, _19171_, _19169_);
  nor (_19173_, _03101_, _01632_);
  nor (_19174_, _19173_, _18009_);
  nand (_19175_, _19174_, _19172_);
  nor (_19176_, _04897_, _04641_);
  nor (_19177_, _19176_, _04908_);
  and (_19178_, _19177_, _19175_);
  nor (_19180_, _19115_, _04905_);
  or (_19181_, _19180_, _01931_);
  nor (_19182_, _19181_, _19178_);
  and (_19183_, _04642_, _01931_);
  or (_19184_, _19183_, _19182_);
  nand (_19185_, _19184_, _01618_);
  and (_19186_, _03101_, _17710_);
  nor (_19187_, _19186_, _01930_);
  and (_19188_, _19187_, _19185_);
  and (_19189_, _04641_, _01930_);
  or (_19191_, _19189_, _19188_);
  nand (_19192_, _19191_, _04928_);
  nor (_19193_, _19115_, _04928_);
  nor (_19194_, _19193_, _04932_);
  nand (_19195_, _19194_, _19192_);
  and (_19196_, _04642_, _04932_);
  nor (_19197_, _19196_, _01611_);
  nand (_19198_, _19197_, _19195_);
  and (_19199_, _19041_, _01611_);
  nor (_19200_, _19199_, _01924_);
  and (_19202_, _19200_, _19198_);
  or (_19203_, _19202_, _19056_);
  nand (_19204_, _19203_, _07270_);
  and (_19205_, _03101_, _01606_);
  nor (_19206_, _19205_, _02001_);
  nand (_19207_, _19206_, _19204_);
  and (_19208_, _03103_, _02001_);
  nor (_19209_, _19208_, _04953_);
  nand (_19210_, _19209_, _19207_);
  nor (_19211_, _04952_, _04641_);
  nor (_19213_, _19211_, _01602_);
  nand (_19214_, _19213_, _19210_);
  nor (_19215_, _04960_, _03103_);
  or (_19216_, _19215_, _17728_);
  and (_19217_, _19216_, _19214_);
  and (_19218_, _19115_, _04960_);
  or (_19219_, _19218_, _19217_);
  nand (_19220_, _19219_, _02519_);
  and (_19221_, _04642_, _01920_);
  nor (_19222_, _19221_, _01654_);
  and (_19224_, _19222_, _19220_);
  nor (_19225_, _03101_, _17739_);
  or (_19226_, _19225_, _19224_);
  nand (_19227_, _19226_, _04969_);
  and (_19228_, _19048_, _04968_);
  nor (_19229_, _19228_, _02859_);
  nand (_19230_, _19229_, _19227_);
  and (_19231_, _02859_, _04642_);
  nor (_19232_, _19231_, _02019_);
  nand (_19233_, _19232_, _19230_);
  and (_19235_, _03103_, _02019_);
  nor (_19236_, _19235_, _02853_);
  nand (_19237_, _19236_, _19233_);
  and (_19238_, _04642_, _02853_);
  nor (_19239_, _19238_, _04984_);
  nand (_19240_, _19239_, _19237_);
  and (_19241_, _05002_, _04999_);
  nor (_19242_, _19241_, _05003_);
  and (_19243_, _19242_, _04984_);
  nor (_19244_, _19243_, _01919_);
  and (_19246_, _19244_, _19240_);
  and (_19247_, _04642_, _01919_);
  or (_19248_, _19247_, _19246_);
  nand (_19249_, _19248_, _01651_);
  and (_19250_, _03101_, _01650_);
  nor (_19251_, _19250_, _05026_);
  and (_19252_, _19251_, _19249_);
  or (_19253_, _19252_, _19055_);
  nand (_19254_, _19253_, _02830_);
  nor (_19255_, _19115_, _02830_);
  nor (_19257_, _19255_, _05047_);
  nand (_19258_, _19257_, _19254_);
  and (_19259_, _05047_, _04642_);
  nor (_19260_, _19259_, _02018_);
  and (_19261_, _19260_, _19258_);
  and (_19262_, _03103_, _02018_);
  or (_19263_, _19262_, _02135_);
  nor (_19264_, _19263_, _19261_);
  and (_19265_, _04642_, _02135_);
  or (_19266_, _19265_, _19264_);
  nand (_19268_, _19266_, _17617_);
  and (_19269_, _03101_, _01653_);
  nor (_19270_, _19269_, _05059_);
  nand (_19271_, _19270_, _19268_);
  nand (_19272_, _05040_, _04641_);
  nand (_19273_, _19048_, _05038_);
  and (_19274_, _19273_, _19272_);
  or (_19275_, _19274_, _05060_);
  nand (_19276_, _19275_, _19271_);
  nand (_19277_, _19276_, _05070_);
  and (_19279_, _19041_, _05069_);
  nor (_19280_, _19279_, _05072_);
  nand (_19281_, _19280_, _19277_);
  and (_19282_, _04642_, _05072_);
  nor (_19283_, _19282_, _02039_);
  and (_19284_, _19283_, _19281_);
  and (_19285_, _03103_, _02039_);
  or (_19286_, _19285_, _02130_);
  nor (_19287_, _19286_, _19284_);
  and (_19288_, _04642_, _02130_);
  or (_19290_, _19288_, _19287_);
  nand (_19291_, _19290_, _17614_);
  and (_19292_, _03101_, _01666_);
  nor (_19293_, _19292_, _05086_);
  nand (_19294_, _19293_, _19291_);
  nand (_19295_, _04641_, \oc8051_golden_model_1.PSW [7]);
  nand (_19296_, _19048_, _05092_);
  and (_19297_, _19296_, _19295_);
  or (_19298_, _19297_, _05087_);
  nand (_19299_, _19298_, _19294_);
  nand (_19301_, _19299_, _05098_);
  and (_19302_, _19041_, _05097_);
  nor (_19303_, _19302_, _05101_);
  nand (_19304_, _19303_, _19301_);
  and (_19305_, _05101_, _04642_);
  nor (_19306_, _19305_, _02016_);
  nand (_19307_, _19306_, _19304_);
  and (_19308_, _03103_, _02016_);
  nor (_19309_, _19308_, _02126_);
  and (_19310_, _19309_, _19307_);
  and (_19312_, _04642_, _02126_);
  or (_19313_, _19312_, _19310_);
  nand (_19314_, _19313_, _17611_);
  and (_19315_, _03101_, _01663_);
  nor (_19316_, _19315_, _05114_);
  and (_19317_, _19316_, _19314_);
  or (_19318_, _19317_, _19051_);
  nand (_19319_, _19318_, _05139_);
  nor (_19320_, _19115_, _05139_);
  nor (_19321_, _19320_, _02273_);
  nand (_19323_, _19321_, _19319_);
  and (_19324_, _04642_, _02273_);
  nor (_19325_, _19324_, _05145_);
  nand (_19326_, _19325_, _19323_);
  and (_19327_, _19041_, _05145_);
  nor (_19328_, _19327_, _02146_);
  and (_19329_, _19328_, _19326_);
  nor (_19330_, _03903_, _02718_);
  or (_19331_, _19330_, _19329_);
  nand (_19332_, _19331_, _05157_);
  and (_19334_, _03101_, _01660_);
  nor (_19335_, _19334_, _02015_);
  and (_19336_, _19335_, _19332_);
  nor (_19337_, _05386_, _03104_);
  and (_19338_, _19060_, _05386_);
  nor (_19339_, _19338_, _19337_);
  nor (_19340_, _19339_, _02153_);
  or (_19341_, _19340_, _19336_);
  nand (_19342_, _19341_, _02818_);
  nor (_19343_, _19115_, _02818_);
  nor (_19345_, _19343_, _02788_);
  nand (_19346_, _19345_, _19342_);
  and (_19347_, _04642_, _02788_);
  nor (_19348_, _19347_, _05396_);
  nand (_19349_, _19348_, _19346_);
  and (_19350_, _19041_, _05396_);
  nor (_19351_, _19350_, _01585_);
  nand (_19352_, _19351_, _19349_);
  nor (_19353_, _03903_, _01596_);
  nor (_19354_, _19353_, _01581_);
  and (_19356_, _19354_, _19352_);
  nor (_19357_, _03101_, _05407_);
  or (_19358_, _19357_, _02022_);
  or (_19359_, _19358_, _19356_);
  and (_19360_, _05386_, _03104_);
  nor (_19361_, _19060_, _05386_);
  nor (_19362_, _19361_, _19360_);
  nor (_19363_, _19362_, _02558_);
  nor (_19364_, _19363_, _05419_);
  nand (_19365_, _19364_, _19359_);
  nor (_19367_, _19115_, _05418_);
  nor (_19368_, _19367_, _02164_);
  nand (_19369_, _19368_, _19365_);
  and (_19370_, _04642_, _02164_);
  nor (_19371_, _19370_, _05426_);
  nand (_19372_, _19371_, _19369_);
  and (_19373_, _19041_, _05426_);
  nor (_19374_, _19373_, _06467_);
  and (_19375_, _19374_, _19372_);
  or (_19376_, _19375_, _19044_);
  nand (_19378_, _19376_, _02377_);
  nor (_19379_, _19362_, _02377_);
  nor (_19380_, _19379_, _05446_);
  nand (_19381_, _19380_, _19378_);
  nor (_19382_, _19115_, _05445_);
  nor (_19383_, _19382_, _01594_);
  nand (_19384_, _19383_, _19381_);
  and (_19385_, _04642_, _01594_);
  nor (_19386_, _19385_, _05453_);
  nand (_19387_, _19386_, _19384_);
  and (_19389_, _19041_, _05453_);
  nor (_19390_, _19389_, _17605_);
  nand (_19391_, _19390_, _19387_);
  and (_19392_, _17605_, _03101_);
  nor (_19393_, _19392_, _05464_);
  nand (_19394_, _19393_, _19391_);
  and (_19395_, _19394_, _19043_);
  nand (_19396_, _19395_, _26505_);
  or (_19397_, _26505_, \oc8051_golden_model_1.PC [4]);
  and (_19398_, _19397_, _25964_);
  and (_27920_, _19398_, _19396_);
  nor (_19400_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_19401_, _04636_, _01325_);
  nor (_19402_, _19401_, _19400_);
  and (_19403_, _19402_, _05464_);
  not (_19404_, _19403_);
  and (_19405_, _04636_, _01594_);
  and (_19406_, _04636_, _02164_);
  nor (_19407_, _03850_, _01596_);
  nor (_19408_, _19402_, _02818_);
  nor (_19410_, _03850_, _02718_);
  nor (_19411_, _19402_, _05139_);
  not (_19412_, _19402_);
  and (_19413_, _19412_, _05097_);
  and (_19414_, _19412_, _05069_);
  nor (_19415_, _19402_, _02830_);
  not (_19416_, _01919_);
  and (_19417_, _04637_, _01924_);
  nor (_19418_, _19402_, _04928_);
  nor (_19419_, _04897_, _04636_);
  or (_19421_, _03070_, _03069_);
  not (_19422_, _19421_);
  nor (_19423_, _19422_, _03133_);
  and (_19424_, _19422_, _03133_);
  nor (_19425_, _19424_, _19423_);
  nor (_19426_, _19425_, _04874_);
  and (_19427_, _04874_, _03067_);
  nor (_19428_, _19427_, _19426_);
  or (_19429_, _19428_, _02378_);
  and (_19430_, _04085_, _03067_);
  nor (_19432_, _19425_, _04085_);
  or (_19433_, _19432_, _19430_);
  nor (_19434_, _19433_, _04090_);
  and (_19435_, _04553_, _03067_);
  not (_19436_, _19425_);
  and (_19437_, _19436_, _04551_);
  or (_19438_, _19437_, _02438_);
  or (_19439_, _19438_, _19435_);
  and (_19440_, _04710_, _04636_);
  or (_19441_, _04639_, _04638_);
  not (_19443_, _19441_);
  nor (_19444_, _19443_, _04664_);
  and (_19445_, _19443_, _04664_);
  nor (_19446_, _19445_, _19444_);
  nor (_19447_, _19446_, _04710_);
  or (_19448_, _19447_, _19440_);
  nor (_19449_, _19448_, _04709_);
  nor (_19450_, _03064_, _01625_);
  and (_19451_, _04571_, _04637_);
  nor (_19452_, _19451_, _04559_);
  and (_19454_, _18340_, \oc8051_golden_model_1.PC [5]);
  or (_19455_, _19454_, _04571_);
  and (_19456_, _19455_, _19452_);
  nor (_19457_, _19412_, _04561_);
  or (_19458_, _19457_, _04563_);
  or (_19459_, _19458_, _19456_);
  and (_19460_, _19459_, _01625_);
  nor (_19461_, _19460_, _19450_);
  and (_19462_, _19412_, _04563_);
  nor (_19463_, _19462_, _01971_);
  not (_19465_, _19463_);
  nor (_19466_, _19465_, _19461_);
  and (_19467_, _04636_, _01971_);
  or (_19468_, _19467_, _19466_);
  and (_19469_, _19468_, _17894_);
  and (_19470_, _19402_, _04562_);
  or (_19471_, _19470_, _19469_);
  and (_19472_, _19471_, _01627_);
  nor (_19473_, _03064_, _01627_);
  nor (_19474_, _19473_, _04557_);
  not (_19476_, _19474_);
  nor (_19477_, _19476_, _19472_);
  or (_19478_, _19477_, _04715_);
  nor (_19479_, _19478_, _19449_);
  and (_19480_, _19402_, _04715_);
  or (_19481_, _19480_, _01969_);
  or (_19482_, _19481_, _19479_);
  and (_19483_, _19482_, _19439_);
  nor (_19484_, _19483_, _04094_);
  and (_19485_, _19412_, _04094_);
  nor (_19487_, _19485_, _01959_);
  not (_19488_, _19487_);
  nor (_19489_, _19488_, _19484_);
  and (_19490_, _04636_, _01959_);
  nor (_19491_, _19490_, _19489_);
  or (_19492_, _19491_, _06363_);
  or (_19493_, _03064_, _01621_);
  and (_19494_, _19493_, _19492_);
  or (_19495_, _19494_, _01967_);
  and (_19496_, _04636_, _01967_);
  nor (_19499_, _19496_, _04725_);
  nand (_19500_, _19499_, _19495_);
  and (_19501_, _19412_, _04725_);
  nor (_19502_, _19501_, _01963_);
  nand (_19503_, _19502_, _19500_);
  and (_19504_, _04636_, _01963_);
  nor (_19505_, _19504_, _04734_);
  nand (_19506_, _19505_, _19503_);
  and (_19507_, _19412_, _04734_);
  nor (_19508_, _19507_, _01957_);
  nand (_19510_, _19508_, _19506_);
  and (_19511_, _04636_, _01957_);
  nor (_19512_, _19511_, _17638_);
  nand (_19513_, _19512_, _19510_);
  and (_19514_, _03064_, _17638_);
  nor (_19515_, _19514_, _01953_);
  nand (_19516_, _19515_, _19513_);
  and (_19517_, _04636_, _01953_);
  nor (_19518_, _19517_, _04089_);
  and (_19519_, _19518_, _19516_);
  or (_19522_, _19519_, _19434_);
  and (_19523_, _19522_, _03187_);
  and (_19524_, _03909_, _03067_);
  nor (_19525_, _19425_, _03909_);
  or (_19526_, _19525_, _19524_);
  nor (_19527_, _19526_, _03187_);
  or (_19528_, _19527_, _19523_);
  or (_19529_, _19528_, _01951_);
  and (_19530_, _19529_, _19429_);
  or (_19531_, _19530_, _03179_);
  nand (_19533_, _03067_, _02912_);
  or (_19534_, _19425_, _02912_);
  and (_19535_, _19534_, _19533_);
  or (_19536_, _19535_, _04749_);
  and (_19537_, _19536_, _19531_);
  or (_19538_, _19537_, _02880_);
  nand (_19539_, _19402_, _02880_);
  and (_19540_, _19539_, _19538_);
  nand (_19541_, _19540_, _04885_);
  and (_19542_, _04637_, _01946_);
  nor (_19545_, _19542_, _06393_);
  nand (_19546_, _19545_, _19541_);
  nor (_19547_, _03064_, _01632_);
  nor (_19548_, _19547_, _18009_);
  and (_19549_, _19548_, _19546_);
  or (_19550_, _19549_, _19419_);
  nand (_19551_, _19550_, _04905_);
  nor (_19552_, _19402_, _04905_);
  nor (_19553_, _19552_, _01931_);
  nand (_19554_, _19553_, _19551_);
  and (_19556_, _04636_, _01931_);
  nor (_19557_, _19556_, _17710_);
  nand (_19558_, _19557_, _19554_);
  and (_19559_, _03064_, _17710_);
  nor (_19560_, _19559_, _01930_);
  nand (_19561_, _19560_, _19558_);
  and (_19562_, _04636_, _01930_);
  nor (_19563_, _19562_, _04933_);
  and (_19564_, _19563_, _19561_);
  or (_19565_, _19564_, _19418_);
  nand (_19568_, _19565_, _04937_);
  and (_19569_, _04637_, _04932_);
  nor (_19570_, _19569_, _01611_);
  nand (_19571_, _19570_, _19568_);
  and (_19572_, _19402_, _01611_);
  nor (_19573_, _19572_, _01924_);
  and (_19574_, _19573_, _19571_);
  or (_19575_, _19574_, _19417_);
  nand (_19576_, _19575_, _07270_);
  and (_19577_, _03064_, _01606_);
  nor (_19579_, _19577_, _02001_);
  nand (_19580_, _19579_, _19576_);
  and (_19581_, _03067_, _02001_);
  nor (_19582_, _19581_, _04953_);
  nand (_19583_, _19582_, _19580_);
  nor (_19584_, _04952_, _04636_);
  nor (_19585_, _19584_, _01602_);
  and (_19586_, _19585_, _19583_);
  nor (_19587_, _04960_, _03067_);
  nor (_19588_, _19587_, _17728_);
  or (_19590_, _19588_, _19586_);
  and (_19591_, _19412_, _04960_);
  nor (_19592_, _19591_, _01920_);
  and (_19593_, _19592_, _19590_);
  and (_19594_, _04636_, _01920_);
  or (_19595_, _19594_, _01654_);
  or (_19596_, _19595_, _19593_);
  and (_19597_, _03064_, _01654_);
  nor (_19598_, _19597_, _04968_);
  nand (_19599_, _19598_, _19596_);
  nor (_19601_, _19446_, _04969_);
  nor (_19602_, _19601_, _02859_);
  nand (_19603_, _19602_, _19599_);
  and (_19604_, _02859_, _04637_);
  nor (_19605_, _19604_, _02019_);
  nand (_19606_, _19605_, _19603_);
  and (_19607_, _03067_, _02019_);
  nor (_19608_, _19607_, _02853_);
  nand (_19609_, _19608_, _19606_);
  and (_19610_, _04637_, _02853_);
  nor (_19612_, _19610_, _04984_);
  and (_19613_, _19612_, _19609_);
  and (_19614_, _05004_, _04997_);
  not (_19615_, _19614_);
  nor (_19616_, _05005_, _04985_);
  and (_19617_, _19616_, _19615_);
  or (_19618_, _19617_, _19613_);
  and (_19619_, _19618_, _19416_);
  and (_19620_, _04636_, _01919_);
  or (_19621_, _19620_, _01650_);
  or (_19623_, _19621_, _19619_);
  and (_19624_, _03064_, _01650_);
  nor (_19625_, _19624_, _05026_);
  nand (_19626_, _19625_, _19623_);
  and (_19627_, _05038_, _04636_);
  nor (_19628_, _19446_, _05038_);
  or (_19629_, _19628_, _19627_);
  and (_19630_, _19629_, _05026_);
  nor (_19631_, _19630_, _05031_);
  and (_19632_, _19631_, _19626_);
  or (_19634_, _19632_, _19415_);
  nand (_19635_, _19634_, _05050_);
  and (_19636_, _05047_, _04637_);
  nor (_19637_, _19636_, _02018_);
  and (_19638_, _19637_, _19635_);
  and (_19639_, _03067_, _02018_);
  or (_19640_, _19639_, _02135_);
  nor (_19641_, _19640_, _19638_);
  and (_19642_, _04637_, _02135_);
  or (_19643_, _19642_, _19641_);
  nand (_19645_, _19643_, _17617_);
  and (_19646_, _03064_, _01653_);
  nor (_19647_, _19646_, _05059_);
  nand (_19648_, _19647_, _19645_);
  and (_19649_, _05040_, _04636_);
  nor (_19650_, _19446_, _05040_);
  or (_19651_, _19650_, _19649_);
  and (_19652_, _19651_, _05059_);
  nor (_19653_, _19652_, _05069_);
  and (_19654_, _19653_, _19648_);
  or (_19656_, _19654_, _19414_);
  nand (_19657_, _19656_, _05077_);
  and (_19658_, _04637_, _05072_);
  nor (_19659_, _19658_, _02039_);
  and (_19660_, _19659_, _19657_);
  and (_19661_, _03067_, _02039_);
  or (_19662_, _19661_, _02130_);
  nor (_19663_, _19662_, _19660_);
  and (_19664_, _04637_, _02130_);
  or (_19665_, _19664_, _19663_);
  nand (_19667_, _19665_, _17614_);
  and (_19668_, _03064_, _01666_);
  nor (_19669_, _19668_, _05086_);
  nand (_19670_, _19669_, _19667_);
  and (_19671_, _19446_, _05092_);
  nor (_19672_, _04636_, _05092_);
  nor (_19673_, _19672_, _05087_);
  not (_19674_, _19673_);
  nor (_19675_, _19674_, _19671_);
  nor (_19676_, _19675_, _05097_);
  and (_19678_, _19676_, _19670_);
  or (_19679_, _19678_, _19413_);
  nand (_19680_, _19679_, _05105_);
  and (_19681_, _05101_, _04637_);
  nor (_19682_, _19681_, _02016_);
  and (_19683_, _19682_, _19680_);
  and (_19684_, _03067_, _02016_);
  or (_19685_, _19684_, _02126_);
  nor (_19686_, _19685_, _19683_);
  and (_19687_, _04637_, _02126_);
  or (_19689_, _19687_, _19686_);
  nand (_19690_, _19689_, _17611_);
  and (_19691_, _03064_, _01663_);
  nor (_19692_, _19691_, _05114_);
  nand (_19693_, _19692_, _19690_);
  and (_19694_, _19446_, \oc8051_golden_model_1.PSW [7]);
  nor (_19695_, _04636_, \oc8051_golden_model_1.PSW [7]);
  nor (_19696_, _19695_, _05115_);
  not (_19697_, _19696_);
  nor (_19698_, _19697_, _19694_);
  nor (_19700_, _19698_, _05141_);
  and (_19701_, _19700_, _19693_);
  or (_19702_, _19701_, _19411_);
  nand (_19703_, _19702_, _05147_);
  and (_19704_, _04637_, _02273_);
  nor (_19705_, _19704_, _05145_);
  nand (_19706_, _19705_, _19703_);
  and (_19707_, _19402_, _05145_);
  nor (_19708_, _19707_, _02146_);
  and (_19709_, _19708_, _19706_);
  or (_19711_, _19709_, _19410_);
  nand (_19712_, _19711_, _05157_);
  and (_19713_, _03064_, _01660_);
  nor (_19714_, _19713_, _02015_);
  nand (_19715_, _19714_, _19712_);
  and (_19716_, _19425_, _05386_);
  nor (_19717_, _05386_, _03067_);
  or (_19718_, _19717_, _02153_);
  nor (_19719_, _19718_, _19716_);
  nor (_19720_, _19719_, _05161_);
  and (_19722_, _19720_, _19715_);
  or (_19723_, _19722_, _19408_);
  nand (_19724_, _19723_, _05398_);
  and (_19725_, _04637_, _02788_);
  nor (_19726_, _19725_, _05396_);
  nand (_19727_, _19726_, _19724_);
  and (_19728_, _19402_, _05396_);
  nor (_19729_, _19728_, _01585_);
  and (_19730_, _19729_, _19727_);
  or (_19731_, _19730_, _19407_);
  nand (_19733_, _19731_, _05407_);
  and (_19734_, _03064_, _01581_);
  nor (_19735_, _19734_, _02022_);
  nand (_19736_, _19735_, _19733_);
  and (_19737_, _05386_, _03068_);
  nor (_19738_, _19436_, _05386_);
  nor (_19739_, _19738_, _19737_);
  and (_19740_, _19739_, _02022_);
  nor (_19741_, _19740_, _05419_);
  nand (_19742_, _19741_, _19736_);
  nor (_19744_, _19402_, _05418_);
  nor (_19745_, _19744_, _02164_);
  and (_19746_, _19745_, _19742_);
  or (_19747_, _19746_, _19406_);
  nand (_19748_, _19747_, _05430_);
  and (_19749_, _19402_, _05426_);
  nor (_19750_, _19749_, _06467_);
  nand (_19751_, _19750_, _19748_);
  and (_19752_, _06467_, _03064_);
  nor (_19753_, _19752_, _02025_);
  nand (_19755_, _19753_, _19751_);
  and (_19756_, _19739_, _02025_);
  nor (_19757_, _19756_, _05446_);
  nand (_19758_, _19757_, _19755_);
  nor (_19759_, _19402_, _05445_);
  nor (_19760_, _19759_, _01594_);
  and (_19761_, _19760_, _19758_);
  or (_19762_, _19761_, _19405_);
  nand (_19763_, _19762_, _05457_);
  and (_19764_, _19402_, _05453_);
  nor (_19766_, _19764_, _17605_);
  nand (_19767_, _19766_, _19763_);
  and (_19768_, _17605_, _03064_);
  nor (_19769_, _19768_, _05464_);
  nand (_19770_, _19769_, _19767_);
  and (_19771_, _19770_, _19404_);
  nand (_19772_, _19771_, _26505_);
  or (_19773_, _26505_, \oc8051_golden_model_1.PC [5]);
  and (_19774_, _19773_, _25964_);
  and (_27921_, _19774_, _19772_);
  nor (_19776_, _02791_, \oc8051_golden_model_1.PC [6]);
  nor (_19777_, _19776_, _02792_);
  and (_19778_, _19777_, _05464_);
  not (_19779_, _19778_);
  and (_19780_, _06467_, _03025_);
  not (_19781_, _01930_);
  and (_19782_, _04874_, _03028_);
  and (_19783_, _03135_, _03033_);
  nor (_19784_, _19783_, _03136_);
  not (_19785_, _19784_);
  nor (_19787_, _19785_, _04874_);
  nor (_19788_, _19787_, _19782_);
  or (_19789_, _19788_, _02378_);
  and (_19790_, _04628_, _01959_);
  or (_19791_, _04551_, _03028_);
  or (_19792_, _19784_, _04553_);
  and (_19793_, _19792_, _19791_);
  nor (_19794_, _19793_, _02438_);
  or (_19795_, _04707_, _04629_);
  and (_19796_, _04666_, _04633_);
  nor (_19798_, _19796_, _04667_);
  nand (_19799_, _19798_, _04707_);
  and (_19800_, _19799_, _04557_);
  nand (_19801_, _19800_, _19795_);
  and (_19802_, _03025_, _04568_);
  and (_19803_, _04571_, _04629_);
  nor (_19804_, _19803_, _04559_);
  and (_19805_, _18340_, \oc8051_golden_model_1.PC [6]);
  or (_19806_, _19805_, _04571_);
  and (_19807_, _19806_, _19804_);
  not (_19809_, _19777_);
  nor (_19810_, _19809_, _04561_);
  or (_19811_, _19810_, _04568_);
  nor (_19812_, _19811_, _19807_);
  nor (_19813_, _19812_, _04563_);
  not (_19814_, _19813_);
  nor (_19815_, _19814_, _19802_);
  and (_19816_, _19777_, _04563_);
  or (_19817_, _19816_, _01971_);
  or (_19818_, _19817_, _19815_);
  nand (_19820_, _04629_, _01971_);
  and (_19821_, _19820_, _19818_);
  and (_19822_, _19821_, _17894_);
  and (_19823_, _19777_, _04562_);
  or (_19824_, _19823_, _19822_);
  and (_19825_, _19824_, _01627_);
  nor (_19826_, _03025_, _01627_);
  nor (_19827_, _19826_, _04557_);
  not (_19828_, _19827_);
  nor (_19829_, _19828_, _19825_);
  nor (_19831_, _19829_, _04715_);
  nand (_19832_, _19831_, _19801_);
  and (_19833_, _19777_, _04715_);
  nor (_19834_, _19833_, _01969_);
  and (_19835_, _19834_, _19832_);
  or (_19836_, _19835_, _19794_);
  nand (_19837_, _19836_, _17940_);
  and (_19838_, _19809_, _04094_);
  nor (_19839_, _19838_, _01959_);
  and (_19840_, _19839_, _19837_);
  or (_19842_, _19840_, _19790_);
  and (_19843_, _19842_, _01621_);
  nor (_19844_, _03025_, _01621_);
  or (_19845_, _19844_, _01967_);
  or (_19846_, _19845_, _19843_);
  and (_19847_, _04629_, _01967_);
  nor (_19848_, _19847_, _04725_);
  nand (_19849_, _19848_, _19846_);
  and (_19850_, _19777_, _04725_);
  nor (_19851_, _19850_, _01963_);
  nand (_19853_, _19851_, _19849_);
  and (_19854_, _04629_, _01963_);
  nor (_19855_, _19854_, _04734_);
  and (_19856_, _19855_, _19853_);
  and (_19857_, _19777_, _04734_);
  or (_19858_, _19857_, _01957_);
  or (_19859_, _19858_, _19856_);
  and (_19860_, _04629_, _01957_);
  nor (_19861_, _19860_, _17638_);
  and (_19862_, _19861_, _19859_);
  nor (_19864_, _03025_, _01630_);
  or (_19865_, _19864_, _19862_);
  nand (_19866_, _19865_, _02457_);
  and (_19867_, _04628_, _01953_);
  nor (_19868_, _19867_, _04089_);
  and (_19869_, _19868_, _19866_);
  and (_19870_, _04085_, _03028_);
  nor (_19871_, _19785_, _04085_);
  or (_19872_, _19871_, _19870_);
  nor (_19873_, _19872_, _04090_);
  or (_19875_, _19873_, _19869_);
  and (_19876_, _19875_, _03187_);
  and (_19877_, _03909_, _03028_);
  nor (_19878_, _19785_, _03909_);
  or (_19879_, _19878_, _03187_);
  nor (_19880_, _19879_, _19877_);
  or (_19881_, _19880_, _19876_);
  or (_19882_, _19881_, _01951_);
  and (_19883_, _19882_, _19789_);
  or (_19884_, _19883_, _03179_);
  nand (_19886_, _03028_, _02912_);
  nand (_19887_, _19784_, _19160_);
  and (_19888_, _19887_, _19886_);
  or (_19889_, _19888_, _04749_);
  and (_19890_, _19889_, _19884_);
  or (_19891_, _19890_, _02880_);
  nand (_19892_, _19777_, _02880_);
  and (_19893_, _19892_, _19891_);
  nand (_19894_, _19893_, _04885_);
  and (_19895_, _04629_, _01946_);
  nor (_19897_, _19895_, _06393_);
  nand (_19898_, _19897_, _19894_);
  nor (_19899_, _03025_, _01632_);
  nor (_19900_, _19899_, _18009_);
  nand (_19901_, _19900_, _19898_);
  nor (_19902_, _04897_, _04628_);
  nor (_19903_, _19902_, _04908_);
  nand (_19904_, _19903_, _19901_);
  nor (_19905_, _19809_, _04905_);
  nor (_19906_, _19905_, _01931_);
  nand (_19908_, _19906_, _19904_);
  and (_19909_, _04629_, _01931_);
  nor (_19910_, _19909_, _17710_);
  and (_19911_, _19910_, _19908_);
  nor (_19912_, _03025_, _01618_);
  or (_19913_, _19912_, _19911_);
  and (_19914_, _19913_, _19781_);
  and (_19915_, _04628_, _01930_);
  or (_19916_, _19915_, _19914_);
  and (_19917_, _19916_, _04928_);
  nor (_19919_, _19809_, _04928_);
  or (_19920_, _19919_, _19917_);
  and (_19921_, _19920_, _04937_);
  and (_19922_, _04628_, _04932_);
  or (_19923_, _19922_, _19921_);
  and (_19924_, _19923_, _01616_);
  and (_19925_, _19777_, _01611_);
  or (_19926_, _19925_, _01924_);
  or (_19927_, _19926_, _19924_);
  and (_19928_, _04629_, _01924_);
  nor (_19930_, _19928_, _01606_);
  nand (_19931_, _19930_, _19927_);
  nor (_19932_, _03025_, _07270_);
  nor (_19933_, _19932_, _02001_);
  nand (_19934_, _19933_, _19931_);
  and (_19935_, _03029_, _02001_);
  nor (_19936_, _19935_, _04953_);
  nand (_19937_, _19936_, _19934_);
  nor (_19938_, _04952_, _04629_);
  nor (_19939_, _19938_, _01602_);
  and (_19941_, _19939_, _19937_);
  nor (_19942_, _04960_, _03029_);
  nor (_19943_, _19942_, _17728_);
  or (_19944_, _19943_, _19941_);
  and (_19945_, _19777_, _04960_);
  nor (_19946_, _19945_, _01920_);
  nand (_19947_, _19946_, _19944_);
  and (_19948_, _04629_, _01920_);
  nor (_19949_, _19948_, _01654_);
  nand (_19950_, _19949_, _19947_);
  nor (_19952_, _03025_, _17739_);
  nor (_19953_, _19952_, _04968_);
  nand (_19954_, _19953_, _19950_);
  nor (_19955_, _19798_, _04969_);
  nor (_19956_, _19955_, _02859_);
  and (_19957_, _19956_, _19954_);
  and (_19958_, _02859_, _04628_);
  or (_19959_, _19958_, _02019_);
  or (_19960_, _19959_, _19957_);
  and (_19961_, _03029_, _02019_);
  nor (_19963_, _19961_, _02853_);
  nand (_19964_, _19963_, _19960_);
  and (_19965_, _04628_, _02853_);
  nor (_19966_, _19965_, _04984_);
  nand (_19967_, _19966_, _19964_);
  and (_19968_, _05006_, _04993_);
  nor (_19969_, _19968_, _05007_);
  nor (_19970_, _19969_, _04985_);
  nor (_19971_, _19970_, _01919_);
  nand (_19972_, _19971_, _19967_);
  and (_19974_, _04628_, _01919_);
  nor (_19975_, _19974_, _01650_);
  nand (_19976_, _19975_, _19972_);
  and (_19977_, _03025_, _01650_);
  nor (_19978_, _19977_, _05026_);
  nand (_19979_, _19978_, _19976_);
  and (_19980_, _05038_, _04628_);
  and (_19981_, _19798_, _05040_);
  or (_19982_, _19981_, _19980_);
  and (_19983_, _19982_, _05026_);
  nor (_19985_, _19983_, _05031_);
  nand (_19986_, _19985_, _19979_);
  nor (_19987_, _19777_, _02830_);
  nor (_19988_, _19987_, _05047_);
  and (_19989_, _19988_, _19986_);
  and (_19990_, _05047_, _04628_);
  or (_19991_, _19990_, _02018_);
  or (_19992_, _19991_, _19989_);
  and (_19993_, _03029_, _02018_);
  nor (_19994_, _19993_, _02135_);
  and (_19996_, _19994_, _19992_);
  and (_19997_, _04628_, _02135_);
  or (_19998_, _19997_, _01653_);
  or (_19999_, _19998_, _19996_);
  and (_20000_, _03025_, _01653_);
  nor (_20001_, _20000_, _05059_);
  nand (_20002_, _20001_, _19999_);
  and (_20003_, _05040_, _04628_);
  and (_20004_, _19798_, _05038_);
  or (_20005_, _20004_, _20003_);
  and (_20007_, _20005_, _05059_);
  nor (_20008_, _20007_, _05069_);
  nand (_20009_, _20008_, _20002_);
  and (_20010_, _19809_, _05069_);
  nor (_20011_, _20010_, _05072_);
  and (_20012_, _20011_, _20009_);
  and (_20013_, _04628_, _05072_);
  or (_20014_, _20013_, _20012_);
  and (_20015_, _20014_, _05076_);
  and (_20016_, _03028_, _02039_);
  or (_20018_, _20016_, _02130_);
  nor (_20019_, _20018_, _20015_);
  and (_20020_, _04629_, _02130_);
  or (_20021_, _20020_, _20019_);
  nand (_20022_, _20021_, _17614_);
  and (_20023_, _03025_, _01666_);
  nor (_20024_, _20023_, _05086_);
  nand (_20025_, _20024_, _20022_);
  nor (_20026_, _19798_, \oc8051_golden_model_1.PSW [7]);
  nor (_20027_, _04628_, _05092_);
  nor (_20029_, _20027_, _05087_);
  not (_20030_, _20029_);
  nor (_20031_, _20030_, _20026_);
  nor (_20032_, _20031_, _05097_);
  nand (_20033_, _20032_, _20025_);
  and (_20034_, _19809_, _05097_);
  nor (_20035_, _20034_, _05101_);
  and (_20036_, _20035_, _20033_);
  and (_20037_, _05101_, _04628_);
  or (_20038_, _20037_, _20036_);
  nand (_20040_, _20038_, _05104_);
  and (_20041_, _03028_, _02016_);
  nor (_20042_, _20041_, _02126_);
  and (_20043_, _20042_, _20040_);
  and (_20044_, _04629_, _02126_);
  or (_20045_, _20044_, _20043_);
  nand (_20046_, _20045_, _17611_);
  and (_20047_, _03025_, _01663_);
  nor (_20048_, _20047_, _05114_);
  nand (_20049_, _20048_, _20046_);
  nor (_20051_, _19798_, _05092_);
  nor (_20052_, _04628_, \oc8051_golden_model_1.PSW [7]);
  nor (_20053_, _20052_, _05115_);
  not (_20054_, _20053_);
  nor (_20055_, _20054_, _20051_);
  nor (_20056_, _20055_, _05141_);
  nand (_20057_, _20056_, _20049_);
  nor (_20058_, _19777_, _05139_);
  nor (_20059_, _20058_, _02273_);
  and (_20060_, _20059_, _20057_);
  and (_20062_, _04628_, _02273_);
  or (_20063_, _20062_, _20060_);
  and (_20064_, _20063_, _05146_);
  and (_20065_, _19777_, _05145_);
  or (_20066_, _20065_, _20064_);
  nand (_20067_, _20066_, _02718_);
  and (_20068_, _03748_, _02146_);
  nor (_20069_, _20068_, _01660_);
  nand (_20070_, _20069_, _20067_);
  and (_20071_, _03025_, _01660_);
  nor (_20073_, _20071_, _02015_);
  nand (_20074_, _20073_, _20070_);
  nor (_20075_, _05386_, _03028_);
  and (_20076_, _19785_, _05386_);
  or (_20077_, _20076_, _02153_);
  nor (_20078_, _20077_, _20075_);
  nor (_20079_, _20078_, _05161_);
  nand (_20080_, _20079_, _20074_);
  nor (_20081_, _19777_, _02818_);
  nor (_20082_, _20081_, _02788_);
  and (_20084_, _20082_, _20080_);
  and (_20085_, _04628_, _02788_);
  or (_20086_, _20085_, _20084_);
  nand (_20087_, _20086_, _05397_);
  and (_20088_, _19777_, _05396_);
  nor (_20089_, _20088_, _01585_);
  nand (_20090_, _20089_, _20087_);
  nor (_20091_, _03748_, _01596_);
  nor (_20092_, _20091_, _01581_);
  nand (_20093_, _20092_, _20090_);
  nor (_20095_, _03025_, _05407_);
  nor (_20096_, _20095_, _02022_);
  and (_20097_, _20096_, _20093_);
  and (_20098_, _05386_, _03029_);
  nor (_20099_, _19784_, _05386_);
  nor (_20100_, _20099_, _20098_);
  nor (_20101_, _20100_, _02558_);
  nor (_20102_, _20101_, _20097_);
  nand (_20103_, _20102_, _05418_);
  nor (_20104_, _19809_, _05418_);
  nor (_20106_, _20104_, _02164_);
  nand (_20107_, _20106_, _20103_);
  and (_20108_, _04629_, _02164_);
  nor (_20109_, _20108_, _05426_);
  nand (_20110_, _20109_, _20107_);
  and (_20111_, _19777_, _05426_);
  nor (_20112_, _20111_, _06467_);
  and (_20113_, _20112_, _20110_);
  or (_20114_, _20113_, _19780_);
  nand (_20115_, _20114_, _02377_);
  nor (_20117_, _20100_, _02377_);
  nor (_20118_, _20117_, _05446_);
  nand (_20119_, _20118_, _20115_);
  nor (_20120_, _19809_, _05445_);
  nor (_20121_, _20120_, _01594_);
  nand (_20122_, _20121_, _20119_);
  and (_20123_, _04629_, _01594_);
  nor (_20124_, _20123_, _05453_);
  nand (_20125_, _20124_, _20122_);
  and (_20126_, _19777_, _05453_);
  nor (_20128_, _20126_, _17605_);
  nand (_20129_, _20128_, _20125_);
  and (_20130_, _17605_, _03025_);
  nor (_20131_, _20130_, _05464_);
  nand (_20132_, _20131_, _20129_);
  and (_20133_, _20132_, _19779_);
  nand (_20134_, _20133_, _26505_);
  or (_20135_, _26505_, \oc8051_golden_model_1.PC [6]);
  and (_20136_, _20135_, _25964_);
  and (_27922_, _20136_, _20134_);
  and (_20138_, _02988_, _02789_);
  and (_20139_, _20138_, \oc8051_golden_model_1.PC [7]);
  nor (_20140_, _20138_, \oc8051_golden_model_1.PC [7]);
  nor (_20141_, _20140_, _20139_);
  and (_20142_, _20141_, _05464_);
  and (_20143_, _04622_, _01594_);
  nor (_20144_, _20141_, _02818_);
  nor (_20145_, _20141_, _05139_);
  not (_20146_, _20141_);
  and (_20147_, _20146_, _05097_);
  and (_20149_, _20146_, _05069_);
  nor (_20150_, _20141_, _02830_);
  and (_20151_, _04623_, _01924_);
  nor (_20152_, _20141_, _04928_);
  nor (_20153_, _02943_, _01632_);
  and (_20154_, _20146_, _02880_);
  and (_20155_, _04085_, _02991_);
  or (_20156_, _02993_, _02994_);
  not (_20157_, _20156_);
  nor (_20158_, _20157_, _03137_);
  and (_20160_, _20157_, _03137_);
  nor (_20161_, _20160_, _20158_);
  nor (_20162_, _20161_, _04085_);
  or (_20163_, _20162_, _20155_);
  nor (_20164_, _20163_, _04090_);
  and (_20165_, _04553_, _02991_);
  not (_20166_, _20161_);
  and (_20167_, _20166_, _04551_);
  or (_20168_, _20167_, _02438_);
  or (_20169_, _20168_, _20165_);
  and (_20171_, _04710_, _04622_);
  or (_20172_, _04624_, _04625_);
  not (_20173_, _20172_);
  nor (_20174_, _20173_, _04668_);
  and (_20175_, _20173_, _04668_);
  nor (_20176_, _20175_, _20174_);
  nor (_20177_, _20176_, _04710_);
  or (_20178_, _20177_, _20171_);
  nor (_20179_, _20178_, _04709_);
  and (_20180_, _20146_, _04563_);
  nor (_20182_, _02943_, _01625_);
  and (_20183_, _04571_, _04623_);
  nor (_20184_, _20183_, _04559_);
  and (_20185_, _18340_, \oc8051_golden_model_1.PC [7]);
  or (_20186_, _20185_, _04571_);
  and (_20187_, _20186_, _20184_);
  nor (_20188_, _20146_, _04561_);
  or (_20189_, _20188_, _04563_);
  or (_20190_, _20189_, _20187_);
  and (_20191_, _20190_, _01625_);
  nor (_20193_, _20191_, _20182_);
  or (_20194_, _20193_, _01971_);
  nor (_20195_, _20194_, _20180_);
  and (_20196_, _04622_, _01971_);
  or (_20197_, _20196_, _20195_);
  and (_20198_, _20197_, _17894_);
  and (_20199_, _20141_, _04562_);
  or (_20200_, _20199_, _20198_);
  and (_20201_, _20200_, _01627_);
  nor (_20202_, _02943_, _01627_);
  nor (_20204_, _20202_, _04557_);
  not (_20205_, _20204_);
  nor (_20206_, _20205_, _20201_);
  or (_20207_, _20206_, _04715_);
  nor (_20208_, _20207_, _20179_);
  and (_20209_, _20141_, _04715_);
  or (_20210_, _20209_, _01969_);
  or (_20211_, _20210_, _20208_);
  and (_20212_, _20211_, _20169_);
  nor (_20213_, _20212_, _04094_);
  and (_20215_, _20146_, _04094_);
  nor (_20216_, _20215_, _01959_);
  not (_20217_, _20216_);
  nor (_20218_, _20217_, _20213_);
  and (_20219_, _04622_, _01959_);
  nor (_20220_, _20219_, _20218_);
  or (_20221_, _20220_, _06363_);
  or (_20222_, _02943_, _01621_);
  and (_20223_, _20222_, _20221_);
  or (_20224_, _20223_, _01967_);
  and (_20226_, _04622_, _01967_);
  nor (_20227_, _20226_, _04725_);
  nand (_20228_, _20227_, _20224_);
  and (_20229_, _20146_, _04725_);
  nor (_20230_, _20229_, _01963_);
  nand (_20231_, _20230_, _20228_);
  and (_20232_, _04622_, _01963_);
  nor (_20233_, _20232_, _04734_);
  nand (_20234_, _20233_, _20231_);
  and (_20235_, _20146_, _04734_);
  nor (_20237_, _20235_, _01957_);
  nand (_20238_, _20237_, _20234_);
  and (_20239_, _04622_, _01957_);
  nor (_20240_, _20239_, _17638_);
  nand (_20241_, _20240_, _20238_);
  and (_20242_, _02943_, _17638_);
  nor (_20243_, _20242_, _01953_);
  nand (_20244_, _20243_, _20241_);
  and (_20245_, _04622_, _01953_);
  nor (_20246_, _20245_, _04089_);
  and (_20248_, _20246_, _20244_);
  or (_20249_, _20248_, _20164_);
  and (_20250_, _20249_, _03187_);
  nor (_20251_, _20166_, _03909_);
  and (_20252_, _03909_, _02992_);
  nor (_20253_, _20252_, _20251_);
  nor (_20254_, _20253_, _03187_);
  or (_20255_, _20254_, _20250_);
  or (_20256_, _20255_, _01951_);
  nor (_20257_, _20161_, _04874_);
  and (_20259_, _04874_, _02991_);
  nor (_20260_, _20259_, _20257_);
  or (_20261_, _20260_, _02378_);
  and (_20262_, _20261_, _20256_);
  or (_20263_, _20262_, _03179_);
  and (_20264_, _02991_, _02912_);
  nor (_20265_, _20161_, _02912_);
  or (_20266_, _20265_, _20264_);
  and (_20267_, _20266_, _03179_);
  nor (_20268_, _20267_, _02880_);
  and (_20270_, _20268_, _20263_);
  or (_20271_, _20270_, _20154_);
  nand (_20272_, _20271_, _04885_);
  and (_20273_, _04623_, _01946_);
  nor (_20274_, _20273_, _06393_);
  nand (_20275_, _20274_, _20272_);
  nand (_20276_, _20275_, _04897_);
  nor (_20277_, _20276_, _20153_);
  nor (_20278_, _04897_, _04622_);
  or (_20279_, _20278_, _20277_);
  nand (_20281_, _20279_, _04905_);
  nor (_20282_, _20141_, _04905_);
  nor (_20283_, _20282_, _01931_);
  nand (_20284_, _20283_, _20281_);
  and (_20285_, _04622_, _01931_);
  nor (_20286_, _20285_, _17710_);
  nand (_20287_, _20286_, _20284_);
  and (_20288_, _02943_, _17710_);
  nor (_20289_, _20288_, _01930_);
  nand (_20290_, _20289_, _20287_);
  and (_20292_, _04622_, _01930_);
  nor (_20293_, _20292_, _04933_);
  and (_20294_, _20293_, _20290_);
  or (_20295_, _20294_, _20152_);
  nand (_20296_, _20295_, _04937_);
  and (_20297_, _04623_, _04932_);
  nor (_20298_, _20297_, _01611_);
  nand (_20299_, _20298_, _20296_);
  and (_20300_, _20141_, _01611_);
  nor (_20301_, _20300_, _01924_);
  and (_20303_, _20301_, _20299_);
  or (_20304_, _20303_, _20151_);
  nand (_20305_, _20304_, _07270_);
  and (_20306_, _02943_, _01606_);
  nor (_20307_, _20306_, _02001_);
  nand (_20308_, _20307_, _20305_);
  and (_20309_, _02991_, _02001_);
  nor (_20310_, _20309_, _04953_);
  nand (_20311_, _20310_, _20308_);
  nor (_20312_, _04952_, _04622_);
  nor (_20314_, _20312_, _01602_);
  and (_20315_, _20314_, _20311_);
  and (_20316_, _02991_, _01602_);
  or (_20317_, _20316_, _04960_);
  or (_20318_, _20317_, _20315_);
  and (_20319_, _20146_, _04960_);
  nor (_20320_, _20319_, _01920_);
  nand (_20321_, _20320_, _20318_);
  and (_20322_, _04622_, _01920_);
  nor (_20323_, _20322_, _01654_);
  nand (_20325_, _20323_, _20321_);
  and (_20326_, _02943_, _01654_);
  nor (_20327_, _20326_, _04968_);
  nand (_20328_, _20327_, _20325_);
  nor (_20329_, _20176_, _04969_);
  nor (_20330_, _20329_, _02859_);
  nand (_20331_, _20330_, _20328_);
  and (_20332_, _02859_, _04623_);
  nor (_20333_, _20332_, _02019_);
  nand (_20334_, _20333_, _20331_);
  and (_20336_, _02991_, _02019_);
  nor (_20337_, _20336_, _02853_);
  nand (_20338_, _20337_, _20334_);
  and (_20339_, _04623_, _02853_);
  nor (_20340_, _20339_, _04984_);
  nand (_20341_, _20340_, _20338_);
  or (_20342_, _04988_, _04989_);
  nor (_20343_, _20342_, _05008_);
  and (_20344_, _20342_, _05008_);
  or (_20345_, _20344_, _04985_);
  or (_20347_, _20345_, _20343_);
  nand (_20348_, _20347_, _20341_);
  and (_20349_, _20348_, _19416_);
  and (_20350_, _04622_, _01919_);
  or (_20351_, _20350_, _01650_);
  or (_20352_, _20351_, _20349_);
  and (_20353_, _02943_, _01650_);
  nor (_20354_, _20353_, _05026_);
  nand (_20355_, _20354_, _20352_);
  and (_20356_, _05038_, _04622_);
  nor (_20358_, _20176_, _05038_);
  or (_20359_, _20358_, _20356_);
  and (_20360_, _20359_, _05026_);
  nor (_20361_, _20360_, _05031_);
  and (_20362_, _20361_, _20355_);
  or (_20363_, _20362_, _20150_);
  nand (_20364_, _20363_, _05050_);
  and (_20365_, _05047_, _04623_);
  nor (_20366_, _20365_, _02018_);
  and (_20367_, _20366_, _20364_);
  and (_20369_, _02991_, _02018_);
  or (_20370_, _20369_, _02135_);
  nor (_20371_, _20370_, _20367_);
  and (_20372_, _04623_, _02135_);
  or (_20373_, _20372_, _20371_);
  nand (_20374_, _20373_, _17617_);
  and (_20375_, _02943_, _01653_);
  nor (_20376_, _20375_, _05059_);
  nand (_20377_, _20376_, _20374_);
  and (_20378_, _05040_, _04622_);
  nor (_20380_, _20176_, _05040_);
  or (_20381_, _20380_, _20378_);
  and (_20382_, _20381_, _05059_);
  nor (_20383_, _20382_, _05069_);
  and (_20384_, _20383_, _20377_);
  or (_20385_, _20384_, _20149_);
  nand (_20386_, _20385_, _05077_);
  and (_20387_, _04623_, _05072_);
  nor (_20388_, _20387_, _02039_);
  and (_20389_, _20388_, _20386_);
  and (_20391_, _02991_, _02039_);
  or (_20392_, _20391_, _02130_);
  nor (_20393_, _20392_, _20389_);
  and (_20394_, _04623_, _02130_);
  or (_20395_, _20394_, _20393_);
  nand (_20396_, _20395_, _17614_);
  and (_20397_, _02943_, _01666_);
  nor (_20398_, _20397_, _05086_);
  nand (_20399_, _20398_, _20396_);
  and (_20400_, _20176_, _05092_);
  nor (_20402_, _04622_, _05092_);
  nor (_20403_, _20402_, _05087_);
  not (_20404_, _20403_);
  nor (_20405_, _20404_, _20400_);
  nor (_20406_, _20405_, _05097_);
  and (_20407_, _20406_, _20399_);
  or (_20408_, _20407_, _20147_);
  nand (_20409_, _20408_, _05105_);
  and (_20410_, _05101_, _04623_);
  nor (_20411_, _20410_, _02016_);
  and (_20413_, _20411_, _20409_);
  and (_20414_, _02991_, _02016_);
  or (_20415_, _20414_, _02126_);
  nor (_20416_, _20415_, _20413_);
  and (_20417_, _04623_, _02126_);
  or (_20418_, _20417_, _20416_);
  nand (_20419_, _20418_, _17611_);
  and (_20420_, _02943_, _01663_);
  nor (_20421_, _20420_, _05114_);
  nand (_20422_, _20421_, _20419_);
  and (_20424_, _04622_, _05092_);
  nor (_20425_, _20176_, _05092_);
  or (_20426_, _20425_, _20424_);
  and (_20427_, _20426_, _05114_);
  nor (_20428_, _20427_, _05141_);
  and (_20429_, _20428_, _20422_);
  or (_20430_, _20429_, _20145_);
  nand (_20431_, _20430_, _05147_);
  and (_20432_, _04623_, _02273_);
  nor (_20433_, _20432_, _05145_);
  nand (_20435_, _20433_, _20431_);
  and (_20436_, _20141_, _05145_);
  nor (_20437_, _20436_, _02146_);
  and (_20438_, _20437_, _20435_);
  nor (_20439_, _03796_, _02718_);
  or (_20440_, _20439_, _20438_);
  nand (_20441_, _20440_, _05157_);
  and (_20442_, _02943_, _01660_);
  nor (_20443_, _20442_, _02015_);
  nand (_20444_, _20443_, _20441_);
  and (_20446_, _20161_, _05386_);
  nor (_20447_, _05386_, _02991_);
  or (_20448_, _20447_, _02153_);
  or (_20449_, _20448_, _20446_);
  and (_20450_, _20449_, _02818_);
  and (_20451_, _20450_, _20444_);
  or (_20452_, _20451_, _20144_);
  nand (_20453_, _20452_, _05398_);
  and (_20454_, _04623_, _02788_);
  nor (_20455_, _20454_, _05396_);
  nand (_20457_, _20455_, _20453_);
  and (_20458_, _20141_, _05396_);
  nor (_20459_, _20458_, _01585_);
  and (_20460_, _20459_, _20457_);
  nor (_20461_, _03796_, _01596_);
  or (_20462_, _20461_, _20460_);
  nand (_20463_, _20462_, _05407_);
  and (_20464_, _02943_, _01581_);
  nor (_20465_, _20464_, _02022_);
  nand (_20466_, _20465_, _20463_);
  and (_20468_, _05386_, _02992_);
  nor (_20469_, _20166_, _05386_);
  nor (_20470_, _20469_, _20468_);
  and (_20471_, _20470_, _02022_);
  nor (_20472_, _20471_, _05419_);
  nand (_20473_, _20472_, _20466_);
  nor (_20474_, _20141_, _05418_);
  nor (_20475_, _20474_, _02164_);
  nand (_20476_, _20475_, _20473_);
  and (_20477_, _04622_, _02164_);
  nor (_20479_, _20477_, _05426_);
  and (_20480_, _20479_, _20476_);
  and (_20481_, _20146_, _05426_);
  or (_20482_, _20481_, _20480_);
  nand (_20483_, _20482_, _06466_);
  and (_20484_, _06467_, _02943_);
  nor (_20485_, _20484_, _02025_);
  nand (_20486_, _20485_, _20483_);
  and (_20487_, _20470_, _02025_);
  nor (_20488_, _20487_, _05446_);
  nand (_20490_, _20488_, _20486_);
  nor (_20491_, _20141_, _05445_);
  nor (_20492_, _20491_, _01594_);
  and (_20493_, _20492_, _20490_);
  or (_20494_, _20493_, _20143_);
  nand (_20495_, _20494_, _05457_);
  and (_20496_, _20141_, _05453_);
  nor (_20497_, _20496_, _17605_);
  nand (_20498_, _20497_, _20495_);
  and (_20499_, _17605_, _02943_);
  nor (_20501_, _20499_, _05464_);
  and (_20502_, _20501_, _20498_);
  or (_20503_, _20502_, _20142_);
  or (_20504_, _20503_, _26506_);
  or (_20505_, _26505_, \oc8051_golden_model_1.PC [7]);
  and (_20506_, _20505_, _25964_);
  and (_27923_, _20506_, _20504_);
  nor (_20507_, _02409_, _05456_);
  nor (_20508_, _02409_, _05429_);
  nor (_20509_, _20139_, \oc8051_golden_model_1.PC [8]);
  and (_20511_, _20139_, \oc8051_golden_model_1.PC [8]);
  nor (_20512_, _20511_, _20509_);
  nor (_20513_, _20512_, _02818_);
  nor (_20514_, _20512_, _05139_);
  not (_20515_, _20512_);
  and (_20516_, _20515_, _05097_);
  and (_20517_, _20515_, _05069_);
  and (_20518_, _03141_, _02018_);
  nor (_20519_, _20512_, _02830_);
  nor (_20520_, _04968_, _01654_);
  nor (_20522_, _20512_, _04928_);
  and (_20523_, _04672_, _01953_);
  and (_20524_, _04672_, _01957_);
  and (_20525_, _04672_, _01967_);
  and (_20526_, _04672_, _01959_);
  and (_20527_, _04553_, _03141_);
  nor (_20528_, _03145_, _03139_);
  nor (_20529_, _20528_, _03146_);
  and (_20530_, _20529_, _04551_);
  or (_20531_, _20530_, _02438_);
  or (_20533_, _20531_, _20527_);
  and (_20534_, _04710_, _04672_);
  nor (_20535_, _04676_, _04670_);
  nor (_20536_, _20535_, _04677_);
  and (_20537_, _20536_, _04707_);
  or (_20538_, _20537_, _20534_);
  nor (_20539_, _20538_, _04709_);
  nor (_20540_, _04571_, _01971_);
  or (_20541_, _20540_, _04673_);
  or (_20542_, _20515_, _04561_);
  and (_20544_, _20515_, _04563_);
  and (_20545_, _05488_, \oc8051_golden_model_1.PC [8]);
  nand (_20546_, _20545_, _04561_);
  and (_20547_, _20546_, _18344_);
  or (_20548_, _20547_, _20544_);
  and (_20549_, _20548_, _20542_);
  or (_20550_, _20549_, _01971_);
  and (_20551_, _20550_, _20541_);
  nor (_20552_, _20551_, _04562_);
  and (_20553_, _20512_, _04562_);
  nor (_20555_, _04557_, _04558_);
  not (_20556_, _20555_);
  nor (_20557_, _20556_, _20553_);
  not (_20558_, _20557_);
  nor (_20559_, _20558_, _20552_);
  or (_20560_, _20559_, _04715_);
  nor (_20561_, _20560_, _20539_);
  and (_20562_, _20512_, _04715_);
  or (_20563_, _20562_, _01969_);
  or (_20564_, _20563_, _20561_);
  and (_20566_, _20564_, _20533_);
  nor (_20567_, _20566_, _04094_);
  and (_20568_, _20515_, _04094_);
  nor (_20569_, _20568_, _01959_);
  not (_20570_, _20569_);
  nor (_20571_, _20570_, _20567_);
  nor (_20572_, _20571_, _20526_);
  nor (_20573_, _20572_, _06363_);
  and (_20574_, _20573_, _05487_);
  or (_20575_, _20574_, _04725_);
  nor (_20577_, _20575_, _20525_);
  and (_20578_, _20515_, _04725_);
  nor (_20579_, _20578_, _01963_);
  not (_20580_, _20579_);
  nor (_20581_, _20580_, _20577_);
  and (_20582_, _04672_, _01963_);
  nor (_20583_, _20582_, _04734_);
  not (_20584_, _20583_);
  nor (_20585_, _20584_, _20581_);
  and (_20586_, _20515_, _04734_);
  nor (_20588_, _20586_, _01957_);
  not (_20589_, _20588_);
  nor (_20590_, _20589_, _20585_);
  nor (_20591_, _20590_, _20524_);
  nor (_20592_, _20591_, _17638_);
  and (_20593_, _20592_, _02457_);
  or (_20594_, _20593_, _04089_);
  nor (_20595_, _20594_, _20523_);
  not (_20596_, _20529_);
  nor (_20597_, _20596_, _04085_);
  not (_20599_, _20597_);
  and (_20600_, _04085_, _03141_);
  nor (_20601_, _20600_, _04090_);
  and (_20602_, _20601_, _20599_);
  nor (_20603_, _20602_, _20595_);
  nor (_20604_, _20603_, _03185_);
  nor (_20605_, _20529_, _03909_);
  and (_20606_, _03909_, _03142_);
  nor (_20607_, _20606_, _20605_);
  nor (_20608_, _20607_, _03187_);
  nor (_20610_, _20608_, _20604_);
  and (_20611_, _20610_, _02378_);
  nor (_20612_, _20596_, _04874_);
  and (_20613_, _04874_, _03141_);
  or (_20614_, _20613_, _20612_);
  and (_20615_, _20614_, _01951_);
  or (_20616_, _20615_, _20611_);
  and (_20617_, _20616_, _04749_);
  and (_20618_, _03141_, _02912_);
  and (_20619_, _20529_, _19160_);
  or (_20621_, _20619_, _20618_);
  and (_20622_, _20621_, _03179_);
  nor (_20623_, _20622_, _20617_);
  or (_20624_, _20623_, _02880_);
  nand (_20625_, _20512_, _02880_);
  and (_20626_, _20625_, _20624_);
  or (_20627_, _20626_, _01946_);
  and (_20628_, _04672_, _01946_);
  not (_20629_, _20628_);
  and (_20630_, _20629_, _04898_);
  and (_20632_, _20630_, _20627_);
  nor (_20633_, _04897_, _04672_);
  or (_20634_, _20633_, _20632_);
  nand (_20635_, _20634_, _04905_);
  nor (_20636_, _20512_, _04905_);
  nor (_20637_, _20636_, _01931_);
  nand (_20638_, _20637_, _20635_);
  and (_20639_, _04672_, _01931_);
  nor (_20640_, _20639_, _17710_);
  nand (_20641_, _20640_, _20638_);
  nand (_20643_, _20641_, _19781_);
  and (_20644_, _04672_, _01930_);
  nor (_20645_, _20644_, _04933_);
  and (_20646_, _20645_, _20643_);
  or (_20647_, _20646_, _20522_);
  nand (_20648_, _20647_, _04937_);
  and (_20649_, _04673_, _04932_);
  nor (_20650_, _20649_, _01611_);
  nand (_20651_, _20650_, _20648_);
  and (_20652_, _20512_, _01611_);
  nor (_20654_, _20652_, _01924_);
  nand (_20655_, _20654_, _20651_);
  nor (_20656_, _02001_, _01606_);
  not (_20657_, _20656_);
  and (_20658_, _04673_, _01924_);
  nor (_20659_, _20658_, _20657_);
  nand (_20660_, _20659_, _20655_);
  and (_20661_, _03141_, _02001_);
  nor (_20662_, _20661_, _04953_);
  nand (_20663_, _20662_, _20660_);
  nor (_20665_, _04952_, _04672_);
  nor (_20666_, _20665_, _01602_);
  and (_20667_, _20666_, _20663_);
  nor (_20668_, _04960_, _03141_);
  nor (_20669_, _20668_, _17728_);
  or (_20670_, _20669_, _20667_);
  and (_20671_, _20515_, _04960_);
  nor (_20672_, _20671_, _01920_);
  and (_20673_, _20672_, _20670_);
  and (_20674_, _04672_, _01920_);
  or (_20676_, _20674_, _20673_);
  nand (_20677_, _20676_, _20520_);
  and (_20678_, _20536_, _04968_);
  nor (_20679_, _20678_, _02859_);
  nand (_20680_, _20679_, _20677_);
  and (_20681_, _02859_, _04673_);
  nor (_20682_, _20681_, _02019_);
  nand (_20683_, _20682_, _20680_);
  and (_20684_, _03141_, _02019_);
  nor (_20685_, _20684_, _02853_);
  nand (_20687_, _20685_, _20683_);
  and (_20688_, _04673_, _02853_);
  nor (_20689_, _20688_, _04984_);
  and (_20690_, _20689_, _20687_);
  nor (_20691_, _05010_, \oc8051_golden_model_1.DPH [0]);
  not (_20692_, _20691_);
  nor (_20693_, _05011_, _04985_);
  and (_20694_, _20693_, _20692_);
  or (_20695_, _20694_, _20690_);
  nand (_20696_, _20695_, _19416_);
  and (_20698_, _04672_, _01919_);
  nor (_20699_, _20698_, _01650_);
  nand (_20700_, _20699_, _20696_);
  nand (_20701_, _20700_, _05027_);
  and (_20702_, _05038_, _04672_);
  and (_20703_, _20536_, _05040_);
  or (_20704_, _20703_, _20702_);
  and (_20705_, _20704_, _05026_);
  nor (_20706_, _20705_, _05031_);
  and (_20707_, _20706_, _20701_);
  or (_20709_, _20707_, _20519_);
  nand (_20710_, _20709_, _05050_);
  and (_20711_, _05047_, _04673_);
  nor (_20712_, _20711_, _02018_);
  and (_20713_, _20712_, _20710_);
  or (_20714_, _20713_, _20518_);
  nand (_20715_, _20714_, _02136_);
  and (_20716_, _04672_, _02135_);
  nor (_20717_, _20716_, _01653_);
  nand (_20718_, _20717_, _20715_);
  nand (_20720_, _20718_, _05060_);
  and (_20721_, _05040_, _04672_);
  and (_20722_, _20536_, _05038_);
  or (_20723_, _20722_, _20721_);
  and (_20724_, _20723_, _05059_);
  nor (_20725_, _20724_, _05069_);
  and (_20726_, _20725_, _20720_);
  or (_20727_, _20726_, _20517_);
  nand (_20728_, _20727_, _05077_);
  and (_20729_, _04673_, _05072_);
  nor (_20731_, _20729_, _02039_);
  nand (_20732_, _20731_, _20728_);
  and (_20733_, _03141_, _02039_);
  nor (_20734_, _20733_, _02130_);
  nand (_20735_, _20734_, _20732_);
  and (_20736_, _04673_, _02130_);
  nor (_20737_, _05086_, _01666_);
  not (_20738_, _20737_);
  nor (_20739_, _20738_, _20736_);
  nand (_20740_, _20739_, _20735_);
  nor (_20742_, _20536_, \oc8051_golden_model_1.PSW [7]);
  nor (_20743_, _04672_, _05092_);
  nor (_20744_, _20743_, _05087_);
  not (_20745_, _20744_);
  nor (_20746_, _20745_, _20742_);
  nor (_20747_, _20746_, _05097_);
  and (_20748_, _20747_, _20740_);
  or (_20749_, _20748_, _20516_);
  nand (_20750_, _20749_, _05105_);
  and (_20751_, _05101_, _04673_);
  nor (_20753_, _20751_, _02016_);
  and (_20754_, _20753_, _20750_);
  and (_20755_, _03141_, _02016_);
  or (_20756_, _20755_, _02126_);
  or (_20757_, _20756_, _20754_);
  and (_20758_, _04673_, _02126_);
  nor (_20759_, _05114_, _01663_);
  not (_20760_, _20759_);
  nor (_20761_, _20760_, _20758_);
  nand (_20762_, _20761_, _20757_);
  and (_20764_, _04672_, _05092_);
  and (_20765_, _20536_, \oc8051_golden_model_1.PSW [7]);
  or (_20766_, _20765_, _20764_);
  and (_20767_, _20766_, _05114_);
  nor (_20768_, _20767_, _05141_);
  and (_20769_, _20768_, _20762_);
  or (_20770_, _20769_, _20514_);
  nand (_20771_, _20770_, _05147_);
  and (_20772_, _04673_, _02273_);
  nor (_20773_, _20772_, _05145_);
  and (_20775_, _20773_, _20771_);
  and (_20776_, _20512_, _05145_);
  or (_20777_, _20776_, _20775_);
  nand (_20778_, _20777_, _02718_);
  and (_20779_, _03334_, _02146_);
  nor (_20780_, _20779_, _01660_);
  nand (_20781_, _20780_, _20778_);
  nand (_20782_, _20781_, _02153_);
  and (_20783_, _20596_, _05386_);
  nor (_20784_, _05386_, _03141_);
  or (_20786_, _20784_, _02153_);
  nor (_20787_, _20786_, _20783_);
  nor (_20788_, _20787_, _05161_);
  and (_20789_, _20788_, _20782_);
  or (_20790_, _20789_, _20513_);
  nand (_20791_, _20790_, _05398_);
  and (_20792_, _04673_, _02788_);
  nor (_20793_, _20792_, _05396_);
  and (_20794_, _20793_, _20791_);
  and (_20795_, _20512_, _05396_);
  or (_20797_, _20795_, _20794_);
  nand (_20798_, _20797_, _01596_);
  and (_20799_, _03334_, _01585_);
  nor (_20800_, _20799_, _01581_);
  nand (_20801_, _20800_, _20798_);
  nand (_20802_, _20801_, _02558_);
  and (_20803_, _05386_, _03142_);
  nor (_20804_, _20529_, _05386_);
  nor (_20805_, _20804_, _20803_);
  and (_20806_, _20805_, _02022_);
  nor (_20808_, _20806_, _05419_);
  nand (_20809_, _20808_, _20802_);
  nor (_20810_, _20512_, _05418_);
  nor (_20811_, _20810_, _02164_);
  nand (_20812_, _20811_, _20809_);
  and (_20813_, _04672_, _02164_);
  nor (_20814_, _20813_, _05426_);
  nand (_20815_, _20814_, _20812_);
  and (_20816_, _20515_, _05426_);
  nor (_20817_, _20816_, _02023_);
  and (_20819_, _20817_, _20815_);
  or (_20820_, _20819_, _20508_);
  nor (_20821_, _02025_, _01670_);
  nand (_20822_, _20821_, _20820_);
  and (_20823_, _20805_, _02025_);
  nor (_20824_, _20823_, _05446_);
  nand (_20825_, _20824_, _20822_);
  nor (_20826_, _20512_, _05445_);
  nor (_20827_, _20826_, _01594_);
  nand (_20828_, _20827_, _20825_);
  and (_20830_, _04672_, _01594_);
  nor (_20831_, _20830_, _05453_);
  nand (_20832_, _20831_, _20828_);
  and (_20833_, _20515_, _05453_);
  nor (_20834_, _20833_, _02026_);
  and (_20835_, _20834_, _20832_);
  or (_20836_, _20835_, _20507_);
  nor (_20837_, _01657_, _05464_);
  nand (_20838_, _20837_, _20836_);
  and (_20839_, _20512_, _05464_);
  not (_20841_, _20839_);
  and (_20842_, _20841_, _20838_);
  nand (_20843_, _20842_, _26505_);
  or (_20844_, _26505_, \oc8051_golden_model_1.PC [8]);
  and (_20845_, _20844_, _25964_);
  and (_27924_, _20845_, _20843_);
  nor (_20846_, _02643_, _05456_);
  nor (_20847_, _02643_, _05429_);
  not (_20848_, \oc8051_golden_model_1.PC [9]);
  and (_20849_, _02835_, _02789_);
  and (_20851_, _20849_, \oc8051_golden_model_1.PC [8]);
  nor (_20852_, _20851_, _20848_);
  and (_20853_, _20851_, _20848_);
  or (_20854_, _20853_, _20852_);
  nor (_20855_, _20854_, _02818_);
  nor (_20856_, _20854_, _05139_);
  and (_20857_, _02983_, _02016_);
  not (_20858_, _20854_);
  and (_20859_, _20858_, _05097_);
  and (_20860_, _02983_, _02039_);
  and (_20862_, _20858_, _05069_);
  and (_20863_, _02983_, _02018_);
  nor (_20864_, _20854_, _02830_);
  and (_20865_, _04615_, _01920_);
  and (_20866_, _04615_, _01930_);
  nor (_20867_, _01930_, _17710_);
  nor (_20868_, _20854_, _04905_);
  and (_20869_, _04615_, _01953_);
  and (_20870_, _04615_, _01967_);
  nor (_20871_, _20540_, _04616_);
  nor (_20873_, _20858_, _04561_);
  and (_20874_, _20858_, _04563_);
  not (_20875_, _18344_);
  nor (_20876_, _04571_, _20848_);
  and (_20877_, _20876_, _04561_);
  nor (_20878_, _20877_, _20875_);
  nor (_20879_, _20878_, _20874_);
  nor (_20880_, _20879_, _20873_);
  nor (_20881_, _20880_, _01971_);
  nor (_20882_, _20881_, _20871_);
  nor (_20884_, _20882_, _04562_);
  and (_20885_, _20854_, _04562_);
  or (_20886_, _20885_, _20556_);
  nor (_20887_, _20886_, _20884_);
  and (_20888_, _04710_, _04615_);
  nor (_20889_, _04677_, _04674_);
  and (_20890_, _20889_, _04619_);
  nor (_20891_, _20889_, _04619_);
  nor (_20892_, _20891_, _20890_);
  nor (_20893_, _20892_, _04710_);
  or (_20895_, _20893_, _20888_);
  nor (_20896_, _20895_, _04709_);
  nor (_20897_, _20896_, _20887_);
  nor (_20898_, _20897_, _04715_);
  and (_20899_, _20858_, _04715_);
  or (_20900_, _20899_, _01969_);
  nor (_20901_, _20900_, _20898_);
  nor (_20902_, _03146_, _03143_);
  and (_20903_, _20902_, _02987_);
  nor (_20904_, _20902_, _02987_);
  nor (_20906_, _20904_, _20903_);
  and (_20907_, _20906_, _04551_);
  and (_20908_, _04553_, _02984_);
  or (_20909_, _20908_, _02438_);
  nor (_20910_, _20909_, _20907_);
  or (_20911_, _20910_, _04094_);
  nor (_20912_, _20911_, _20901_);
  and (_20913_, _20858_, _04094_);
  nor (_20914_, _20913_, _01959_);
  not (_20915_, _20914_);
  nor (_20917_, _20915_, _20912_);
  and (_20918_, _04615_, _01959_);
  or (_20919_, _20918_, _06363_);
  nor (_20920_, _20919_, _20917_);
  nor (_20921_, _20920_, _01967_);
  or (_20922_, _20921_, _04725_);
  nor (_20923_, _20922_, _20870_);
  and (_20924_, _20858_, _04725_);
  nor (_20925_, _20924_, _01963_);
  not (_20926_, _20925_);
  nor (_20928_, _20926_, _20923_);
  and (_20929_, _04615_, _01963_);
  nor (_20930_, _20929_, _04734_);
  not (_20931_, _20930_);
  nor (_20932_, _20931_, _20928_);
  and (_20933_, _20858_, _04734_);
  nor (_20934_, _20933_, _01957_);
  not (_20935_, _20934_);
  nor (_20936_, _20935_, _20932_);
  and (_20937_, _04615_, _01957_);
  or (_20939_, _20937_, _17638_);
  nor (_20940_, _20939_, _20936_);
  nor (_20941_, _20940_, _01953_);
  or (_20942_, _20941_, _04089_);
  nor (_20943_, _20942_, _20869_);
  and (_20944_, _04085_, _02983_);
  nor (_20945_, _20906_, _04085_);
  or (_20946_, _20945_, _04090_);
  nor (_20947_, _20946_, _20944_);
  nor (_20948_, _20947_, _20943_);
  or (_20950_, _20948_, _03185_);
  and (_20951_, _03909_, _02983_);
  nor (_20952_, _20906_, _03909_);
  or (_20953_, _20952_, _03187_);
  or (_20954_, _20953_, _20951_);
  and (_20955_, _20954_, _20950_);
  and (_20956_, _20955_, _02378_);
  and (_20957_, _04874_, _02983_);
  nor (_20958_, _20906_, _04874_);
  or (_20959_, _20958_, _20957_);
  and (_20961_, _20959_, _01951_);
  or (_20962_, _20961_, _20956_);
  and (_20963_, _20962_, _04749_);
  and (_20964_, _02983_, _02912_);
  nor (_20965_, _20906_, _02912_);
  or (_20966_, _20965_, _20964_);
  and (_20967_, _20966_, _03179_);
  or (_20968_, _20967_, _20963_);
  and (_20969_, _20968_, _02881_);
  and (_20970_, _20854_, _02880_);
  or (_20972_, _20970_, _20969_);
  nor (_20973_, _20972_, _01946_);
  and (_20974_, _04898_, _04615_);
  nor (_20975_, _20974_, _04899_);
  nor (_20976_, _20975_, _20973_);
  nor (_20977_, _04897_, _04616_);
  nor (_20978_, _20977_, _04908_);
  not (_20979_, _20978_);
  nor (_20980_, _20979_, _20976_);
  or (_20981_, _20980_, _01931_);
  nor (_20983_, _20981_, _20868_);
  and (_20984_, _04615_, _01931_);
  or (_20985_, _20984_, _20983_);
  and (_20986_, _20985_, _20867_);
  or (_20987_, _20986_, _20866_);
  nand (_20988_, _20987_, _04928_);
  nor (_20989_, _20858_, _04928_);
  nor (_20990_, _20989_, _04932_);
  nand (_20991_, _20990_, _20988_);
  and (_20992_, _04616_, _04932_);
  nor (_20994_, _20992_, _01611_);
  nand (_20995_, _20994_, _20991_);
  and (_20996_, _20854_, _01611_);
  nor (_20997_, _20996_, _01924_);
  nand (_20998_, _20997_, _20995_);
  and (_20999_, _04616_, _01924_);
  nor (_21000_, _20999_, _20657_);
  nand (_21001_, _21000_, _20998_);
  and (_21002_, _02983_, _02001_);
  nor (_21003_, _21002_, _04953_);
  nand (_21005_, _21003_, _21001_);
  nor (_21006_, _04952_, _04615_);
  nor (_21007_, _21006_, _01602_);
  and (_21008_, _21007_, _21005_);
  nor (_21009_, _04960_, _02983_);
  nor (_21010_, _21009_, _17728_);
  or (_21011_, _21010_, _21008_);
  and (_21012_, _20858_, _04960_);
  nor (_21013_, _21012_, _01920_);
  and (_21014_, _21013_, _21011_);
  or (_21016_, _21014_, _20865_);
  nand (_21017_, _21016_, _20520_);
  nor (_21018_, _20892_, _04969_);
  nor (_21019_, _21018_, _02859_);
  nand (_21020_, _21019_, _21017_);
  and (_21021_, _02859_, _04616_);
  nor (_21022_, _21021_, _02019_);
  nand (_21023_, _21022_, _21020_);
  and (_21024_, _02983_, _02019_);
  nor (_21025_, _21024_, _02853_);
  nand (_21027_, _21025_, _21023_);
  and (_21028_, _04616_, _02853_);
  nor (_21029_, _21028_, _04984_);
  and (_21030_, _21029_, _21027_);
  nor (_21031_, _05011_, \oc8051_golden_model_1.DPH [1]);
  not (_21032_, _21031_);
  nor (_21033_, _05012_, _04985_);
  and (_21034_, _21033_, _21032_);
  or (_21035_, _21034_, _21030_);
  nand (_21036_, _21035_, _19416_);
  and (_21038_, _04615_, _01919_);
  nor (_21039_, _21038_, _01650_);
  nand (_21040_, _21039_, _21036_);
  nand (_21041_, _21040_, _05027_);
  and (_21042_, _20892_, _05040_);
  nor (_21043_, _05040_, _04615_);
  nor (_21044_, _21043_, _05027_);
  not (_21045_, _21044_);
  nor (_21046_, _21045_, _21042_);
  nor (_21047_, _21046_, _05031_);
  and (_21049_, _21047_, _21041_);
  or (_21050_, _21049_, _20864_);
  nand (_21051_, _21050_, _05050_);
  and (_21052_, _05047_, _04616_);
  nor (_21053_, _21052_, _02018_);
  and (_21054_, _21053_, _21051_);
  or (_21055_, _21054_, _20863_);
  nand (_21056_, _21055_, _02136_);
  and (_21057_, _04615_, _02135_);
  nor (_21058_, _21057_, _01653_);
  nand (_21060_, _21058_, _21056_);
  nand (_21061_, _21060_, _05060_);
  and (_21062_, _05040_, _04615_);
  nor (_21063_, _20892_, _05040_);
  or (_21064_, _21063_, _21062_);
  and (_21065_, _21064_, _05059_);
  nor (_21066_, _21065_, _05069_);
  and (_21067_, _21066_, _21061_);
  or (_21068_, _21067_, _20862_);
  nand (_21069_, _21068_, _05077_);
  and (_21071_, _04616_, _05072_);
  nor (_21072_, _21071_, _02039_);
  and (_21073_, _21072_, _21069_);
  or (_21074_, _21073_, _20860_);
  nand (_21075_, _21074_, _02131_);
  and (_21076_, _04615_, _02130_);
  nor (_21077_, _21076_, _01666_);
  nand (_21078_, _21077_, _21075_);
  nand (_21079_, _21078_, _05087_);
  and (_21080_, _20892_, _05092_);
  nor (_21082_, _04615_, _05092_);
  nor (_21083_, _21082_, _05087_);
  not (_21084_, _21083_);
  nor (_21085_, _21084_, _21080_);
  nor (_21086_, _21085_, _05097_);
  and (_21087_, _21086_, _21079_);
  or (_21088_, _21087_, _20859_);
  nand (_21089_, _21088_, _05105_);
  and (_21090_, _05101_, _04616_);
  nor (_21091_, _21090_, _02016_);
  and (_21093_, _21091_, _21089_);
  or (_21094_, _21093_, _20857_);
  nand (_21095_, _21094_, _05474_);
  and (_21096_, _04615_, _02126_);
  nor (_21097_, _21096_, _01663_);
  nand (_21098_, _21097_, _21095_);
  nand (_21099_, _21098_, _05115_);
  and (_21100_, _04615_, _05092_);
  nor (_21101_, _20892_, _05092_);
  or (_21102_, _21101_, _21100_);
  and (_21104_, _21102_, _05114_);
  nor (_21105_, _21104_, _05141_);
  and (_21106_, _21105_, _21099_);
  or (_21107_, _21106_, _20856_);
  nand (_21108_, _21107_, _05147_);
  and (_21109_, _04616_, _02273_);
  nor (_21110_, _21109_, _05145_);
  nand (_21111_, _21110_, _21108_);
  and (_21112_, _20854_, _05145_);
  nor (_21113_, _21112_, _02146_);
  nand (_21115_, _21113_, _21111_);
  nor (_21116_, _02015_, _01660_);
  not (_21117_, _21116_);
  and (_21118_, _03393_, _02146_);
  nor (_21119_, _21118_, _21117_);
  nand (_21120_, _21119_, _21115_);
  nor (_21121_, _05386_, _02983_);
  and (_21122_, _20906_, _05386_);
  or (_21123_, _21122_, _02153_);
  nor (_21124_, _21123_, _21121_);
  nor (_21126_, _21124_, _05161_);
  and (_21127_, _21126_, _21120_);
  or (_21128_, _21127_, _20855_);
  nand (_21129_, _21128_, _05398_);
  and (_21130_, _04616_, _02788_);
  nor (_21131_, _21130_, _05396_);
  nand (_21132_, _21131_, _21129_);
  and (_21133_, _20854_, _05396_);
  nor (_21134_, _21133_, _01585_);
  nand (_21135_, _21134_, _21132_);
  nor (_21137_, _02022_, _01581_);
  not (_21138_, _21137_);
  and (_21139_, _03393_, _01585_);
  nor (_21140_, _21139_, _21138_);
  nand (_21141_, _21140_, _21135_);
  and (_21142_, _05386_, _02983_);
  nor (_21143_, _20906_, _05386_);
  or (_21144_, _21143_, _21142_);
  and (_21145_, _21144_, _02022_);
  nor (_21146_, _21145_, _05419_);
  nand (_21148_, _21146_, _21141_);
  nor (_21149_, _20854_, _05418_);
  nor (_21150_, _21149_, _02164_);
  nand (_21151_, _21150_, _21148_);
  and (_21152_, _04615_, _02164_);
  nor (_21153_, _21152_, _05426_);
  nand (_21154_, _21153_, _21151_);
  and (_21155_, _20858_, _05426_);
  nor (_21156_, _21155_, _02023_);
  and (_21157_, _21156_, _21154_);
  or (_21159_, _21157_, _20847_);
  nand (_21160_, _21159_, _20821_);
  and (_21161_, _21144_, _02025_);
  nor (_21162_, _21161_, _05446_);
  nand (_21163_, _21162_, _21160_);
  nor (_21164_, _20854_, _05445_);
  nor (_21165_, _21164_, _01594_);
  nand (_21166_, _21165_, _21163_);
  and (_21167_, _04615_, _01594_);
  nor (_21168_, _21167_, _05453_);
  nand (_21170_, _21168_, _21166_);
  and (_21171_, _20858_, _05453_);
  nor (_21172_, _21171_, _02026_);
  and (_21173_, _21172_, _21170_);
  or (_21174_, _21173_, _20846_);
  nand (_21175_, _21174_, _20837_);
  and (_21176_, _20854_, _05464_);
  not (_21177_, _21176_);
  and (_21178_, _21177_, _21175_);
  nand (_21179_, _21178_, _26505_);
  or (_21181_, _26505_, \oc8051_golden_model_1.PC [9]);
  and (_21182_, _21181_, _25964_);
  and (_27925_, _21182_, _21179_);
  and (_21183_, _02833_, _20139_);
  nor (_21184_, _02795_, \oc8051_golden_model_1.PC [10]);
  nor (_21185_, _21184_, _21183_);
  and (_21186_, _21185_, _05464_);
  not (_21187_, _21186_);
  and (_21188_, _02263_, _02026_);
  nor (_21189_, _21185_, _05445_);
  and (_21191_, _02263_, _02023_);
  nor (_21192_, _21185_, _05418_);
  and (_21193_, _04600_, _02135_);
  and (_21194_, _21185_, _04960_);
  not (_21195_, _21185_);
  nor (_21196_, _21195_, _04905_);
  and (_21197_, _04874_, _02967_);
  not (_21198_, _02980_);
  nor (_21199_, _03150_, _03147_);
  nor (_21200_, _21199_, _21198_);
  and (_21202_, _21199_, _21198_);
  nor (_21203_, _21202_, _21200_);
  not (_21204_, _21203_);
  nor (_21205_, _21204_, _04874_);
  nor (_21206_, _21205_, _21197_);
  nor (_21207_, _21206_, _02378_);
  nor (_21208_, _21203_, _03909_);
  and (_21209_, _03909_, _02968_);
  nor (_21210_, _21209_, _21208_);
  and (_21211_, _21210_, _03185_);
  and (_21213_, _04601_, _01967_);
  or (_21214_, _04551_, _02968_);
  or (_21215_, _21204_, _04553_);
  and (_21216_, _21215_, _01969_);
  and (_21217_, _21216_, _21214_);
  and (_21218_, _04710_, _04600_);
  not (_21219_, _04612_);
  nor (_21220_, _04681_, _04678_);
  nor (_21221_, _21220_, _21219_);
  and (_21222_, _21220_, _21219_);
  nor (_21224_, _21222_, _21221_);
  and (_21225_, _21224_, _04707_);
  nor (_21226_, _21225_, _21218_);
  nand (_21227_, _21226_, _04557_);
  and (_21228_, _21185_, _04562_);
  and (_21229_, _21195_, _04563_);
  nor (_21230_, _21185_, _04561_);
  and (_21231_, _04571_, _04601_);
  or (_21232_, _04571_, \oc8051_golden_model_1.PC [10]);
  nor (_21233_, _21232_, _04560_);
  or (_21235_, _21233_, _21231_);
  and (_21236_, _21235_, _17901_);
  nor (_21237_, _21236_, _21230_);
  nor (_21238_, _21237_, _20875_);
  nor (_21239_, _21238_, _21229_);
  and (_21240_, _21239_, _02424_);
  and (_21241_, _04600_, _01971_);
  or (_21242_, _21241_, _21240_);
  and (_21243_, _21242_, _17894_);
  or (_21244_, _21243_, _20556_);
  nor (_21246_, _21244_, _21228_);
  nor (_21247_, _21246_, _04715_);
  nand (_21248_, _21247_, _21227_);
  and (_21249_, _21185_, _04715_);
  nor (_21250_, _21249_, _01969_);
  and (_21251_, _21250_, _21248_);
  or (_21252_, _21251_, _21217_);
  nand (_21253_, _21252_, _17940_);
  and (_21254_, _21195_, _04094_);
  nor (_21255_, _21254_, _01959_);
  nand (_21257_, _21255_, _21253_);
  and (_21258_, _04600_, _01959_);
  nor (_21259_, _21258_, _06363_);
  and (_21260_, _21259_, _05487_);
  and (_21261_, _21260_, _21257_);
  or (_21262_, _21261_, _21213_);
  or (_21263_, _21262_, _04725_);
  nand (_21264_, _21185_, _04725_);
  and (_21265_, _21264_, _01964_);
  nand (_21266_, _21265_, _21263_);
  and (_21268_, _04601_, _01963_);
  nor (_21269_, _21268_, _04734_);
  and (_21270_, _21269_, _21266_);
  and (_21271_, _21185_, _04734_);
  or (_21272_, _21271_, _21270_);
  nand (_21273_, _21272_, _06229_);
  and (_21274_, _21273_, _01630_);
  or (_21275_, _21274_, _01953_);
  or (_21276_, _04601_, _02455_);
  and (_21277_, _21276_, _04090_);
  nand (_21279_, _21277_, _21275_);
  and (_21280_, _04085_, _02967_);
  nor (_21281_, _21204_, _04085_);
  or (_21282_, _21281_, _04090_);
  nor (_21283_, _21282_, _21280_);
  nor (_21284_, _21283_, _03185_);
  and (_21285_, _21284_, _21279_);
  or (_21286_, _21285_, _21211_);
  and (_21287_, _21286_, _02378_);
  or (_21288_, _21287_, _21207_);
  nand (_21290_, _21288_, _04749_);
  nand (_21291_, _02967_, _02912_);
  nand (_21292_, _21203_, _19160_);
  and (_21293_, _21292_, _21291_);
  or (_21294_, _21293_, _04749_);
  and (_21295_, _21294_, _21290_);
  or (_21296_, _21295_, _02880_);
  nand (_21297_, _21185_, _02880_);
  and (_21298_, _21297_, _21296_);
  nor (_21299_, _21298_, _01946_);
  and (_21301_, _04600_, _01946_);
  nor (_21302_, _21301_, _21299_);
  nand (_21303_, _21302_, _04898_);
  nor (_21304_, _04897_, _04600_);
  nor (_21305_, _21304_, _04908_);
  and (_21306_, _21305_, _21303_);
  or (_21307_, _21306_, _21196_);
  nand (_21308_, _21307_, _01932_);
  nor (_21309_, _04601_, _01932_);
  nor (_21310_, _21309_, _17710_);
  and (_21312_, _21310_, _04928_);
  nand (_21313_, _21312_, _21308_);
  nor (_21314_, _21185_, _04928_);
  nor (_21315_, _21314_, _04932_);
  and (_21316_, _21315_, _21313_);
  and (_21317_, _04600_, _04932_);
  or (_21318_, _21317_, _01611_);
  or (_21319_, _21318_, _21316_);
  and (_21320_, _21195_, _01611_);
  nor (_21321_, _21320_, _01924_);
  nand (_21323_, _21321_, _21319_);
  and (_21324_, _04600_, _01924_);
  nor (_21325_, _21324_, _20657_);
  nand (_21326_, _21325_, _21323_);
  and (_21327_, _02968_, _02001_);
  nor (_21328_, _21327_, _04953_);
  nand (_21329_, _21328_, _21326_);
  nor (_21330_, _04952_, _04601_);
  nor (_21331_, _21330_, _01602_);
  and (_21332_, _21331_, _21329_);
  nor (_21334_, _04960_, _02968_);
  nor (_21335_, _21334_, _17728_);
  nor (_21336_, _21335_, _21332_);
  or (_21337_, _21336_, _21194_);
  nand (_21338_, _21337_, _02519_);
  and (_21339_, _04600_, _01920_);
  not (_21340_, _21339_);
  and (_21341_, _21340_, _20520_);
  nand (_21342_, _21341_, _21338_);
  nor (_21343_, _21224_, _04969_);
  nor (_21345_, _21343_, _02859_);
  and (_21346_, _21345_, _21342_);
  and (_21347_, _02859_, _04600_);
  or (_21348_, _21347_, _02019_);
  or (_21349_, _21348_, _21346_);
  and (_21350_, _02968_, _02019_);
  nor (_21351_, _21350_, _02853_);
  nand (_21352_, _21351_, _21349_);
  and (_21353_, _04600_, _02853_);
  nor (_21354_, _21353_, _04984_);
  nand (_21356_, _21354_, _21352_);
  nor (_21357_, _05012_, \oc8051_golden_model_1.DPH [2]);
  nor (_21358_, _21357_, _05013_);
  nor (_21359_, _21358_, _04985_);
  nor (_21360_, _21359_, _01919_);
  and (_21361_, _21360_, _21356_);
  and (_21362_, _04600_, _01919_);
  or (_21363_, _21362_, _21361_);
  nor (_21364_, _05026_, _01650_);
  nand (_21365_, _21364_, _21363_);
  nand (_21367_, _05038_, _04600_);
  nand (_21368_, _21224_, _05040_);
  and (_21369_, _21368_, _21367_);
  or (_21370_, _21369_, _05027_);
  nand (_21371_, _21370_, _21365_);
  and (_21372_, _21371_, _02830_);
  nor (_21373_, _21195_, _02830_);
  nor (_21374_, _21373_, _21372_);
  or (_21375_, _21374_, _05047_);
  nand (_21376_, _05047_, _04600_);
  and (_21378_, _21376_, _05049_);
  nand (_21379_, _21378_, _21375_);
  and (_21380_, _02968_, _02018_);
  nor (_21381_, _21380_, _02135_);
  and (_21382_, _21381_, _21379_);
  or (_21383_, _21382_, _21193_);
  nor (_21384_, _05059_, _01653_);
  nand (_21385_, _21384_, _21383_);
  nand (_21386_, _05040_, _04600_);
  nand (_21387_, _21224_, _05038_);
  and (_21389_, _21387_, _21386_);
  or (_21390_, _21389_, _05060_);
  nand (_21391_, _21390_, _21385_);
  and (_21392_, _21391_, _05070_);
  and (_21393_, _21185_, _05069_);
  nor (_21394_, _21393_, _21392_);
  or (_21395_, _21394_, _05072_);
  nand (_21396_, _04600_, _05072_);
  and (_21397_, _21396_, _05076_);
  nand (_21398_, _21397_, _21395_);
  and (_21400_, _02968_, _02039_);
  nor (_21401_, _21400_, _02130_);
  and (_21402_, _21401_, _21398_);
  and (_21403_, _04600_, _02130_);
  or (_21404_, _21403_, _21402_);
  nand (_21405_, _21404_, _20737_);
  nor (_21406_, _21224_, \oc8051_golden_model_1.PSW [7]);
  nor (_21407_, _04600_, _05092_);
  nor (_21408_, _21407_, _05087_);
  not (_21409_, _21408_);
  nor (_21411_, _21409_, _21406_);
  nor (_21412_, _21411_, _05097_);
  nand (_21413_, _21412_, _21405_);
  and (_21414_, _21195_, _05097_);
  nor (_21415_, _21414_, _05101_);
  and (_21416_, _21415_, _21413_);
  and (_21417_, _05101_, _04600_);
  or (_21418_, _21417_, _21416_);
  and (_21419_, _21418_, _05104_);
  and (_21420_, _02967_, _02016_);
  or (_21422_, _21420_, _02126_);
  or (_21423_, _21422_, _21419_);
  and (_21424_, _04601_, _02126_);
  nor (_21425_, _21424_, _20760_);
  nand (_21426_, _21425_, _21423_);
  and (_21427_, _04600_, _05092_);
  and (_21428_, _21224_, \oc8051_golden_model_1.PSW [7]);
  or (_21429_, _21428_, _21427_);
  and (_21430_, _21429_, _05114_);
  nor (_21431_, _21430_, _05141_);
  nand (_21433_, _21431_, _21426_);
  nor (_21434_, _21185_, _05139_);
  nor (_21435_, _21434_, _02273_);
  and (_21436_, _21435_, _21433_);
  and (_21437_, _04600_, _02273_);
  or (_21438_, _21437_, _21436_);
  and (_21439_, _21438_, _05146_);
  and (_21440_, _21185_, _05145_);
  or (_21441_, _21440_, _02146_);
  or (_21442_, _21441_, _21439_);
  and (_21444_, _03272_, _02146_);
  nor (_21445_, _21444_, _21117_);
  and (_21446_, _21445_, _21442_);
  or (_21447_, _05386_, _02967_);
  nand (_21448_, _21204_, _05386_);
  and (_21449_, _21448_, _02015_);
  and (_21450_, _21449_, _21447_);
  or (_21451_, _21450_, _05161_);
  nor (_21452_, _21451_, _21446_);
  nor (_21453_, _21185_, _02818_);
  or (_21455_, _21453_, _21452_);
  or (_21456_, _21455_, _02788_);
  nand (_21457_, _04600_, _02788_);
  and (_21458_, _21457_, _05397_);
  and (_21459_, _21458_, _21456_);
  and (_21460_, _21195_, _05396_);
  or (_21461_, _21460_, _21459_);
  nand (_21462_, _21461_, _01596_);
  and (_21463_, _03272_, _01585_);
  nor (_21464_, _21463_, _21138_);
  nand (_21466_, _21464_, _21462_);
  nor (_21467_, _21203_, _05386_);
  and (_21468_, _05386_, _02968_);
  nor (_21469_, _21468_, _21467_);
  and (_21470_, _21469_, _02022_);
  nor (_21471_, _21470_, _05419_);
  and (_21472_, _21471_, _21466_);
  or (_21473_, _21472_, _21192_);
  nand (_21474_, _21473_, _02168_);
  and (_21475_, _04601_, _02164_);
  nor (_21477_, _21475_, _05426_);
  nand (_21478_, _21477_, _21474_);
  and (_21479_, _21185_, _05426_);
  nor (_21480_, _21479_, _02023_);
  nand (_21481_, _21480_, _21478_);
  nand (_21482_, _21481_, _20821_);
  or (_21483_, _21482_, _21191_);
  and (_21484_, _21469_, _02025_);
  nor (_21485_, _21484_, _05446_);
  and (_21486_, _21485_, _21483_);
  or (_21488_, _21486_, _21189_);
  nand (_21489_, _21488_, _01595_);
  and (_21490_, _04601_, _01594_);
  nor (_21491_, _21490_, _05453_);
  nand (_21492_, _21491_, _21489_);
  and (_21493_, _21185_, _05453_);
  nor (_21494_, _21493_, _02026_);
  nand (_21495_, _21494_, _21492_);
  nand (_21496_, _21495_, _20837_);
  or (_21497_, _21496_, _21188_);
  and (_21499_, _21497_, _21187_);
  nand (_21500_, _21499_, _26505_);
  or (_21501_, _26505_, \oc8051_golden_model_1.PC [10]);
  and (_21502_, _21501_, _25964_);
  and (_27926_, _21502_, _21500_);
  and (_21503_, _03473_, _01585_);
  nor (_21504_, _21183_, _02971_);
  and (_21505_, _21183_, _02971_);
  or (_21506_, _21505_, _21504_);
  nor (_21507_, _21506_, _02818_);
  and (_21509_, _03473_, _02146_);
  and (_21510_, _04606_, _05092_);
  nor (_21511_, _21221_, _04602_);
  nor (_21512_, _21511_, _04610_);
  and (_21513_, _21511_, _04610_);
  or (_21514_, _21513_, _21512_);
  and (_21515_, _21514_, \oc8051_golden_model_1.PSW [7]);
  or (_21516_, _21515_, _21510_);
  and (_21517_, _21516_, _05114_);
  not (_21518_, _21506_);
  and (_21520_, _21518_, _05097_);
  and (_21521_, _05040_, _04606_);
  and (_21522_, _21514_, _05038_);
  or (_21523_, _21522_, _21521_);
  and (_21524_, _21523_, _05059_);
  nor (_21525_, _21506_, _02830_);
  and (_21526_, _02974_, _02912_);
  nor (_21527_, _21200_, _02969_);
  and (_21528_, _21527_, _02978_);
  nor (_21529_, _21527_, _02978_);
  nor (_21531_, _21529_, _21528_);
  nor (_21532_, _21531_, _02912_);
  or (_21533_, _21532_, _21526_);
  and (_21534_, _21533_, _03179_);
  and (_21535_, _03909_, _02974_);
  nor (_21536_, _21531_, _03909_);
  or (_21537_, _21536_, _21535_);
  nor (_21538_, _21537_, _03187_);
  and (_21539_, _04085_, _02974_);
  nor (_21540_, _21531_, _04085_);
  or (_21542_, _21540_, _21539_);
  nor (_21543_, _21542_, _04090_);
  and (_21544_, _04606_, _01963_);
  not (_21545_, _21531_);
  and (_21546_, _21545_, _04551_);
  and (_21547_, _04553_, _02974_);
  or (_21548_, _21547_, _02438_);
  or (_21549_, _21548_, _21546_);
  nor (_21550_, _04607_, _01627_);
  nor (_21551_, _21506_, _18336_);
  not (_21553_, _21551_);
  and (_21554_, _04571_, _04607_);
  nor (_21555_, _04571_, \oc8051_golden_model_1.PC [11]);
  and (_21556_, _21555_, _18340_);
  nor (_21557_, _21556_, _21554_);
  nor (_21558_, _21557_, _18347_);
  nor (_21559_, _04606_, _01625_);
  nor (_21560_, _21559_, _01971_);
  not (_21561_, _21560_);
  nor (_21562_, _21561_, _21558_);
  and (_21564_, _21562_, _21553_);
  and (_21565_, _04606_, _01971_);
  or (_21566_, _21565_, _21564_);
  and (_21567_, _21566_, _17894_);
  and (_21568_, _21506_, _04562_);
  or (_21569_, _21568_, _21567_);
  and (_21570_, _21569_, _01627_);
  or (_21571_, _21570_, _04557_);
  nor (_21572_, _21571_, _21550_);
  and (_21573_, _04710_, _04606_);
  and (_21575_, _21514_, _04707_);
  or (_21576_, _21575_, _04709_);
  nor (_21577_, _21576_, _21573_);
  nor (_21578_, _21577_, _21572_);
  or (_21579_, _21578_, _04716_);
  and (_21580_, _21579_, _21549_);
  or (_21581_, _21580_, _04094_);
  or (_21582_, _21506_, _04721_);
  and (_21583_, _21582_, _04720_);
  and (_21584_, _21583_, _21581_);
  nor (_21586_, _04720_, _04607_);
  or (_21587_, _21586_, _04725_);
  nor (_21588_, _21587_, _21584_);
  and (_21589_, _21518_, _04725_);
  nor (_21590_, _21589_, _01963_);
  not (_21591_, _21590_);
  nor (_21592_, _21591_, _21588_);
  nor (_21593_, _21592_, _21544_);
  nor (_21594_, _21593_, _04734_);
  and (_21595_, _21506_, _04734_);
  nor (_21597_, _21595_, _04739_);
  not (_21598_, _21597_);
  nor (_21599_, _21598_, _21594_);
  nor (_21600_, _04738_, _04606_);
  nor (_21601_, _21600_, _21599_);
  nor (_21602_, _21601_, _04089_);
  nor (_21603_, _21602_, _21543_);
  nor (_21604_, _21603_, _03185_);
  nor (_21605_, _21604_, _21538_);
  and (_21606_, _21605_, _02378_);
  nor (_21608_, _21531_, _04874_);
  and (_21609_, _04874_, _02974_);
  or (_21610_, _21609_, _21608_);
  and (_21611_, _21610_, _01951_);
  or (_21612_, _21611_, _21606_);
  and (_21613_, _21612_, _04749_);
  nor (_21614_, _21613_, _21534_);
  nor (_21615_, _21614_, _02880_);
  and (_21616_, _21506_, _02880_);
  not (_21617_, _21616_);
  and (_21619_, _21617_, _04899_);
  not (_21620_, _21619_);
  nor (_21621_, _21620_, _21615_);
  nor (_21622_, _04899_, _04606_);
  nor (_21623_, _21622_, _04908_);
  not (_21624_, _21623_);
  nor (_21625_, _21624_, _21621_);
  nor (_21626_, _21518_, _04905_);
  or (_21627_, _21626_, _04911_);
  or (_21628_, _21627_, _21625_);
  or (_21630_, _04910_, _04606_);
  and (_21631_, _21630_, _04928_);
  and (_21632_, _21631_, _21628_);
  nor (_21633_, _21518_, _04928_);
  nor (_21634_, _21633_, _04932_);
  not (_21635_, _21634_);
  nor (_21636_, _21635_, _21632_);
  and (_21637_, _04607_, _04932_);
  nor (_21638_, _21637_, _01611_);
  not (_21639_, _21638_);
  nor (_21641_, _21639_, _21636_);
  and (_21642_, _21506_, _01611_);
  nor (_21643_, _21642_, _04943_);
  not (_21644_, _21643_);
  nor (_21645_, _21644_, _21641_);
  nor (_21646_, _04942_, _04606_);
  nor (_21647_, _21646_, _02001_);
  not (_21648_, _21647_);
  nor (_21649_, _21648_, _21645_);
  and (_21650_, _02974_, _02001_);
  nor (_21652_, _21650_, _04953_);
  not (_21653_, _21652_);
  or (_21654_, _21653_, _21649_);
  nor (_21655_, _04952_, _04606_);
  nor (_21656_, _21655_, _01602_);
  and (_21657_, _21656_, _21654_);
  nor (_21658_, _04960_, _02974_);
  nor (_21659_, _21658_, _17728_);
  nor (_21660_, _21659_, _21657_);
  and (_21661_, _21518_, _04960_);
  or (_21663_, _21661_, _21660_);
  nand (_21664_, _21663_, _04963_);
  nor (_21665_, _04963_, _04606_);
  nor (_21666_, _21665_, _04968_);
  nand (_21667_, _21666_, _21664_);
  and (_21668_, _21514_, _04968_);
  nor (_21669_, _21668_, _02859_);
  nand (_21670_, _21669_, _21667_);
  and (_21671_, _02859_, _04607_);
  nor (_21672_, _21671_, _02019_);
  nand (_21674_, _21672_, _21670_);
  and (_21675_, _02974_, _02019_);
  nor (_21676_, _21675_, _02853_);
  nand (_21677_, _21676_, _21674_);
  and (_21678_, _04607_, _02853_);
  nor (_21679_, _21678_, _04984_);
  nand (_21680_, _21679_, _21677_);
  nor (_21681_, _05013_, \oc8051_golden_model_1.DPH [3]);
  or (_21682_, _21681_, _04985_);
  or (_21683_, _21682_, _05014_);
  and (_21685_, _21683_, _05022_);
  nand (_21686_, _21685_, _21680_);
  nor (_21687_, _05022_, _04606_);
  nor (_21688_, _21687_, _05026_);
  nand (_21689_, _21688_, _21686_);
  and (_21690_, _05038_, _04606_);
  and (_21691_, _21514_, _05040_);
  or (_21692_, _21691_, _21690_);
  and (_21693_, _21692_, _05026_);
  nor (_21694_, _21693_, _05031_);
  and (_21696_, _21694_, _21689_);
  or (_21697_, _21696_, _21525_);
  nand (_21698_, _21697_, _05050_);
  and (_21699_, _05047_, _04607_);
  nor (_21700_, _21699_, _02018_);
  nand (_21701_, _21700_, _21698_);
  and (_21702_, _02974_, _02018_);
  nor (_21703_, _21702_, _05056_);
  nand (_21704_, _21703_, _21701_);
  nor (_21705_, _05055_, _04606_);
  nor (_21707_, _21705_, _05059_);
  and (_21708_, _21707_, _21704_);
  or (_21709_, _21708_, _21524_);
  nand (_21710_, _21709_, _05070_);
  and (_21711_, _21506_, _05069_);
  nor (_21712_, _21711_, _05072_);
  nand (_21713_, _21712_, _21710_);
  and (_21714_, _04607_, _05072_);
  nor (_21715_, _21714_, _02039_);
  nand (_21716_, _21715_, _21713_);
  and (_21718_, _02974_, _02039_);
  nor (_21719_, _21718_, _05083_);
  nand (_21720_, _21719_, _21716_);
  nor (_21721_, _05082_, _04606_);
  nor (_21722_, _21721_, _05086_);
  nand (_21723_, _21722_, _21720_);
  nor (_21724_, _21514_, \oc8051_golden_model_1.PSW [7]);
  nor (_21725_, _04606_, _05092_);
  nor (_21726_, _21725_, _05087_);
  not (_21727_, _21726_);
  nor (_21729_, _21727_, _21724_);
  nor (_21730_, _21729_, _05097_);
  and (_21731_, _21730_, _21723_);
  or (_21732_, _21731_, _21520_);
  nand (_21733_, _21732_, _05105_);
  and (_21734_, _05101_, _04607_);
  nor (_21735_, _21734_, _02016_);
  nand (_21736_, _21735_, _21733_);
  and (_21737_, _02974_, _02016_);
  nor (_21738_, _21737_, _05111_);
  nand (_21740_, _21738_, _21736_);
  nor (_21741_, _05110_, _04606_);
  nor (_21742_, _21741_, _05114_);
  and (_21743_, _21742_, _21740_);
  or (_21744_, _21743_, _21517_);
  nand (_21745_, _21744_, _05139_);
  nor (_21746_, _21518_, _05139_);
  nor (_21747_, _21746_, _02273_);
  nand (_21748_, _21747_, _21745_);
  and (_21749_, _04607_, _02273_);
  nor (_21751_, _21749_, _05145_);
  nand (_21752_, _21751_, _21748_);
  and (_21753_, _21506_, _05145_);
  nor (_21754_, _21753_, _02146_);
  and (_21755_, _21754_, _21752_);
  or (_21756_, _21755_, _21509_);
  nand (_21757_, _21756_, _05157_);
  and (_21758_, _04607_, _01660_);
  nor (_21759_, _21758_, _02015_);
  nand (_21760_, _21759_, _21757_);
  nor (_21762_, _05386_, _02974_);
  and (_21763_, _21531_, _05386_);
  or (_21764_, _21763_, _02153_);
  nor (_21765_, _21764_, _21762_);
  nor (_21766_, _21765_, _05161_);
  and (_21767_, _21766_, _21760_);
  or (_21768_, _21767_, _21507_);
  nand (_21769_, _21768_, _05398_);
  and (_21770_, _04607_, _02788_);
  nor (_21771_, _21770_, _05396_);
  nand (_21773_, _21771_, _21769_);
  and (_21774_, _21506_, _05396_);
  nor (_21775_, _21774_, _01585_);
  and (_21776_, _21775_, _21773_);
  or (_21777_, _21776_, _21503_);
  nand (_21778_, _21777_, _05407_);
  and (_21779_, _04607_, _01581_);
  nor (_21780_, _21779_, _02022_);
  nand (_21781_, _21780_, _21778_);
  nor (_21782_, _21545_, _05386_);
  and (_21784_, _05386_, _02975_);
  nor (_21785_, _21784_, _21782_);
  and (_21786_, _21785_, _02022_);
  nor (_21787_, _21786_, _05419_);
  nand (_21788_, _21787_, _21781_);
  nor (_21789_, _21506_, _05418_);
  nor (_21790_, _21789_, _02164_);
  nand (_21791_, _21790_, _21788_);
  and (_21792_, _04606_, _02164_);
  nor (_21793_, _21792_, _05426_);
  nand (_21795_, _21793_, _21791_);
  and (_21796_, _21518_, _05426_);
  nor (_21797_, _21796_, _02023_);
  nand (_21798_, _21797_, _21795_);
  and (_21799_, _02023_, _01916_);
  nor (_21800_, _21799_, _01670_);
  nand (_21801_, _21800_, _21798_);
  and (_21802_, _04607_, _01670_);
  nor (_21803_, _21802_, _02025_);
  nand (_21804_, _21803_, _21801_);
  and (_21806_, _21785_, _02025_);
  nor (_21807_, _21806_, _05446_);
  nand (_21808_, _21807_, _21804_);
  nor (_21809_, _21506_, _05445_);
  nor (_21810_, _21809_, _01594_);
  nand (_21811_, _21810_, _21808_);
  and (_21812_, _04606_, _01594_);
  nor (_21813_, _21812_, _05453_);
  nand (_21814_, _21813_, _21811_);
  and (_21815_, _21518_, _05453_);
  nor (_21817_, _21815_, _02026_);
  nand (_21818_, _21817_, _21814_);
  and (_21819_, _02026_, _01916_);
  nor (_21820_, _21819_, _01657_);
  and (_21821_, _21820_, _21818_);
  and (_21822_, _04607_, _01657_);
  nor (_21823_, _21822_, _21821_);
  nand (_21824_, _21823_, _05465_);
  and (_21825_, _21506_, _05464_);
  not (_21826_, _21825_);
  and (_21828_, _21826_, _21824_);
  nand (_21829_, _21828_, _26505_);
  or (_21830_, _26505_, \oc8051_golden_model_1.PC [11]);
  and (_21831_, _21830_, _25964_);
  and (_27927_, _21831_, _21829_);
  and (_21832_, _21183_, \oc8051_golden_model_1.PC [11]);
  nor (_21833_, _21832_, \oc8051_golden_model_1.PC [12]);
  nor (_21834_, _21833_, _02798_);
  or (_21835_, _21834_, _05445_);
  nand (_21836_, _04024_, _02146_);
  nor (_21838_, _04688_, _04686_);
  nor (_21839_, _21838_, _04689_);
  or (_21840_, _21839_, _05092_);
  or (_21841_, _04596_, \oc8051_golden_model_1.PSW [7]);
  and (_21842_, _21841_, _05114_);
  and (_21843_, _21842_, _21840_);
  and (_21844_, _02964_, _01602_);
  and (_21845_, _03909_, _02964_);
  not (_21846_, _03909_);
  nor (_21847_, _03158_, _03156_);
  nor (_21849_, _21847_, _03159_);
  and (_21850_, _21849_, _21846_);
  or (_21851_, _21850_, _21845_);
  or (_21852_, _21851_, _03187_);
  and (_21853_, _04085_, _02964_);
  not (_21854_, _04085_);
  and (_21855_, _21849_, _21854_);
  or (_21856_, _21855_, _21853_);
  or (_21857_, _21856_, _04090_);
  not (_21858_, _04720_);
  or (_21860_, _21834_, _04721_);
  or (_21861_, _21849_, _04553_);
  or (_21862_, _04551_, _02964_);
  and (_21863_, _21862_, _21861_);
  or (_21864_, _21863_, _02438_);
  and (_21865_, _21834_, _04559_);
  and (_21866_, _04561_, \oc8051_golden_model_1.PC [12]);
  and (_21867_, _21834_, _04560_);
  or (_21868_, _21867_, _21866_);
  and (_21869_, _21868_, _05488_);
  or (_21871_, _21869_, _21865_);
  and (_21872_, _21871_, _01625_);
  and (_21873_, _04578_, _04596_);
  or (_21874_, _21873_, _21872_);
  and (_21875_, _21874_, _18334_);
  and (_21876_, _21834_, _04563_);
  or (_21877_, _21876_, _01971_);
  or (_21878_, _21877_, _21875_);
  nand (_21879_, _04597_, _01971_);
  and (_21880_, _21879_, _21878_);
  or (_21882_, _21880_, _04562_);
  or (_21883_, _21834_, _17894_);
  and (_21884_, _21883_, _01627_);
  and (_21885_, _21884_, _21882_);
  nor (_21886_, _04597_, _01627_);
  or (_21887_, _21886_, _04557_);
  or (_21888_, _21887_, _21885_);
  and (_21889_, _04710_, _04596_);
  and (_21890_, _21839_, _04707_);
  or (_21891_, _21890_, _04709_);
  or (_21893_, _21891_, _21889_);
  and (_21894_, _21893_, _21888_);
  or (_21895_, _21894_, _04716_);
  and (_21896_, _21895_, _21864_);
  or (_21897_, _21896_, _04094_);
  and (_21898_, _21897_, _21860_);
  or (_21899_, _21898_, _21858_);
  or (_21900_, _04720_, _04596_);
  and (_21901_, _21900_, _04729_);
  and (_21902_, _21901_, _21899_);
  and (_21904_, _21834_, _04725_);
  or (_21905_, _21904_, _01963_);
  or (_21906_, _21905_, _21902_);
  and (_21907_, _04597_, _01963_);
  nor (_21908_, _21907_, _04734_);
  and (_21909_, _21908_, _21906_);
  nand (_21910_, _21834_, _04734_);
  nand (_21911_, _21910_, _04738_);
  or (_21912_, _21911_, _21909_);
  or (_21913_, _04738_, _04596_);
  and (_21915_, _21913_, _21912_);
  or (_21916_, _21915_, _04089_);
  and (_21917_, _21916_, _21857_);
  or (_21918_, _21917_, _03185_);
  and (_21919_, _21918_, _21852_);
  or (_21920_, _21919_, _01951_);
  and (_21921_, _04874_, _02964_);
  and (_21922_, _21849_, _04875_);
  or (_21923_, _21922_, _02378_);
  or (_21924_, _21923_, _21921_);
  and (_21926_, _21924_, _04749_);
  and (_21927_, _21926_, _21920_);
  or (_21928_, _21849_, _02912_);
  or (_21929_, _02964_, _19160_);
  and (_21930_, _21929_, _03179_);
  and (_21931_, _21930_, _21928_);
  or (_21932_, _21931_, _21927_);
  and (_21933_, _21932_, _02881_);
  nand (_21934_, _21834_, _02880_);
  nand (_21935_, _21934_, _04899_);
  or (_21937_, _21935_, _21933_);
  or (_21938_, _04899_, _04596_);
  and (_21939_, _21938_, _04905_);
  and (_21940_, _21939_, _21937_);
  and (_21941_, _21834_, _04908_);
  or (_21942_, _21941_, _04911_);
  or (_21943_, _21942_, _21940_);
  or (_21944_, _04910_, _04596_);
  and (_21945_, _21944_, _04928_);
  and (_21946_, _21945_, _21943_);
  and (_21948_, _21834_, _04933_);
  or (_21949_, _21948_, _04932_);
  or (_21950_, _21949_, _21946_);
  nand (_21951_, _04597_, _04932_);
  and (_21952_, _21951_, _01616_);
  and (_21953_, _21952_, _21950_);
  nand (_21954_, _21834_, _01611_);
  nand (_21955_, _21954_, _04942_);
  or (_21956_, _21955_, _21953_);
  or (_21957_, _04942_, _04596_);
  and (_21959_, _21957_, _02002_);
  and (_21960_, _21959_, _21956_);
  nand (_21961_, _02964_, _02001_);
  nand (_21962_, _21961_, _04952_);
  or (_21963_, _21962_, _21960_);
  or (_21964_, _04952_, _04596_);
  and (_21965_, _21964_, _01923_);
  and (_21966_, _21965_, _21963_);
  or (_21967_, _21966_, _21844_);
  and (_21968_, _21967_, _04961_);
  and (_21970_, _21834_, _04960_);
  or (_21971_, _21970_, _04964_);
  or (_21972_, _21971_, _21968_);
  or (_21973_, _04963_, _04596_);
  and (_21974_, _21973_, _04969_);
  and (_21975_, _21974_, _21972_);
  and (_21976_, _21839_, _04968_);
  or (_21977_, _21976_, _02859_);
  or (_21978_, _21977_, _21975_);
  nor (_21979_, _04597_, _02019_);
  or (_21981_, _21979_, _07508_);
  and (_21982_, _21981_, _21978_);
  and (_21983_, _02964_, _02019_);
  or (_21984_, _21983_, _02853_);
  or (_21985_, _21984_, _21982_);
  nand (_21986_, _04597_, _02853_);
  and (_21987_, _21986_, _04985_);
  and (_21988_, _21987_, _21985_);
  nor (_21989_, _05014_, \oc8051_golden_model_1.DPH [4]);
  nor (_21990_, _21989_, _05015_);
  and (_21992_, _21990_, _04984_);
  or (_21993_, _21992_, _05023_);
  or (_21994_, _21993_, _21988_);
  or (_21995_, _05022_, _04596_);
  and (_21996_, _21995_, _05027_);
  and (_21997_, _21996_, _21994_);
  or (_21998_, _21839_, _05038_);
  or (_21999_, _05040_, _04596_);
  and (_22000_, _21999_, _05026_);
  and (_22001_, _22000_, _21998_);
  or (_22003_, _22001_, _21997_);
  and (_22004_, _22003_, _02830_);
  and (_22005_, _21834_, _05031_);
  or (_22006_, _22005_, _05047_);
  or (_22007_, _22006_, _22004_);
  nand (_22008_, _05047_, _04597_);
  and (_22009_, _22008_, _05049_);
  and (_22010_, _22009_, _22007_);
  nand (_22011_, _02964_, _02018_);
  nand (_22012_, _22011_, _05055_);
  or (_22014_, _22012_, _22010_);
  or (_22015_, _05055_, _04596_);
  and (_22016_, _22015_, _05060_);
  and (_22017_, _22016_, _22014_);
  or (_22018_, _21839_, _05040_);
  or (_22019_, _05038_, _04596_);
  and (_22020_, _22019_, _05059_);
  and (_22021_, _22020_, _22018_);
  or (_22022_, _22021_, _22017_);
  and (_22023_, _22022_, _05070_);
  and (_22025_, _21834_, _05069_);
  or (_22026_, _22025_, _05072_);
  or (_22027_, _22026_, _22023_);
  nand (_22028_, _04597_, _05072_);
  and (_22029_, _22028_, _05076_);
  and (_22030_, _22029_, _22027_);
  nand (_22031_, _02964_, _02039_);
  nand (_22032_, _22031_, _05082_);
  or (_22033_, _22032_, _22030_);
  or (_22034_, _05082_, _04596_);
  and (_22036_, _22034_, _05087_);
  and (_22037_, _22036_, _22033_);
  or (_22038_, _21839_, \oc8051_golden_model_1.PSW [7]);
  or (_22039_, _04596_, _05092_);
  and (_22040_, _22039_, _05086_);
  and (_22041_, _22040_, _22038_);
  or (_22042_, _22041_, _22037_);
  and (_22043_, _22042_, _05098_);
  and (_22044_, _21834_, _05097_);
  or (_22045_, _22044_, _05101_);
  or (_22047_, _22045_, _22043_);
  nand (_22048_, _05101_, _04597_);
  and (_22049_, _22048_, _05104_);
  and (_22050_, _22049_, _22047_);
  nand (_22051_, _02964_, _02016_);
  nand (_22052_, _22051_, _05110_);
  or (_22053_, _22052_, _22050_);
  or (_22054_, _05110_, _04596_);
  and (_22055_, _22054_, _05115_);
  and (_22056_, _22055_, _22053_);
  or (_22058_, _22056_, _21843_);
  and (_22059_, _22058_, _05139_);
  and (_22060_, _21834_, _05141_);
  or (_22061_, _22060_, _02273_);
  or (_22062_, _22061_, _22059_);
  nand (_22063_, _04597_, _02273_);
  and (_22064_, _22063_, _05146_);
  and (_22065_, _22064_, _22062_);
  and (_22066_, _21834_, _05145_);
  or (_22067_, _22066_, _02146_);
  or (_22069_, _22067_, _22065_);
  and (_22070_, _22069_, _21836_);
  or (_22071_, _22070_, _01660_);
  nand (_22072_, _04597_, _01660_);
  and (_22073_, _22072_, _02153_);
  and (_22074_, _22073_, _22071_);
  or (_22075_, _21849_, _05387_);
  or (_22076_, _05386_, _02964_);
  and (_22077_, _22076_, _02015_);
  and (_22078_, _22077_, _22075_);
  or (_22080_, _22078_, _22074_);
  and (_22081_, _22080_, _02818_);
  and (_22082_, _21834_, _05161_);
  or (_22083_, _22082_, _02788_);
  or (_22084_, _22083_, _22081_);
  nand (_22085_, _04597_, _02788_);
  and (_22086_, _22085_, _05397_);
  and (_22087_, _22086_, _22084_);
  and (_22088_, _21834_, _05396_);
  or (_22089_, _22088_, _01585_);
  or (_22091_, _22089_, _22087_);
  nand (_22092_, _04024_, _01585_);
  and (_22093_, _22092_, _05407_);
  and (_22094_, _22093_, _22091_);
  and (_22095_, _04596_, _01581_);
  or (_22096_, _22095_, _02022_);
  or (_22097_, _22096_, _22094_);
  or (_22098_, _05387_, _02964_);
  or (_22099_, _21849_, _05386_);
  and (_22100_, _22099_, _22098_);
  or (_22102_, _22100_, _02558_);
  and (_22103_, _22102_, _05418_);
  and (_22104_, _22103_, _22097_);
  and (_22105_, _21834_, _05419_);
  or (_22106_, _22105_, _02164_);
  or (_22107_, _22106_, _22104_);
  nand (_22108_, _04597_, _02164_);
  and (_22109_, _22108_, _22107_);
  or (_22110_, _22109_, _05426_);
  or (_22111_, _21834_, _05430_);
  and (_22113_, _22111_, _22110_);
  or (_22114_, _22113_, _02023_);
  nand (_22115_, _02606_, _02023_);
  and (_22116_, _22115_, _01671_);
  and (_22117_, _22116_, _22114_);
  and (_22118_, _04596_, _01670_);
  or (_22119_, _22118_, _02025_);
  or (_22120_, _22119_, _22117_);
  or (_22121_, _22100_, _02377_);
  and (_22122_, _22121_, _22120_);
  or (_22124_, _22122_, _05446_);
  and (_22125_, _22124_, _21835_);
  or (_22126_, _22125_, _01594_);
  and (_22127_, _04597_, _01594_);
  nor (_22128_, _22127_, _05453_);
  and (_22129_, _22128_, _22126_);
  and (_22130_, _21834_, _05453_);
  or (_22131_, _22130_, _02026_);
  or (_22132_, _22131_, _22129_);
  nand (_22133_, _02606_, _02026_);
  and (_22135_, _22133_, _22132_);
  or (_22136_, _22135_, _01657_);
  nand (_22137_, _04597_, _01657_);
  and (_22138_, _22137_, _05465_);
  and (_22139_, _22138_, _22136_);
  and (_22140_, _21834_, _05464_);
  or (_22141_, _22140_, _22139_);
  or (_22142_, _22141_, _26506_);
  or (_22143_, _26505_, \oc8051_golden_model_1.PC [12]);
  and (_22144_, _22143_, _25964_);
  and (_27928_, _22144_, _22142_);
  nor (_22146_, _02798_, \oc8051_golden_model_1.PC [13]);
  nor (_22147_, _22146_, _02799_);
  and (_22148_, _22147_, _05464_);
  nand (_22149_, _03976_, _01585_);
  or (_22150_, _22147_, _02818_);
  nand (_22151_, _03976_, _02146_);
  or (_22152_, _22147_, _05098_);
  or (_22153_, _22147_, _05070_);
  or (_22154_, _22147_, _02830_);
  or (_22156_, _02961_, _02960_);
  nand (_22157_, _22156_, _03161_);
  or (_22158_, _22156_, _03161_);
  and (_22159_, _22158_, _22157_);
  or (_22160_, _22159_, _03909_);
  nand (_22161_, _03909_, _02959_);
  and (_22162_, _22161_, _22160_);
  or (_22163_, _22162_, _03187_);
  or (_22164_, _22159_, _04085_);
  nand (_22165_, _04085_, _02959_);
  and (_22167_, _22165_, _22164_);
  or (_22168_, _22167_, _04090_);
  and (_22169_, _04592_, _01963_);
  and (_22170_, _22159_, _04551_);
  and (_22171_, _04553_, _02958_);
  or (_22172_, _22171_, _02438_);
  or (_22173_, _22172_, _22170_);
  or (_22174_, _22147_, _18336_);
  nor (_22175_, _04571_, \oc8051_golden_model_1.PC [13]);
  nand (_22176_, _22175_, _18345_);
  or (_22178_, _22176_, _04560_);
  and (_22179_, _22178_, _22174_);
  or (_22180_, _22179_, _01971_);
  or (_22181_, _04579_, _04592_);
  and (_22182_, _22181_, _22180_);
  or (_22183_, _22182_, _04562_);
  or (_22184_, _22147_, _17894_);
  and (_22185_, _22184_, _01627_);
  and (_22186_, _22185_, _22183_);
  and (_22187_, _04592_, _04558_);
  or (_22189_, _22187_, _04557_);
  or (_22190_, _22189_, _22186_);
  or (_22191_, _04594_, _04593_);
  nand (_22192_, _22191_, _04690_);
  or (_22193_, _22191_, _04690_);
  and (_22194_, _22193_, _22192_);
  and (_22195_, _22194_, _04707_);
  and (_22196_, _04710_, _04592_);
  or (_22197_, _22196_, _04709_);
  or (_22198_, _22197_, _22195_);
  and (_22200_, _22198_, _22190_);
  or (_22201_, _22200_, _04716_);
  and (_22202_, _22201_, _22173_);
  or (_22203_, _22202_, _04094_);
  or (_22204_, _22147_, _04721_);
  and (_22205_, _22204_, _04720_);
  and (_22206_, _22205_, _22203_);
  and (_22207_, _21858_, _04592_);
  or (_22208_, _22207_, _04725_);
  or (_22209_, _22208_, _22206_);
  or (_22211_, _22147_, _04729_);
  and (_22212_, _22211_, _01964_);
  and (_22213_, _22212_, _22209_);
  or (_22214_, _22213_, _22169_);
  and (_22215_, _22214_, _04735_);
  nand (_22216_, _22147_, _04734_);
  nand (_22217_, _22216_, _04738_);
  or (_22218_, _22217_, _22215_);
  or (_22219_, _04738_, _04592_);
  and (_22220_, _22219_, _22218_);
  or (_22222_, _22220_, _04089_);
  and (_22223_, _22222_, _22168_);
  or (_22224_, _22223_, _03185_);
  and (_22225_, _22224_, _22163_);
  or (_22226_, _22225_, _01951_);
  and (_22227_, _22159_, _04875_);
  and (_22228_, _04874_, _02958_);
  or (_22229_, _22228_, _02378_);
  or (_22230_, _22229_, _22227_);
  and (_22231_, _22230_, _04749_);
  and (_22233_, _22231_, _22226_);
  or (_22234_, _22159_, _02912_);
  nand (_22235_, _02959_, _02912_);
  and (_22236_, _22235_, _03179_);
  and (_22237_, _22236_, _22234_);
  or (_22238_, _22237_, _22233_);
  and (_22239_, _22238_, _02881_);
  nand (_22240_, _22147_, _02880_);
  nand (_22241_, _22240_, _04899_);
  or (_22242_, _22241_, _22239_);
  or (_22244_, _04899_, _04592_);
  and (_22245_, _22244_, _04905_);
  and (_22246_, _22245_, _22242_);
  and (_22247_, _22147_, _04908_);
  or (_22248_, _22247_, _04911_);
  or (_22249_, _22248_, _22246_);
  or (_22250_, _04910_, _04592_);
  and (_22251_, _22250_, _04928_);
  and (_22252_, _22251_, _22249_);
  and (_22253_, _22147_, _04933_);
  or (_22255_, _22253_, _04932_);
  or (_22256_, _22255_, _22252_);
  or (_22257_, _04592_, _04937_);
  and (_22258_, _22257_, _01616_);
  and (_22259_, _22258_, _22256_);
  and (_22260_, _22147_, _01611_);
  or (_22261_, _22260_, _04943_);
  or (_22262_, _22261_, _22259_);
  or (_22263_, _04942_, _04592_);
  and (_22264_, _22263_, _02002_);
  and (_22266_, _22264_, _22262_);
  nand (_22267_, _02958_, _02001_);
  nand (_22268_, _22267_, _04952_);
  or (_22269_, _22268_, _22266_);
  or (_22270_, _04952_, _04592_);
  and (_22271_, _22270_, _01923_);
  and (_22272_, _22271_, _22269_);
  nor (_22273_, _04960_, _02958_);
  nor (_22274_, _22273_, _17728_);
  or (_22275_, _22274_, _22272_);
  or (_22277_, _22147_, _04961_);
  and (_22278_, _22277_, _22275_);
  or (_22279_, _22278_, _04964_);
  or (_22280_, _04963_, _04592_);
  and (_22281_, _22280_, _04969_);
  and (_22282_, _22281_, _22279_);
  and (_22283_, _22194_, _04968_);
  or (_22284_, _22283_, _02859_);
  or (_22285_, _22284_, _22282_);
  and (_22286_, _04592_, _04979_);
  or (_22288_, _22286_, _07508_);
  and (_22289_, _22288_, _22285_);
  and (_22290_, _02958_, _02019_);
  or (_22291_, _22290_, _02853_);
  or (_22292_, _22291_, _22289_);
  or (_22293_, _04592_, _04978_);
  and (_22294_, _22293_, _04985_);
  and (_22295_, _22294_, _22292_);
  or (_22296_, _05015_, \oc8051_golden_model_1.DPH [5]);
  nor (_22297_, _05016_, _04985_);
  and (_22299_, _22297_, _22296_);
  or (_22300_, _22299_, _05023_);
  or (_22301_, _22300_, _22295_);
  or (_22302_, _05022_, _04592_);
  and (_22303_, _22302_, _05027_);
  and (_22304_, _22303_, _22301_);
  or (_22305_, _22194_, _05038_);
  or (_22306_, _05040_, _04592_);
  and (_22307_, _22306_, _05026_);
  and (_22308_, _22307_, _22305_);
  or (_22310_, _22308_, _05031_);
  or (_22311_, _22310_, _22304_);
  and (_22312_, _22311_, _22154_);
  or (_22313_, _22312_, _05047_);
  or (_22314_, _05050_, _04592_);
  and (_22315_, _22314_, _05049_);
  and (_22316_, _22315_, _22313_);
  nand (_22317_, _02958_, _02018_);
  nand (_22318_, _22317_, _05055_);
  or (_22319_, _22318_, _22316_);
  or (_22321_, _05055_, _04592_);
  and (_22322_, _22321_, _05060_);
  and (_22323_, _22322_, _22319_);
  or (_22324_, _22194_, _05040_);
  or (_22325_, _05038_, _04592_);
  and (_22326_, _22325_, _05059_);
  and (_22327_, _22326_, _22324_);
  or (_22328_, _22327_, _05069_);
  or (_22329_, _22328_, _22323_);
  and (_22330_, _22329_, _22153_);
  or (_22332_, _22330_, _05072_);
  or (_22333_, _04592_, _05077_);
  and (_22334_, _22333_, _05076_);
  and (_22335_, _22334_, _22332_);
  nand (_22336_, _02958_, _02039_);
  nand (_22337_, _22336_, _05082_);
  or (_22338_, _22337_, _22335_);
  or (_22339_, _05082_, _04592_);
  and (_22340_, _22339_, _05087_);
  and (_22341_, _22340_, _22338_);
  or (_22343_, _22194_, \oc8051_golden_model_1.PSW [7]);
  or (_22344_, _04592_, _05092_);
  and (_22345_, _22344_, _05086_);
  and (_22346_, _22345_, _22343_);
  or (_22347_, _22346_, _05097_);
  or (_22348_, _22347_, _22341_);
  and (_22349_, _22348_, _22152_);
  or (_22350_, _22349_, _05101_);
  or (_22351_, _05105_, _04592_);
  and (_22352_, _22351_, _05104_);
  and (_22354_, _22352_, _22350_);
  nand (_22355_, _02958_, _02016_);
  nand (_22356_, _22355_, _05110_);
  or (_22357_, _22356_, _22354_);
  or (_22358_, _05110_, _04592_);
  and (_22359_, _22358_, _05115_);
  and (_22360_, _22359_, _22357_);
  or (_22361_, _22194_, _05092_);
  or (_22362_, _04592_, \oc8051_golden_model_1.PSW [7]);
  and (_22363_, _22362_, _05114_);
  and (_22365_, _22363_, _22361_);
  or (_22366_, _22365_, _22360_);
  and (_22367_, _22366_, _05139_);
  and (_22368_, _22147_, _05141_);
  or (_22369_, _22368_, _02273_);
  or (_22370_, _22369_, _22367_);
  or (_22371_, _04592_, _05147_);
  and (_22372_, _22371_, _05146_);
  and (_22373_, _22372_, _22370_);
  and (_22374_, _22147_, _05145_);
  or (_22376_, _22374_, _02146_);
  or (_22377_, _22376_, _22373_);
  and (_22378_, _22377_, _22151_);
  or (_22379_, _22378_, _01660_);
  or (_22380_, _04592_, _05157_);
  and (_22381_, _22380_, _02153_);
  and (_22382_, _22381_, _22379_);
  or (_22383_, _22159_, _05387_);
  or (_22384_, _05386_, _02958_);
  and (_22385_, _22384_, _02015_);
  and (_22387_, _22385_, _22383_);
  or (_22388_, _22387_, _05161_);
  or (_22389_, _22388_, _22382_);
  and (_22390_, _22389_, _22150_);
  or (_22391_, _22390_, _02788_);
  or (_22392_, _04592_, _05398_);
  and (_22393_, _22392_, _05397_);
  and (_22394_, _22393_, _22391_);
  and (_22395_, _22147_, _05396_);
  or (_22396_, _22395_, _01585_);
  or (_22398_, _22396_, _22394_);
  and (_22399_, _22398_, _22149_);
  or (_22400_, _22399_, _01581_);
  or (_22401_, _04592_, _05407_);
  and (_22402_, _22401_, _02558_);
  and (_22403_, _22402_, _22400_);
  nand (_22404_, _05386_, _02959_);
  or (_22405_, _22159_, _05386_);
  and (_22406_, _22405_, _22404_);
  and (_22407_, _22406_, _02022_);
  or (_22409_, _22407_, _05419_);
  or (_22410_, _22409_, _22403_);
  or (_22411_, _22147_, _05418_);
  and (_22412_, _22411_, _02168_);
  and (_22413_, _22412_, _22410_);
  and (_22414_, _04592_, _02164_);
  or (_22415_, _22414_, _05426_);
  or (_22416_, _22415_, _22413_);
  or (_22417_, _22147_, _05430_);
  and (_22418_, _22417_, _05429_);
  and (_22420_, _22418_, _22416_);
  nor (_22421_, _02214_, _05429_);
  or (_22422_, _22421_, _01670_);
  or (_22423_, _22422_, _22420_);
  or (_22424_, _04592_, _01671_);
  and (_22425_, _22424_, _02377_);
  and (_22426_, _22425_, _22423_);
  and (_22427_, _22406_, _02025_);
  or (_22428_, _22427_, _05446_);
  or (_22429_, _22428_, _22426_);
  or (_22431_, _22147_, _05445_);
  and (_22432_, _22431_, _01595_);
  and (_22433_, _22432_, _22429_);
  and (_22434_, _04592_, _01594_);
  or (_22435_, _22434_, _05453_);
  or (_22436_, _22435_, _22433_);
  or (_22437_, _22147_, _05457_);
  and (_22438_, _22437_, _05456_);
  and (_22439_, _22438_, _22436_);
  nor (_22440_, _02214_, _05456_);
  or (_22442_, _22440_, _01657_);
  or (_22443_, _22442_, _22439_);
  or (_22444_, _04592_, _01658_);
  and (_22445_, _22444_, _05465_);
  and (_22446_, _22445_, _22443_);
  or (_22447_, _22446_, _22148_);
  or (_22448_, _22447_, _26506_);
  or (_22449_, _26505_, \oc8051_golden_model_1.PC [13]);
  and (_22450_, _22449_, _25964_);
  and (_27929_, _22450_, _22448_);
  and (_22452_, _04586_, _01594_);
  nor (_22453_, _05022_, _04586_);
  and (_22454_, _04874_, _02945_);
  and (_22455_, _03163_, _02950_);
  nor (_22456_, _22455_, _03165_);
  not (_22457_, _22456_);
  nor (_22458_, _22457_, _04874_);
  nor (_22459_, _22458_, _22454_);
  or (_22460_, _22459_, _02378_);
  or (_22461_, _22456_, _03909_);
  nand (_22463_, _03909_, _02946_);
  nand (_22464_, _22463_, _22461_);
  nand (_22465_, _22464_, _03185_);
  and (_22466_, _04085_, _02945_);
  nor (_22467_, _22457_, _04085_);
  or (_22468_, _22467_, _22466_);
  nor (_22469_, _22468_, _04090_);
  nor (_22470_, _02799_, \oc8051_golden_model_1.PC [14]);
  nor (_22471_, _22470_, _02800_);
  and (_22472_, _22471_, _04734_);
  nor (_22474_, _04720_, _04586_);
  nand (_22475_, _04553_, _02945_);
  or (_22476_, _22457_, _04553_);
  and (_22477_, _22476_, _01969_);
  and (_22478_, _22477_, _22475_);
  and (_22479_, _04710_, _04585_);
  and (_22480_, _04692_, _04590_);
  nor (_22481_, _22480_, _04693_);
  and (_22482_, _22481_, _04707_);
  nor (_22483_, _22482_, _22479_);
  nand (_22485_, _22483_, _04557_);
  nor (_22486_, _04586_, _01627_);
  and (_22487_, _04571_, _04586_);
  nand (_22488_, _18340_, \oc8051_golden_model_1.PC [14]);
  and (_22489_, _22488_, _05488_);
  or (_22490_, _04559_, _04563_);
  or (_22491_, _22490_, _22489_);
  and (_22492_, _22491_, _02424_);
  or (_22493_, _22492_, _22487_);
  and (_22494_, _22493_, _01625_);
  or (_22496_, _22494_, _04562_);
  not (_22497_, _22471_);
  or (_22498_, _22497_, _04565_);
  and (_22499_, _22498_, _22496_);
  nor (_22500_, _01971_, _04568_);
  nor (_22501_, _22500_, _04585_);
  or (_22502_, _22501_, _04558_);
  nor (_22503_, _22502_, _22499_);
  or (_22504_, _22503_, _04557_);
  nor (_22505_, _22504_, _22486_);
  nor (_22507_, _22505_, _04715_);
  nand (_22508_, _22507_, _22485_);
  and (_22509_, _22471_, _04715_);
  nor (_22510_, _22509_, _01969_);
  and (_22511_, _22510_, _22508_);
  or (_22512_, _22511_, _22478_);
  nand (_22513_, _22512_, _17940_);
  nor (_22514_, _22471_, _17940_);
  nor (_22515_, _22514_, _21858_);
  and (_22516_, _22515_, _22513_);
  nor (_22518_, _22516_, _22474_);
  or (_22519_, _22518_, _04725_);
  nand (_22520_, _22471_, _04725_);
  and (_22521_, _22520_, _01964_);
  nand (_22522_, _22521_, _22519_);
  and (_22523_, _04586_, _01963_);
  nor (_22524_, _22523_, _04734_);
  and (_22525_, _22524_, _22522_);
  or (_22526_, _22525_, _22472_);
  nand (_22527_, _22526_, _04738_);
  nor (_22529_, _04738_, _04586_);
  nor (_22530_, _22529_, _04089_);
  and (_22531_, _22530_, _22527_);
  or (_22532_, _22531_, _22469_);
  nand (_22533_, _22532_, _03187_);
  nand (_22534_, _22533_, _22465_);
  or (_22535_, _22534_, _01951_);
  and (_22536_, _22535_, _22460_);
  or (_22537_, _22536_, _03179_);
  nand (_22538_, _02945_, _02912_);
  nand (_22540_, _22456_, _19160_);
  and (_22541_, _22540_, _22538_);
  or (_22542_, _22541_, _04749_);
  and (_22543_, _22542_, _22537_);
  or (_22544_, _22543_, _02880_);
  nand (_22545_, _22471_, _02880_);
  and (_22546_, _22545_, _22544_);
  and (_22547_, _22546_, _04899_);
  nor (_22548_, _04899_, _04585_);
  or (_22549_, _22548_, _22547_);
  nand (_22551_, _22549_, _04905_);
  nor (_22552_, _22471_, _04905_);
  nor (_22553_, _22552_, _04911_);
  nand (_22554_, _22553_, _22551_);
  nor (_22555_, _04910_, _04586_);
  nor (_22556_, _22555_, _04933_);
  nand (_22557_, _22556_, _22554_);
  nor (_22558_, _22471_, _04928_);
  nor (_22559_, _22558_, _04932_);
  and (_22560_, _22559_, _22557_);
  and (_22562_, _04585_, _04932_);
  or (_22563_, _22562_, _01611_);
  or (_22564_, _22563_, _22560_);
  nor (_22565_, _22471_, _01616_);
  nor (_22566_, _22565_, _04943_);
  nand (_22567_, _22566_, _22564_);
  nor (_22568_, _04942_, _04586_);
  nor (_22569_, _22568_, _02001_);
  nand (_22570_, _22569_, _22567_);
  and (_22571_, _02946_, _02001_);
  nor (_22573_, _22571_, _04953_);
  nand (_22574_, _22573_, _22570_);
  nor (_22575_, _04952_, _04586_);
  nor (_22576_, _22575_, _01602_);
  and (_22577_, _22576_, _22574_);
  nor (_22578_, _04960_, _02946_);
  nor (_22579_, _22578_, _17728_);
  or (_22580_, _22579_, _22577_);
  and (_22581_, _22471_, _04960_);
  nor (_22582_, _22581_, _04964_);
  nand (_22584_, _22582_, _22580_);
  nor (_22585_, _04963_, _04585_);
  nor (_22586_, _22585_, _04968_);
  nand (_22587_, _22586_, _22584_);
  and (_22588_, _22481_, _04968_);
  nor (_22589_, _22588_, _02859_);
  and (_22590_, _22589_, _22587_);
  and (_22591_, _02859_, _04586_);
  or (_22592_, _22591_, _22590_);
  nand (_22593_, _22592_, _04979_);
  and (_22595_, _02946_, _02019_);
  nor (_22596_, _22595_, _02853_);
  nand (_22597_, _22596_, _22593_);
  and (_22598_, _04585_, _02853_);
  nor (_22599_, _22598_, _04984_);
  nand (_22600_, _22599_, _22597_);
  nor (_22601_, _05016_, \oc8051_golden_model_1.DPH [6]);
  nor (_22602_, _22601_, _05017_);
  nor (_22603_, _22602_, _04985_);
  nor (_22604_, _22603_, _05023_);
  and (_22605_, _22604_, _22600_);
  or (_22606_, _22605_, _22453_);
  nand (_22607_, _22606_, _05027_);
  and (_22608_, _05038_, _04585_);
  and (_22609_, _22481_, _05040_);
  or (_22610_, _22609_, _22608_);
  and (_22611_, _22610_, _05026_);
  nor (_22612_, _22611_, _05031_);
  nand (_22613_, _22612_, _22607_);
  nor (_22614_, _22471_, _02830_);
  nor (_22616_, _22614_, _05047_);
  and (_22617_, _22616_, _22613_);
  and (_22618_, _05047_, _04585_);
  or (_22619_, _22618_, _02018_);
  or (_22620_, _22619_, _22617_);
  and (_22621_, _02946_, _02018_);
  nor (_22622_, _22621_, _05056_);
  and (_22623_, _22622_, _22620_);
  nor (_22624_, _05055_, _04586_);
  or (_22625_, _22624_, _22623_);
  nand (_22627_, _22625_, _05060_);
  and (_22628_, _05040_, _04585_);
  and (_22629_, _22481_, _05038_);
  or (_22630_, _22629_, _22628_);
  and (_22631_, _22630_, _05059_);
  nor (_22632_, _22631_, _05069_);
  nand (_22633_, _22632_, _22627_);
  nor (_22634_, _22471_, _05070_);
  nor (_22635_, _22634_, _05072_);
  and (_22636_, _22635_, _22633_);
  and (_22638_, _04585_, _05072_);
  or (_22639_, _22638_, _02039_);
  or (_22640_, _22639_, _22636_);
  nand (_22641_, _02946_, _02039_);
  and (_22642_, _22641_, _05082_);
  and (_22643_, _22642_, _22640_);
  nor (_22644_, _05082_, _04586_);
  or (_22645_, _22644_, _22643_);
  nand (_22646_, _22645_, _05087_);
  nor (_22647_, _22481_, \oc8051_golden_model_1.PSW [7]);
  nor (_22649_, _04585_, _05092_);
  nor (_22650_, _22649_, _05087_);
  not (_22651_, _22650_);
  nor (_22652_, _22651_, _22647_);
  nor (_22653_, _22652_, _05097_);
  nand (_22654_, _22653_, _22646_);
  nor (_22655_, _22471_, _05098_);
  nor (_22656_, _22655_, _05101_);
  and (_22657_, _22656_, _22654_);
  and (_22658_, _05101_, _04585_);
  or (_22660_, _22658_, _02016_);
  or (_22661_, _22660_, _22657_);
  and (_22662_, _02946_, _02016_);
  nor (_22663_, _22662_, _05111_);
  and (_22664_, _22663_, _22661_);
  nor (_22665_, _05110_, _04586_);
  or (_22666_, _22665_, _22664_);
  nand (_22667_, _22666_, _05115_);
  nor (_22668_, _22481_, _05092_);
  nor (_22669_, _04585_, \oc8051_golden_model_1.PSW [7]);
  nor (_22671_, _22669_, _05115_);
  not (_22672_, _22671_);
  nor (_22673_, _22672_, _22668_);
  nor (_22674_, _22673_, _05141_);
  nand (_22675_, _22674_, _22667_);
  nor (_22676_, _22471_, _05139_);
  nor (_22677_, _22676_, _02273_);
  and (_22678_, _22677_, _22675_);
  and (_22679_, _04585_, _02273_);
  or (_22680_, _22679_, _22678_);
  and (_22682_, _22680_, _05146_);
  and (_22683_, _22471_, _05145_);
  or (_22684_, _22683_, _22682_);
  and (_22685_, _22684_, _02718_);
  nor (_22686_, _04074_, _02718_);
  or (_22687_, _22686_, _01660_);
  or (_22688_, _22687_, _22685_);
  and (_22689_, _04586_, _01660_);
  nor (_22690_, _22689_, _02015_);
  nand (_22691_, _22690_, _22688_);
  and (_22693_, _22457_, _05386_);
  nor (_22694_, _05386_, _02945_);
  or (_22695_, _22694_, _02153_);
  nor (_22696_, _22695_, _22693_);
  nor (_22697_, _22696_, _05161_);
  nand (_22698_, _22697_, _22691_);
  nor (_22699_, _22471_, _02818_);
  nor (_22700_, _22699_, _02788_);
  and (_22701_, _22700_, _22698_);
  and (_22702_, _04585_, _02788_);
  or (_22704_, _22702_, _22701_);
  and (_22705_, _22704_, _05397_);
  and (_22706_, _22471_, _05396_);
  or (_22707_, _22706_, _01585_);
  or (_22708_, _22707_, _22705_);
  and (_22709_, _04074_, _01585_);
  nor (_22710_, _22709_, _01581_);
  and (_22711_, _22710_, _22708_);
  and (_22712_, _04585_, _01581_);
  or (_22713_, _22712_, _02022_);
  nor (_22715_, _22713_, _22711_);
  and (_22716_, _05386_, _02946_);
  nor (_22717_, _22456_, _05386_);
  nor (_22718_, _22717_, _22716_);
  nor (_22719_, _22718_, _02558_);
  or (_22720_, _22719_, _22715_);
  and (_22721_, _22720_, _05418_);
  nor (_22722_, _22471_, _05418_);
  or (_22723_, _22722_, _22721_);
  nand (_22724_, _22723_, _02168_);
  and (_22726_, _04586_, _02164_);
  nor (_22727_, _22726_, _05426_);
  nand (_22728_, _22727_, _22724_);
  and (_22729_, _22471_, _05426_);
  nor (_22730_, _22729_, _02023_);
  nand (_22731_, _22730_, _22728_);
  and (_22732_, _02023_, _01884_);
  nor (_22733_, _22732_, _01670_);
  nand (_22734_, _22733_, _22731_);
  and (_22735_, _04585_, _01670_);
  nor (_22737_, _22735_, _02025_);
  nand (_22738_, _22737_, _22734_);
  nor (_22739_, _22718_, _02377_);
  nor (_22740_, _22739_, _05446_);
  nand (_22741_, _22740_, _22738_);
  and (_22742_, _22471_, _05446_);
  nor (_22743_, _22742_, _01594_);
  and (_22744_, _22743_, _22741_);
  or (_22745_, _22744_, _22452_);
  nand (_22746_, _22745_, _05457_);
  nor (_22748_, _22471_, _05457_);
  nor (_22749_, _22748_, _02026_);
  and (_22750_, _22749_, _22746_);
  and (_22751_, _01884_, _01658_);
  nor (_22752_, _22751_, _17603_);
  or (_22753_, _22752_, _22750_);
  and (_22754_, _04586_, _01657_);
  nor (_22755_, _22754_, _05464_);
  and (_22756_, _22755_, _22753_);
  and (_22757_, _22471_, _05464_);
  or (_22759_, _22757_, _22756_);
  or (_22760_, _22759_, _26506_);
  or (_22761_, _26505_, \oc8051_golden_model_1.PC [14]);
  and (_22762_, _22761_, _25964_);
  and (_27930_, _22762_, _22760_);
  and (_22763_, _26506_, \oc8051_golden_model_1.P0INREG [0]);
  or (_22764_, _22763_, _26557_);
  and (_27931_, _22764_, _25964_);
  and (_22765_, _26506_, \oc8051_golden_model_1.P0INREG [1]);
  or (_22766_, _22765_, _26525_);
  and (_27932_, _22766_, _25964_);
  and (_22768_, _26506_, \oc8051_golden_model_1.P0INREG [2]);
  or (_22769_, _22768_, _26516_);
  and (_27935_, _22769_, _25964_);
  and (_22770_, _26506_, \oc8051_golden_model_1.P0INREG [3]);
  or (_22771_, _22770_, _26548_);
  and (_27936_, _22771_, _25964_);
  and (_22772_, _26506_, \oc8051_golden_model_1.P0INREG [4]);
  or (_22773_, _22772_, _26564_);
  and (_27937_, _22773_, _25964_);
  and (_22775_, _26506_, \oc8051_golden_model_1.P0INREG [5]);
  or (_22776_, _22775_, _26532_);
  and (_27938_, _22776_, _25964_);
  and (_22777_, _26506_, \oc8051_golden_model_1.P0INREG [6]);
  or (_22778_, _22777_, _26508_);
  and (_27939_, _22778_, _25964_);
  and (_22779_, _26506_, \oc8051_golden_model_1.P1INREG [0]);
  or (_22780_, _22779_, _26785_);
  and (_27942_, _22780_, _25964_);
  and (_22781_, _26506_, \oc8051_golden_model_1.P1INREG [1]);
  or (_22783_, _22781_, _26763_);
  and (_27943_, _22783_, _25964_);
  and (_22784_, _26506_, \oc8051_golden_model_1.P1INREG [2]);
  or (_22785_, _22784_, _26778_);
  and (_27944_, _22785_, _25964_);
  and (_22786_, _26506_, \oc8051_golden_model_1.P1INREG [3]);
  or (_22787_, _22786_, _26770_);
  and (_27945_, _22787_, _25964_);
  and (_22788_, _26506_, \oc8051_golden_model_1.P1INREG [4]);
  or (_22789_, _22788_, _26731_);
  and (_27946_, _22789_, _25964_);
  and (_22791_, _26506_, \oc8051_golden_model_1.P1INREG [5]);
  or (_22792_, _22791_, _26746_);
  and (_27947_, _22792_, _25964_);
  and (_22793_, _26506_, \oc8051_golden_model_1.P1INREG [6]);
  or (_22794_, _22793_, _26738_);
  and (_27948_, _22794_, _25964_);
  and (_22795_, _26506_, \oc8051_golden_model_1.P2INREG [0]);
  or (_22796_, _22795_, _26616_);
  and (_27949_, _22796_, _25964_);
  and (_22798_, _26506_, \oc8051_golden_model_1.P2INREG [1]);
  or (_22799_, _22798_, _26600_);
  and (_27950_, _22799_, _25964_);
  and (_22800_, _26506_, \oc8051_golden_model_1.P2INREG [2]);
  or (_22801_, _22800_, _26577_);
  and (_27951_, _22801_, _25964_);
  and (_22802_, _26506_, \oc8051_golden_model_1.P2INREG [3]);
  or (_22803_, _22802_, _26625_);
  and (_27952_, _22803_, _25964_);
  and (_22804_, _26506_, \oc8051_golden_model_1.P2INREG [4]);
  or (_22806_, _22804_, _26609_);
  and (_27955_, _22806_, _25964_);
  and (_22807_, _26506_, \oc8051_golden_model_1.P2INREG [5]);
  or (_22808_, _22807_, _26593_);
  and (_27956_, _22808_, _25964_);
  and (_22809_, _26506_, \oc8051_golden_model_1.P2INREG [6]);
  or (_22810_, _22809_, _26584_);
  and (_27957_, _22810_, _25964_);
  and (_22811_, _26506_, \oc8051_golden_model_1.P3INREG [0]);
  or (_22812_, _22811_, _26841_);
  and (_27960_, _22812_, _25964_);
  and (_22814_, _26506_, \oc8051_golden_model_1.P3INREG [1]);
  or (_22815_, _22814_, _26874_);
  and (_27961_, _22815_, _25964_);
  and (_22816_, _26506_, \oc8051_golden_model_1.P3INREG [2]);
  or (_22817_, _22816_, _26857_);
  and (_27962_, _22817_, _25964_);
  and (_22818_, _26506_, \oc8051_golden_model_1.P3INREG [3]);
  or (_22819_, _22818_, _26867_);
  and (_27963_, _22819_, _25964_);
  and (_22821_, _26506_, \oc8051_golden_model_1.P3INREG [4]);
  or (_22822_, _22821_, _26834_);
  and (_27964_, _22822_, _25964_);
  and (_22823_, _26506_, \oc8051_golden_model_1.P3INREG [5]);
  or (_22824_, _22823_, _26825_);
  and (_27965_, _22824_, _25964_);
  and (_22825_, _26506_, \oc8051_golden_model_1.P3INREG [6]);
  or (_22826_, _22825_, _26850_);
  and (_27966_, _22826_, _25964_);
  and (_00005_[6], _26851_, _25964_);
  and (_00005_[5], _26826_, _25964_);
  and (_00005_[4], _26835_, _25964_);
  and (_00005_[3], _26868_, _25964_);
  and (_00005_[2], _26858_, _25964_);
  and (_00005_[1], _26875_, _25964_);
  and (_00005_[0], _26842_, _25964_);
  and (_00004_[6], _26585_, _25964_);
  and (_00004_[5], _26594_, _25964_);
  and (_00004_[4], _26610_, _25964_);
  and (_00004_[3], _26626_, _25964_);
  and (_00004_[2], _26578_, _25964_);
  and (_00004_[1], _26601_, _25964_);
  and (_00004_[0], _26617_, _25964_);
  and (_00003_[6], _26739_, _25964_);
  and (_00003_[5], _26747_, _25964_);
  and (_00003_[4], _26732_, _25964_);
  and (_00003_[3], _26771_, _25964_);
  and (_00003_[2], _26779_, _25964_);
  and (_00003_[1], _26764_, _25964_);
  and (_00003_[0], _26786_, _25964_);
  and (_00001_[6], _26509_, _25964_);
  and (_00001_[5], _26533_, _25964_);
  and (_00001_[4], _26565_, _25964_);
  and (_00001_[3], _26549_, _25964_);
  and (_00001_[2], _26517_, _25964_);
  and (_00001_[1], _26526_, _25964_);
  and (_00001_[0], _26558_, _25964_);
  and (_00004_[7], _26633_, _25964_);
  and (_00005_[7], _26819_, _25964_);
  nand (_22830_, _18297_, _27466_);
  or (_22832_, _18297_, _27466_);
  and (_22833_, _18673_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_22834_, _19395_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_22835_, _18673_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_22836_, _22835_, _22834_);
  nor (_22837_, _22836_, _22833_);
  or (_22838_, _20133_, _27428_);
  nand (_22839_, _20133_, _27428_);
  nand (_22840_, _22839_, _22838_);
  or (_22841_, _19033_, _27452_);
  and (_22843_, _21178_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_22844_, _21178_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_22845_, _20842_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_22846_, _20842_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_22847_, _21499_, _27423_);
  nand (_22848_, _21499_, _27423_);
  nand (_22849_, _22848_, _22847_);
  or (_22850_, _22759_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_22851_, _22759_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_22852_, _22851_, _22850_);
  and (_22854_, _21828_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_22855_, _21828_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_22856_, _17864_, _27473_);
  and (_22857_, _17864_, _27473_);
  nor (_22858_, _22857_, _22856_);
  and (_22859_, _22447_, _27419_);
  nor (_22860_, _22447_, _27419_);
  or (_22861_, _22860_, _22859_);
  nor (_22862_, _22861_, _22858_);
  nand (_22863_, _22862_, _22855_);
  nor (_22865_, _22863_, _22854_);
  nor (_22866_, _05470_, _27278_);
  and (_22867_, _05470_, _27278_);
  nor (_22868_, _22867_, _22866_);
  and (_22869_, _22868_, _22865_);
  and (_22870_, _22869_, _22852_);
  nor (_22871_, _22141_, _27420_);
  and (_22872_, _22141_, _27420_);
  nor (_22873_, _22872_, _22871_);
  and (_22874_, _22873_, _22870_);
  and (_22876_, _22874_, _22849_);
  nand (_22877_, _22876_, _22846_);
  nor (_22878_, _22877_, _22845_);
  nand (_22879_, _22878_, _22844_);
  nor (_22880_, _22879_, _22843_);
  and (_22881_, _22880_, _22841_);
  or (_22882_, _19771_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_22883_, _20503_, _27425_);
  and (_22884_, _22883_, _22882_);
  and (_22885_, _22884_, _22881_);
  and (_22887_, _22885_, _22840_);
  nand (_22888_, _19395_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_22889_, _19771_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_22890_, _19033_, _27452_);
  nand (_22891_, _20503_, _27425_);
  nand (_22892_, _22891_, _22890_);
  nor (_22893_, _22892_, _22889_);
  and (_22894_, _22893_, _22888_);
  and (_22895_, _22894_, _22887_);
  and (_22896_, _22895_, _22837_);
  and (_22898_, _22896_, _22832_);
  and (_22899_, _22898_, _22830_);
  and (_22900_, _26505_, eq_state);
  and (_22901_, _22900_, _01589_);
  nand (_22902_, _22901_, _02852_);
  nor (property_invalid_pc, _22902_, _22899_);
  nor (_22903_, _11030_, _10315_);
  nor (_22904_, _14350_, _12903_);
  and (_22905_, _22904_, _22903_);
  nor (_22906_, _06583_, _06327_);
  nor (_22908_, _06965_, _06858_);
  and (_22909_, _22908_, _22906_);
  nor (_22910_, _14661_, _13214_);
  nor (_22911_, _11341_, _10626_);
  and (_22912_, _22911_, _22910_);
  nor (_22913_, _12697_, _10824_);
  and (_22914_, _22913_, _14144_);
  nor (_22915_, _06664_, _06200_);
  nor (_22916_, _10109_, _06745_);
  and (_22917_, _22916_, _22915_);
  and (_22919_, _22917_, _22914_);
  and (_22920_, _22919_, _12598_);
  nor (_22921_, _16824_, _16307_);
  nor (_22922_, _17426_, _16913_);
  and (_22923_, _22922_, _22921_);
  nor (_22924_, _15610_, _15051_);
  nor (_22925_, _16219_, _15698_);
  and (_22926_, _22925_, _22924_);
  or (_22927_, _17514_, _17168_);
  or (_22928_, _22927_, _17599_);
  nor (_22930_, _22928_, _11771_);
  nor (_22931_, _12343_, _11851_);
  and (_22932_, _22931_, _22930_);
  and (_22933_, _22932_, _22926_);
  and (_22934_, _22933_, _22923_);
  nor (_22935_, _05930_, _05767_);
  nor (_22936_, _06119_, _06037_);
  and (_22937_, _22936_, _22935_);
  nor (_22938_, _15131_, _14814_);
  nor (_22939_, _15361_, _15209_);
  and (_22941_, _22939_, _22938_);
  nor (_22942_, _12081_, _11929_);
  nor (_22943_, _12501_, _12423_);
  and (_22944_, _22943_, _22942_);
  and (_22945_, _22944_, _22941_);
  nor (_22946_, _16560_, _16394_);
  nor (_22947_, _16998_, _16735_);
  and (_22948_, _22947_, _22946_);
  nor (_22949_, _15784_, _15522_);
  nor (_22950_, _16130_, _15954_);
  and (_22952_, _22950_, _22949_);
  and (_22953_, _22952_, _22948_);
  and (_22954_, _22953_, _22945_);
  and (_22955_, _10725_, _10007_);
  and (_22956_, _22955_, _14046_);
  nor (_22957_, _15867_, _15282_);
  nor (_22958_, _17082_, _16474_);
  and (_22959_, _22958_, _22957_);
  nor (_22960_, \oc8051_golden_model_1.IE [7], \oc8051_golden_model_1.IP [7]);
  nor (_22961_, \oc8051_golden_model_1.SCON [7], \oc8051_golden_model_1.SBUF [7]);
  nor (_22963_, \oc8051_golden_model_1.TL1 [7], \oc8051_golden_model_1.TH1 [7]);
  and (_22964_, _22963_, _22961_);
  and (_22965_, _22964_, _22960_);
  nor (_22966_, \oc8051_golden_model_1.IP [1], \oc8051_golden_model_1.IP [0]);
  nor (_22967_, \oc8051_golden_model_1.IP [2], \oc8051_golden_model_1.PCON [7]);
  and (_22968_, _22967_, _22966_);
  nor (_22969_, \oc8051_golden_model_1.TL0 [7], \oc8051_golden_model_1.TH0 [7]);
  nor (_22970_, \oc8051_golden_model_1.TCON [7], \oc8051_golden_model_1.TMOD [7]);
  and (_22971_, _22970_, _22969_);
  and (_22972_, _22971_, _22968_);
  and (_22974_, _22972_, _22965_);
  nor (_22975_, \oc8051_golden_model_1.SBUF [3], \oc8051_golden_model_1.SBUF [2]);
  nor (_22976_, \oc8051_golden_model_1.SBUF [4], \oc8051_golden_model_1.SBUF [1]);
  and (_22977_, _22976_, _22975_);
  nor (_22978_, \oc8051_golden_model_1.IE [5], \oc8051_golden_model_1.IE [4]);
  nor (_22979_, \oc8051_golden_model_1.SBUF [0], \oc8051_golden_model_1.IE [6]);
  and (_22980_, _22979_, _22978_);
  and (_22981_, _22980_, _22977_);
  nor (_22982_, \oc8051_golden_model_1.IE [1], \oc8051_golden_model_1.IE [0]);
  nor (_22983_, \oc8051_golden_model_1.IE [3], \oc8051_golden_model_1.IE [2]);
  and (_22985_, _22983_, _22982_);
  nor (_22986_, \oc8051_golden_model_1.IP [4], \oc8051_golden_model_1.IP [3]);
  nor (_22987_, \oc8051_golden_model_1.IP [6], \oc8051_golden_model_1.IP [5]);
  and (_22988_, _22987_, _22986_);
  and (_22989_, _22988_, _22985_);
  and (_22990_, _22989_, _22981_);
  and (_22991_, _22990_, _22974_);
  nor (_22992_, \oc8051_golden_model_1.SCON [3], \oc8051_golden_model_1.SCON [2]);
  nor (_22993_, \oc8051_golden_model_1.SCON [5], \oc8051_golden_model_1.SCON [4]);
  and (_22994_, _22993_, _22992_);
  nor (_22996_, \oc8051_golden_model_1.SCON [1], \oc8051_golden_model_1.SCON [0]);
  nor (_22997_, \oc8051_golden_model_1.SBUF [6], \oc8051_golden_model_1.SBUF [5]);
  and (_22998_, _22997_, _22996_);
  and (_22999_, _22998_, _22994_);
  nor (_23000_, \oc8051_golden_model_1.TH1 [5], \oc8051_golden_model_1.TH1 [4]);
  nor (_23001_, \oc8051_golden_model_1.TH1 [6], \oc8051_golden_model_1.TH1 [3]);
  and (_23002_, _23001_, _23000_);
  nor (_23003_, \oc8051_golden_model_1.TH1 [0], \oc8051_golden_model_1.SCON [6]);
  nor (_23004_, \oc8051_golden_model_1.TH1 [2], \oc8051_golden_model_1.TH1 [1]);
  and (_23005_, _23004_, _23003_);
  and (_23007_, _23005_, _23002_);
  and (_23008_, _23007_, _22999_);
  nor (_23009_, \oc8051_golden_model_1.TL1 [1], \oc8051_golden_model_1.TL1 [0]);
  nor (_23010_, \oc8051_golden_model_1.TL1 [3], \oc8051_golden_model_1.TL1 [2]);
  and (_23011_, _23010_, _23009_);
  nor (_23012_, \oc8051_golden_model_1.TL1 [5], \oc8051_golden_model_1.TL1 [4]);
  nor (_23013_, \oc8051_golden_model_1.TH0 [0], \oc8051_golden_model_1.TL1 [6]);
  and (_23014_, _23013_, _23012_);
  and (_23015_, _23014_, _23011_);
  nor (_23016_, \oc8051_golden_model_1.TL0 [1], \oc8051_golden_model_1.TL0 [0]);
  nor (_23018_, \oc8051_golden_model_1.TH0 [6], \oc8051_golden_model_1.TH0 [5]);
  and (_23019_, _23018_, _23016_);
  nor (_23020_, \oc8051_golden_model_1.TH0 [2], \oc8051_golden_model_1.TH0 [1]);
  nor (_23021_, \oc8051_golden_model_1.TH0 [4], \oc8051_golden_model_1.TH0 [3]);
  and (_23022_, _23021_, _23020_);
  and (_23023_, _23022_, _23019_);
  and (_23024_, _23023_, _23015_);
  and (_23025_, _23024_, _23008_);
  nor (_23026_, \oc8051_golden_model_1.PCON [6], \oc8051_golden_model_1.PCON [5]);
  and (_23027_, _23026_, regs_always_zero);
  nor (_23029_, \oc8051_golden_model_1.PCON [3], \oc8051_golden_model_1.PCON [2]);
  nor (_23030_, \oc8051_golden_model_1.PCON [4], \oc8051_golden_model_1.PCON [1]);
  and (_23031_, _23030_, _23029_);
  nor (_23032_, \oc8051_golden_model_1.TCON [5], \oc8051_golden_model_1.TCON [4]);
  nor (_23033_, \oc8051_golden_model_1.PCON [0], \oc8051_golden_model_1.TCON [6]);
  and (_23034_, _23033_, _23032_);
  and (_23035_, _23034_, _23031_);
  and (_23036_, _23035_, _23027_);
  and (_23037_, \oc8051_golden_model_1.TCON [1], _13951_);
  nor (_23038_, \oc8051_golden_model_1.TCON [3], \oc8051_golden_model_1.TCON [2]);
  and (_23040_, _23038_, _23037_);
  nor (_23041_, \oc8051_golden_model_1.TMOD [4], \oc8051_golden_model_1.TMOD [3]);
  nor (_23042_, \oc8051_golden_model_1.TMOD [6], \oc8051_golden_model_1.TMOD [5]);
  and (_23043_, _23042_, _23041_);
  and (_23044_, _23043_, _23040_);
  nor (_23045_, \oc8051_golden_model_1.TMOD [1], \oc8051_golden_model_1.TMOD [0]);
  nor (_23046_, \oc8051_golden_model_1.TMOD [2], \oc8051_golden_model_1.TL0 [6]);
  and (_23047_, _23046_, _23045_);
  nor (_23048_, \oc8051_golden_model_1.TL0 [3], \oc8051_golden_model_1.TL0 [2]);
  nor (_23049_, \oc8051_golden_model_1.TL0 [5], \oc8051_golden_model_1.TL0 [4]);
  and (_23051_, _23049_, _23048_);
  and (_23052_, _23051_, _23047_);
  and (_23053_, _23052_, _23044_);
  and (_23054_, _23053_, _23036_);
  and (_23055_, _23054_, _23025_);
  nand (_23056_, _23055_, _22991_);
  nor (_23057_, _23056_, _11452_);
  nor (_23058_, _14736_, _12003_);
  and (_23059_, _23058_, _23057_);
  and (_23060_, _23059_, _22959_);
  nor (_23062_, _12173_, _11610_);
  and (_23063_, _23062_, _23060_);
  nor (_23064_, _11690_, _11530_);
  and (_23065_, _23064_, _23063_);
  nor (_23066_, _17339_, _17253_);
  nor (_23067_, _16647_, _16041_);
  and (_23068_, _23067_, _23066_);
  nor (_23069_, _14893_, _12263_);
  nor (_23070_, _15440_, _14971_);
  and (_23071_, _23070_, _23069_);
  and (_23073_, _23071_, _23068_);
  and (_23074_, _23073_, _23065_);
  and (_23075_, _23074_, _22956_);
  and (_23076_, _23075_, _22954_);
  and (_23077_, _23076_, _22937_);
  and (_23078_, _23077_, _22934_);
  and (_23079_, _23078_, _22920_);
  and (_23080_, _23079_, _22912_);
  and (_23081_, _23080_, _22909_);
  and (_23082_, _23081_, _22905_);
  nor (_23083_, _14558_, _14454_);
  nor (_23084_, _14247_, _13111_);
  and (_23085_, _23084_, _23083_);
  nor (_23086_, _11238_, _11134_);
  nor (_23087_, _13007_, _12800_);
  and (_23088_, _23087_, _23086_);
  nor (_23089_, _10419_, _10212_);
  nor (_23090_, _10927_, _10523_);
  and (_23091_, _23090_, _23089_);
  and (_23092_, _23091_, _23088_);
  and (_23094_, _23092_, _23085_);
  and (_23095_, _23094_, _23082_);
  or (_00006_, _23095_, rst);
  and (_23096_, _23095_, _06750_);
  and (_00002_, _23096_, _22899_);
  or (_00000_, p1_valid_r, rst);
  and (_00001_[7], _26542_, _25964_);
  and (_00003_[7], _26754_, _25964_);
  buf (_00069_, _25964_);
  buf (_00120_, _25964_);
  buf (_00172_, _25964_);
  buf (_00224_, _25964_);
  buf (_00276_, _25964_);
  buf (_00328_, _25964_);
  buf (_00380_, _25964_);
  buf (_00432_, _25964_);
  buf (_00484_, _25964_);
  buf (_00536_, _25964_);
  buf (_00588_, _25964_);
  buf (_00640_, _25964_);
  buf (_00691_, _25964_);
  buf (_00743_, _25964_);
  buf (_00794_, _25964_);
  buf (_00846_, _25964_);
  buf (_03167_, _00922_);
  buf (_03170_, _00926_);
  buf (_03204_, _00922_);
  buf (_03207_, _00926_);
  buf (_05680_, _01067_);
  buf (_05682_, _01070_);
  buf (_05684_, _01073_);
  buf (_05686_, _01076_);
  buf (_05688_, _01079_);
  buf (_05690_, _01082_);
  buf (_05692_, _01085_);
  buf (_05694_, _01088_);
  buf (_05696_, _01091_);
  buf (_05698_, _01094_);
  buf (_05700_, _01097_);
  buf (_05702_, _01100_);
  buf (_05704_, _01103_);
  buf (_05706_, _01105_);
  buf (_05799_, _01067_);
  buf (_05801_, _01070_);
  buf (_05803_, _01073_);
  buf (_05805_, _01076_);
  buf (_05807_, _01079_);
  buf (_05809_, _01082_);
  buf (_05811_, _01085_);
  buf (_05813_, _01088_);
  buf (_05815_, _01091_);
  buf (_05817_, _01094_);
  buf (_05819_, _01097_);
  buf (_05821_, _01100_);
  buf (_05823_, _01103_);
  buf (_05825_, _01105_);
  buf (_08192_, _01527_);
  buf (_08296_, _01527_);
  dff (p0in_reg[0], _00001_[0]);
  dff (p0in_reg[1], _00001_[1]);
  dff (p0in_reg[2], _00001_[2]);
  dff (p0in_reg[3], _00001_[3]);
  dff (p0in_reg[4], _00001_[4]);
  dff (p0in_reg[5], _00001_[5]);
  dff (p0in_reg[6], _00001_[6]);
  dff (p0in_reg[7], _00001_[7]);
  dff (p1in_reg[0], _00003_[0]);
  dff (p1in_reg[1], _00003_[1]);
  dff (p1in_reg[2], _00003_[2]);
  dff (p1in_reg[3], _00003_[3]);
  dff (p1in_reg[4], _00003_[4]);
  dff (p1in_reg[5], _00003_[5]);
  dff (p1in_reg[6], _00003_[6]);
  dff (p1in_reg[7], _00003_[7]);
  dff (p2in_reg[0], _00004_[0]);
  dff (p2in_reg[1], _00004_[1]);
  dff (p2in_reg[2], _00004_[2]);
  dff (p2in_reg[3], _00004_[3]);
  dff (p2in_reg[4], _00004_[4]);
  dff (p2in_reg[5], _00004_[5]);
  dff (p2in_reg[6], _00004_[6]);
  dff (p2in_reg[7], _00004_[7]);
  dff (p3in_reg[0], _00005_[0]);
  dff (p3in_reg[1], _00005_[1]);
  dff (p3in_reg[2], _00005_[2]);
  dff (p3in_reg[3], _00005_[3]);
  dff (p3in_reg[4], _00005_[4]);
  dff (p3in_reg[5], _00005_[5]);
  dff (p3in_reg[6], _00005_[6]);
  dff (p3in_reg[7], _00005_[7]);
  dff (regs_always_zero, _00006_);
  dff (p1_valid_r, _00002_);
  dff (eq_state, _00000_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _00098_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _00100_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _00102_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _00104_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _00106_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _00108_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _00110_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _00066_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _00069_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _00149_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _00151_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _00153_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _00155_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _00157_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _00159_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _00161_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _00117_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _00120_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _00617_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _00619_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _00621_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _00623_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _00625_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _00627_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _00629_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _00585_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _00588_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _00669_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _00671_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _00673_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _00675_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _00677_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _00679_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _00681_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _00637_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _00640_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _00720_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _00722_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _00724_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _00726_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _00728_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _00730_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _00732_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _00688_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _00691_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _00772_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _00774_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _00776_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _00778_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _00780_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _00782_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _00784_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _00740_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _00743_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _00824_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _00826_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _00827_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _00829_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _00831_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _00833_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _00835_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _00792_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _00794_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _00875_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _00877_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _00879_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _00881_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _00883_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _00885_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _00887_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _00843_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _00846_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _00201_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _00203_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _00205_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _00207_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _00209_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _00211_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _00213_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _00169_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _00172_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _00253_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _00255_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _00257_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _00259_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _00261_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _00263_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _00265_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _00221_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _00224_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _00305_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _00307_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _00309_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _00311_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _00313_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _00315_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _00317_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _00273_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _00276_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _00357_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _00359_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _00361_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _00363_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _00365_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _00367_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _00369_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _00325_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _00328_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _00409_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _00411_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _00413_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _00415_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _00417_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _00419_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _00421_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _00377_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _00380_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _00461_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _00463_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _00465_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _00467_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _00469_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _00471_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _00473_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _00429_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _00432_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _00514_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _00516_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _00517_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _00519_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _00521_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _00523_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _00525_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _00481_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _00484_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _00566_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _00568_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _00570_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _00572_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _00574_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _00575_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _00577_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _00533_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _00536_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _29636_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _29637_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _29638_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _29639_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _29640_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _29641_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _29642_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _29643_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _29682_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _29683_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _29684_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _29685_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _29686_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _29687_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _29688_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _29689_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _29674_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _29675_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _29676_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _29677_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _29678_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _29679_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _29680_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _29681_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _29666_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _29667_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _29668_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _29669_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _29670_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _29671_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _29672_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _29673_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _29658_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _29659_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _29660_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _29661_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _29662_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _29663_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _29664_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _29665_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _29650_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _29651_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _29652_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _29653_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _29654_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _29655_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _29656_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _29657_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _25573_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _25574_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _29644_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _29645_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _29646_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _29647_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _29648_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _29649_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _29722_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _29723_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _29724_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _29725_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _29730_[4]);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _29730_[5]);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _29730_[6]);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _29730_[7]);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _29714_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _29715_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _29716_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _29717_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _29718_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _29719_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _29720_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _29721_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _29706_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _29707_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _29708_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _29709_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _29710_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _29711_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _29712_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _29713_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _29698_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _29699_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _29700_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _29701_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _29702_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _29703_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _29704_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _29705_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _29690_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _29691_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _29692_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _29693_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _29694_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _29695_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _29696_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _29697_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _29729_[0]);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _29729_[1]);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _29729_[2]);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _29729_[3]);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _29729_[4]);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _29729_[5]);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _29729_[6]);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _29729_[7]);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _29728_[0]);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _29728_[1]);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _29728_[2]);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _29728_[3]);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _29728_[4]);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _29728_[5]);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _29728_[6]);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _29728_[7]);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _29727_[0]);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _29727_[1]);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _29727_[2]);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _29727_[3]);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _29727_[4]);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _29727_[5]);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _29727_[6]);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _29727_[7]);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _29726_[0]);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _29726_[1]);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _29726_[2]);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _29726_[3]);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _29726_[4]);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _29726_[5]);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _29726_[6]);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _29726_[7]);
  dff (\oc8051_golden_model_1.B [0], _27719_);
  dff (\oc8051_golden_model_1.B [1], _27720_);
  dff (\oc8051_golden_model_1.B [2], _27723_);
  dff (\oc8051_golden_model_1.B [3], _27724_);
  dff (\oc8051_golden_model_1.B [4], _27725_);
  dff (\oc8051_golden_model_1.B [5], _27726_);
  dff (\oc8051_golden_model_1.B [6], _27727_);
  dff (\oc8051_golden_model_1.B [7], _25338_);
  dff (\oc8051_golden_model_1.ACC [0], _27729_);
  dff (\oc8051_golden_model_1.ACC [1], _27732_);
  dff (\oc8051_golden_model_1.ACC [2], _27733_);
  dff (\oc8051_golden_model_1.ACC [3], _27734_);
  dff (\oc8051_golden_model_1.ACC [4], _27735_);
  dff (\oc8051_golden_model_1.ACC [5], _27736_);
  dff (\oc8051_golden_model_1.ACC [6], _27737_);
  dff (\oc8051_golden_model_1.ACC [7], _25336_);
  dff (\oc8051_golden_model_1.DPL [0], _27739_);
  dff (\oc8051_golden_model_1.DPL [1], _27740_);
  dff (\oc8051_golden_model_1.DPL [2], _27741_);
  dff (\oc8051_golden_model_1.DPL [3], _27742_);
  dff (\oc8051_golden_model_1.DPL [4], _27743_);
  dff (\oc8051_golden_model_1.DPL [5], _27744_);
  dff (\oc8051_golden_model_1.DPL [6], _27745_);
  dff (\oc8051_golden_model_1.DPL [7], _25335_);
  dff (\oc8051_golden_model_1.DPH [0], _27750_);
  dff (\oc8051_golden_model_1.DPH [1], _27751_);
  dff (\oc8051_golden_model_1.DPH [2], _27752_);
  dff (\oc8051_golden_model_1.DPH [3], _27753_);
  dff (\oc8051_golden_model_1.DPH [4], _27754_);
  dff (\oc8051_golden_model_1.DPH [5], _27755_);
  dff (\oc8051_golden_model_1.DPH [6], _27756_);
  dff (\oc8051_golden_model_1.DPH [7], _25334_);
  dff (\oc8051_golden_model_1.IE [0], _27757_);
  dff (\oc8051_golden_model_1.IE [1], _27758_);
  dff (\oc8051_golden_model_1.IE [2], _27759_);
  dff (\oc8051_golden_model_1.IE [3], _27760_);
  dff (\oc8051_golden_model_1.IE [4], _27761_);
  dff (\oc8051_golden_model_1.IE [5], _27764_);
  dff (\oc8051_golden_model_1.IE [6], _27765_);
  dff (\oc8051_golden_model_1.IE [7], _25333_);
  dff (\oc8051_golden_model_1.IP [0], _27766_);
  dff (\oc8051_golden_model_1.IP [1], _27769_);
  dff (\oc8051_golden_model_1.IP [2], _27770_);
  dff (\oc8051_golden_model_1.IP [3], _27771_);
  dff (\oc8051_golden_model_1.IP [4], _27772_);
  dff (\oc8051_golden_model_1.IP [5], _27773_);
  dff (\oc8051_golden_model_1.IP [6], _27774_);
  dff (\oc8051_golden_model_1.IP [7], _25331_);
  dff (\oc8051_golden_model_1.P0 [0], _27777_);
  dff (\oc8051_golden_model_1.P0 [1], _27778_);
  dff (\oc8051_golden_model_1.P0 [2], _27779_);
  dff (\oc8051_golden_model_1.P0 [3], _27780_);
  dff (\oc8051_golden_model_1.P0 [4], _27781_);
  dff (\oc8051_golden_model_1.P0 [5], _27782_);
  dff (\oc8051_golden_model_1.P0 [6], _27783_);
  dff (\oc8051_golden_model_1.P0 [7], _25330_);
  dff (\oc8051_golden_model_1.P1 [0], _27786_);
  dff (\oc8051_golden_model_1.P1 [1], _27787_);
  dff (\oc8051_golden_model_1.P1 [2], _27788_);
  dff (\oc8051_golden_model_1.P1 [3], _27789_);
  dff (\oc8051_golden_model_1.P1 [4], _27790_);
  dff (\oc8051_golden_model_1.P1 [5], _27791_);
  dff (\oc8051_golden_model_1.P1 [6], _27792_);
  dff (\oc8051_golden_model_1.P1 [7], _25328_);
  dff (\oc8051_golden_model_1.P2 [0], _27797_);
  dff (\oc8051_golden_model_1.P2 [1], _27798_);
  dff (\oc8051_golden_model_1.P2 [2], _27799_);
  dff (\oc8051_golden_model_1.P2 [3], _27800_);
  dff (\oc8051_golden_model_1.P2 [4], _27801_);
  dff (\oc8051_golden_model_1.P2 [5], _27802_);
  dff (\oc8051_golden_model_1.P2 [6], _27803_);
  dff (\oc8051_golden_model_1.P2 [7], _25326_);
  dff (\oc8051_golden_model_1.P3 [0], _27806_);
  dff (\oc8051_golden_model_1.P3 [1], _27807_);
  dff (\oc8051_golden_model_1.P3 [2], _27808_);
  dff (\oc8051_golden_model_1.P3 [3], _27809_);
  dff (\oc8051_golden_model_1.P3 [4], _27810_);
  dff (\oc8051_golden_model_1.P3 [5], _27811_);
  dff (\oc8051_golden_model_1.P3 [6], _27812_);
  dff (\oc8051_golden_model_1.P3 [7], _25325_);
  dff (\oc8051_golden_model_1.PSW [0], _27815_);
  dff (\oc8051_golden_model_1.PSW [1], _27816_);
  dff (\oc8051_golden_model_1.PSW [2], _27817_);
  dff (\oc8051_golden_model_1.PSW [3], _27818_);
  dff (\oc8051_golden_model_1.PSW [4], _27819_);
  dff (\oc8051_golden_model_1.PSW [5], _27820_);
  dff (\oc8051_golden_model_1.PSW [6], _27823_);
  dff (\oc8051_golden_model_1.PSW [7], _25324_);
  dff (\oc8051_golden_model_1.PCON [0], _27824_);
  dff (\oc8051_golden_model_1.PCON [1], _27825_);
  dff (\oc8051_golden_model_1.PCON [2], _27828_);
  dff (\oc8051_golden_model_1.PCON [3], _27829_);
  dff (\oc8051_golden_model_1.PCON [4], _27830_);
  dff (\oc8051_golden_model_1.PCON [5], _27831_);
  dff (\oc8051_golden_model_1.PCON [6], _27832_);
  dff (\oc8051_golden_model_1.PCON [7], _25323_);
  dff (\oc8051_golden_model_1.SBUF [0], _27833_);
  dff (\oc8051_golden_model_1.SBUF [1], _27834_);
  dff (\oc8051_golden_model_1.SBUF [2], _27835_);
  dff (\oc8051_golden_model_1.SBUF [3], _27836_);
  dff (\oc8051_golden_model_1.SBUF [4], _27837_);
  dff (\oc8051_golden_model_1.SBUF [5], _27838_);
  dff (\oc8051_golden_model_1.SBUF [6], _27839_);
  dff (\oc8051_golden_model_1.SBUF [7], _25322_);
  dff (\oc8051_golden_model_1.SCON [0], _27842_);
  dff (\oc8051_golden_model_1.SCON [1], _27843_);
  dff (\oc8051_golden_model_1.SCON [2], _27844_);
  dff (\oc8051_golden_model_1.SCON [3], _27845_);
  dff (\oc8051_golden_model_1.SCON [4], _27848_);
  dff (\oc8051_golden_model_1.SCON [5], _27849_);
  dff (\oc8051_golden_model_1.SCON [6], _27850_);
  dff (\oc8051_golden_model_1.SCON [7], _25320_);
  dff (\oc8051_golden_model_1.SP [0], _27852_);
  dff (\oc8051_golden_model_1.SP [1], _27853_);
  dff (\oc8051_golden_model_1.SP [2], _27854_);
  dff (\oc8051_golden_model_1.SP [3], _27855_);
  dff (\oc8051_golden_model_1.SP [4], _27856_);
  dff (\oc8051_golden_model_1.SP [5], _27857_);
  dff (\oc8051_golden_model_1.SP [6], _27858_);
  dff (\oc8051_golden_model_1.SP [7], _25318_);
  dff (\oc8051_golden_model_1.TCON [0], _27861_);
  dff (\oc8051_golden_model_1.TCON [1], _27862_);
  dff (\oc8051_golden_model_1.TCON [2], _27863_);
  dff (\oc8051_golden_model_1.TCON [3], _27864_);
  dff (\oc8051_golden_model_1.TCON [4], _27865_);
  dff (\oc8051_golden_model_1.TCON [5], _27866_);
  dff (\oc8051_golden_model_1.TCON [6], _27868_);
  dff (\oc8051_golden_model_1.TCON [7], _25317_);
  dff (\oc8051_golden_model_1.TH0 [0], _27869_);
  dff (\oc8051_golden_model_1.TH0 [1], _27870_);
  dff (\oc8051_golden_model_1.TH0 [2], _27871_);
  dff (\oc8051_golden_model_1.TH0 [3], _27872_);
  dff (\oc8051_golden_model_1.TH0 [4], _27873_);
  dff (\oc8051_golden_model_1.TH0 [5], _27874_);
  dff (\oc8051_golden_model_1.TH0 [6], _27875_);
  dff (\oc8051_golden_model_1.TH0 [7], _25315_);
  dff (\oc8051_golden_model_1.TH1 [0], _27878_);
  dff (\oc8051_golden_model_1.TH1 [1], _27879_);
  dff (\oc8051_golden_model_1.TH1 [2], _27880_);
  dff (\oc8051_golden_model_1.TH1 [3], _27881_);
  dff (\oc8051_golden_model_1.TH1 [4], _27882_);
  dff (\oc8051_golden_model_1.TH1 [5], _27883_);
  dff (\oc8051_golden_model_1.TH1 [6], _27884_);
  dff (\oc8051_golden_model_1.TH1 [7], _25314_);
  dff (\oc8051_golden_model_1.TL0 [0], _27887_);
  dff (\oc8051_golden_model_1.TL0 [1], _27888_);
  dff (\oc8051_golden_model_1.TL0 [2], _27889_);
  dff (\oc8051_golden_model_1.TL0 [3], _27890_);
  dff (\oc8051_golden_model_1.TL0 [4], _27891_);
  dff (\oc8051_golden_model_1.TL0 [5], _27892_);
  dff (\oc8051_golden_model_1.TL0 [6], _27893_);
  dff (\oc8051_golden_model_1.TL0 [7], _25313_);
  dff (\oc8051_golden_model_1.TL1 [0], _27896_);
  dff (\oc8051_golden_model_1.TL1 [1], _27897_);
  dff (\oc8051_golden_model_1.TL1 [2], _27898_);
  dff (\oc8051_golden_model_1.TL1 [3], _27899_);
  dff (\oc8051_golden_model_1.TL1 [4], _27900_);
  dff (\oc8051_golden_model_1.TL1 [5], _27901_);
  dff (\oc8051_golden_model_1.TL1 [6], _27902_);
  dff (\oc8051_golden_model_1.TL1 [7], _25312_);
  dff (\oc8051_golden_model_1.TMOD [0], _27905_);
  dff (\oc8051_golden_model_1.TMOD [1], _27906_);
  dff (\oc8051_golden_model_1.TMOD [2], _27907_);
  dff (\oc8051_golden_model_1.TMOD [3], _27908_);
  dff (\oc8051_golden_model_1.TMOD [4], _27909_);
  dff (\oc8051_golden_model_1.TMOD [5], _27910_);
  dff (\oc8051_golden_model_1.TMOD [6], _27911_);
  dff (\oc8051_golden_model_1.TMOD [7], _25310_);
  dff (\oc8051_golden_model_1.PC [0], _27914_);
  dff (\oc8051_golden_model_1.PC [1], _27915_);
  dff (\oc8051_golden_model_1.PC [2], _27916_);
  dff (\oc8051_golden_model_1.PC [3], _27917_);
  dff (\oc8051_golden_model_1.PC [4], _27920_);
  dff (\oc8051_golden_model_1.PC [5], _27921_);
  dff (\oc8051_golden_model_1.PC [6], _27922_);
  dff (\oc8051_golden_model_1.PC [7], _27923_);
  dff (\oc8051_golden_model_1.PC [8], _27924_);
  dff (\oc8051_golden_model_1.PC [9], _27925_);
  dff (\oc8051_golden_model_1.PC [10], _27926_);
  dff (\oc8051_golden_model_1.PC [11], _27927_);
  dff (\oc8051_golden_model_1.PC [12], _27928_);
  dff (\oc8051_golden_model_1.PC [13], _27929_);
  dff (\oc8051_golden_model_1.PC [14], _27930_);
  dff (\oc8051_golden_model_1.PC [15], _25309_);
  dff (\oc8051_golden_model_1.P0INREG [0], _27931_);
  dff (\oc8051_golden_model_1.P0INREG [1], _27932_);
  dff (\oc8051_golden_model_1.P0INREG [2], _27935_);
  dff (\oc8051_golden_model_1.P0INREG [3], _27936_);
  dff (\oc8051_golden_model_1.P0INREG [4], _27937_);
  dff (\oc8051_golden_model_1.P0INREG [5], _27938_);
  dff (\oc8051_golden_model_1.P0INREG [6], _27939_);
  dff (\oc8051_golden_model_1.P0INREG [7], _25307_);
  dff (\oc8051_golden_model_1.P1INREG [0], _27942_);
  dff (\oc8051_golden_model_1.P1INREG [1], _27943_);
  dff (\oc8051_golden_model_1.P1INREG [2], _27944_);
  dff (\oc8051_golden_model_1.P1INREG [3], _27945_);
  dff (\oc8051_golden_model_1.P1INREG [4], _27946_);
  dff (\oc8051_golden_model_1.P1INREG [5], _27947_);
  dff (\oc8051_golden_model_1.P1INREG [6], _27948_);
  dff (\oc8051_golden_model_1.P1INREG [7], _25306_);
  dff (\oc8051_golden_model_1.P2INREG [0], _27949_);
  dff (\oc8051_golden_model_1.P2INREG [1], _27950_);
  dff (\oc8051_golden_model_1.P2INREG [2], _27951_);
  dff (\oc8051_golden_model_1.P2INREG [3], _27952_);
  dff (\oc8051_golden_model_1.P2INREG [4], _27955_);
  dff (\oc8051_golden_model_1.P2INREG [5], _27956_);
  dff (\oc8051_golden_model_1.P2INREG [6], _27957_);
  dff (\oc8051_golden_model_1.P2INREG [7], _25304_);
  dff (\oc8051_golden_model_1.P3INREG [0], _27960_);
  dff (\oc8051_golden_model_1.P3INREG [1], _27961_);
  dff (\oc8051_golden_model_1.P3INREG [2], _27962_);
  dff (\oc8051_golden_model_1.P3INREG [3], _27963_);
  dff (\oc8051_golden_model_1.P3INREG [4], _27964_);
  dff (\oc8051_golden_model_1.P3INREG [5], _27965_);
  dff (\oc8051_golden_model_1.P3INREG [6], _27966_);
  dff (\oc8051_golden_model_1.P3INREG [7], _25303_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _01047_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _01050_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _01053_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _01056_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _01058_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _01061_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _01064_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _00918_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _01067_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _01070_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _01073_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _01076_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _01079_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _01082_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _01085_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _00922_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _01088_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _01091_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _01094_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _01097_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _01100_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _01103_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _01105_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _00926_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _12208_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _12210_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _12124_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _12213_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _12216_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _12127_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _12219_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _12130_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _12222_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _12225_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _12228_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _12231_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _12234_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _12237_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _12240_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _12133_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _12136_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _24286_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _12139_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _24287_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _12142_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _24288_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _24289_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _12145_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _24290_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _24291_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _12148_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _24292_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _12151_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _24293_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _24294_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _24295_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _12154_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _24297_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _12157_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _12160_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _08192_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _03626_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _03628_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _03630_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _03632_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _03634_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _03636_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _03638_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _03640_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _03642_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _03644_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _03646_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _03648_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _03650_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _03652_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _03654_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _02771_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _03686_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _03688_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _03690_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _03692_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _03694_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _03696_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _03698_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _03700_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _03702_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _03704_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _03706_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _03708_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _03710_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _03712_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _03714_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _02775_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _05586_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _05588_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _05590_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _05592_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _05594_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _05596_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _05598_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _05600_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _05602_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _05604_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _05606_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _05608_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _05610_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _05612_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _05614_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _05616_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _05618_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _05620_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _05622_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _05624_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _05626_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _05628_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _05630_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _05632_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _05634_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _05636_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _05638_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _05640_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _05642_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _05644_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _05646_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _03224_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _03153_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _05649_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _05652_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _05655_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _05657_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _03160_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _05660_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _05663_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _05666_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _05669_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _05672_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _05675_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _05678_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _03164_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _05680_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _05682_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _05684_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _05686_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _05688_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _05690_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _05692_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _03167_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _05694_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _05696_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _05698_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _05700_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _05702_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _05704_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _05706_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _03170_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _03173_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _03177_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _05708_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _05710_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _05712_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _05714_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _05716_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _05718_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _05720_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _03180_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _05722_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _05724_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _05726_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _05728_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _05730_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _05732_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _05734_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _05736_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _05738_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _05740_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _05742_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _05744_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _05746_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _05748_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _05750_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _03183_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _05752_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _05754_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _05756_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _05758_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _05760_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _05762_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _05764_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _05766_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _05768_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _05770_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _05772_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _05774_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _05775_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _05777_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _05779_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _03186_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _03191_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _03197_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _03194_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _05781_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _05783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _05785_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _05787_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _05789_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _05791_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _05793_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _03200_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _05795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _05797_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _03202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _05799_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _05801_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _05803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _05805_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _05807_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _05809_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _05811_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _03204_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _05813_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _05815_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _05817_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _05819_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _05821_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _05823_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _05825_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _03207_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _03210_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _05827_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _05829_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _05831_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _05833_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _05835_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _05837_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _05839_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _03212_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _03215_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _03218_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _05841_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _05843_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _05845_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _03221_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _05847_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _05849_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _05851_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _05853_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _05855_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _05857_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _05859_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _05861_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _05863_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _05865_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _05867_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _05869_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _05871_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _05873_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _05875_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _05877_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _05879_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _05881_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _05883_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _05885_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _05887_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _05889_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _05891_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _05893_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _05895_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _05897_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _05899_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _05901_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _05903_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _05905_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _05907_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _03226_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _05909_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _05911_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _05913_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _05915_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _05917_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _05919_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _05921_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _03228_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _03230_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _03232_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _05923_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _05925_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _05927_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _05929_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _05931_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _05933_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _05935_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _05937_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _05938_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _05940_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _05942_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _05944_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _05946_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _05948_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _05950_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _03234_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _03236_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _03238_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _03240_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _05952_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _05954_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _05956_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _05958_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _05960_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _05962_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _05964_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _05966_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _05968_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _05970_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _05972_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _05974_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _05976_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _05978_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _05980_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _03242_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _03244_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _08290_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _08451_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _08453_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _08455_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _08457_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _08459_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _08461_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _08463_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _08293_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _08296_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _08465_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _08467_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _08298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _27382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _27388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _27394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _27400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _27406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _27412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _27418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _27421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _27464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _27468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _27472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _27476_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _27480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _27484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _27488_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _27491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _27429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _27433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _27437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _27441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _27445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _27449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _27453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _27456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _27532_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _27536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _27540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _27544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _27548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _27552_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _27556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _27559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _27497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _27501_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _27505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _27509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _27513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _27517_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _27521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _27524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _27694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _27698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _27702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _27706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _27710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _27714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _27718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _27728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _27662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _27666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _27670_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _27674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _27678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _27682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _27686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _27689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _27627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _27631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _27635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _27639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _27643_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _27647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _27651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _27654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _27596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _27600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _27604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _27608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _27612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _27616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _27619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _27622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _27564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _27568_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _27572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _27576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _27580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _27584_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _27588_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _27591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _28077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _28081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _28085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _28089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _28093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _28097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _28101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _27105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _28045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _28049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _28053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _28057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _28061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _28065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _28069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _28072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _28013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _28017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _28021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _28025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _28029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _28033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _28037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _28040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _27981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _27985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _27989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _27993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _27997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _28001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _28005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _28008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _27877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _27895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _27913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _27934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _27954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _27968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _27972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _27975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _27747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _27763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _27776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _27794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _27805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _27822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _27841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _27851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _00046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _00048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _00050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _00052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _00054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _00056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _00058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _27093_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _01520_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _01522_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _02203_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _02205_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _02207_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _02209_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _02211_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _02213_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _02215_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _01524_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _01527_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _08851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _08862_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _08873_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _08884_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _08895_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _08906_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _08917_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _07142_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _23586_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _23596_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _23606_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _23617_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _23627_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _23637_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _23647_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _05323_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _28332_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _28341_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _28349_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _28358_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _28367_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _28376_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _28384_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _27135_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _28393_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _28401_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _28410_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _28418_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _28427_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _28435_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _28444_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _27155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _25964_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _26952_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _26954_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _26956_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _26958_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _26960_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _26962_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _26964_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _25967_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _26966_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _25969_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _25972_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _26968_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _26970_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _25975_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _26972_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _26974_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _25978_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _26976_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _25979_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _26978_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _25981_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _26016_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _26018_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _26020_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _26022_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _26980_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _26982_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _26984_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _26024_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _26986_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _26988_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _26990_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _26991_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _26993_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _26995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _26997_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _26027_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _26999_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _27001_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _27003_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _27005_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _27007_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _27009_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _27011_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _26028_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _25391_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _25393_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _25395_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _25397_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _25399_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _25401_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _25403_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _19486_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _25405_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _25407_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _25409_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _25411_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _25413_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _25415_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _25417_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _19509_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _25419_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _25421_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _25423_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _25425_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _25427_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _25429_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _25431_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _19532_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _25433_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _25435_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _25437_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _25439_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _25441_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _25443_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _25445_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _19555_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _06381_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _06392_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _06403_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _06414_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _06425_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _06436_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _01600_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _25125_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _25133_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _25141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _25149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _25156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _25164_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _25175_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _24137_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _24117_);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.cy_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in , ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in , ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], 1'b0);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], 1'b0);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.desAc , ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_sfr1.desOv , ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [8], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [9], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [10], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [11], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [12], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [13], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [14], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [15], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_data_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_comp1.des [0], ABINPUT[27]);
  buf(\oc8051_top_1.oc8051_comp1.des [1], ABINPUT[28]);
  buf(\oc8051_top_1.oc8051_comp1.des [2], ABINPUT[29]);
  buf(\oc8051_top_1.oc8051_comp1.des [3], ABINPUT[30]);
  buf(\oc8051_top_1.oc8051_comp1.des [4], ABINPUT[31]);
  buf(\oc8051_top_1.oc8051_comp1.des [5], ABINPUT[32]);
  buf(\oc8051_top_1.oc8051_comp1.des [6], ABINPUT[33]);
  buf(\oc8051_top_1.oc8051_comp1.des [7], ABINPUT[34]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.PSW_next [0], ABINPUT008[0]);
  buf(\oc8051_golden_model_1.PSW_next [1], ABINPUT008[1]);
  buf(\oc8051_golden_model_1.PSW_next [2], ABINPUT008[2]);
  buf(\oc8051_golden_model_1.PSW_next [3], ABINPUT008[3]);
  buf(\oc8051_golden_model_1.PSW_next [4], ABINPUT008[4]);
  buf(\oc8051_golden_model_1.PSW_next [5], ABINPUT008[5]);
  buf(\oc8051_golden_model_1.PSW_next [6], ABINPUT008[6]);
  buf(\oc8051_golden_model_1.PSW_next [7], ABINPUT008[7]);
  buf(\oc8051_golden_model_1.ABINPUT007 [0], ABINPUT008[0]);
  buf(\oc8051_golden_model_1.ABINPUT007 [1], ABINPUT008[1]);
  buf(\oc8051_golden_model_1.ABINPUT007 [2], ABINPUT008[2]);
  buf(\oc8051_golden_model_1.ABINPUT007 [3], ABINPUT008[3]);
  buf(\oc8051_golden_model_1.ABINPUT007 [4], ABINPUT008[4]);
  buf(\oc8051_golden_model_1.ABINPUT007 [5], ABINPUT008[5]);
  buf(\oc8051_golden_model_1.ABINPUT007 [6], ABINPUT008[6]);
  buf(\oc8051_golden_model_1.ABINPUT007 [7], ABINPUT008[7]);
  buf(\oc8051_golden_model_1.P2_next [0], ABINPUT006[0]);
  buf(\oc8051_golden_model_1.P2_next [1], ABINPUT006[1]);
  buf(\oc8051_golden_model_1.P2_next [2], ABINPUT006[2]);
  buf(\oc8051_golden_model_1.P2_next [3], ABINPUT006[3]);
  buf(\oc8051_golden_model_1.P2_next [4], ABINPUT006[4]);
  buf(\oc8051_golden_model_1.P2_next [5], ABINPUT006[5]);
  buf(\oc8051_golden_model_1.P2_next [6], ABINPUT006[6]);
  buf(\oc8051_golden_model_1.P2_next [7], ABINPUT006[7]);
  buf(\oc8051_golden_model_1.ABINPUT005 [0], ABINPUT006[0]);
  buf(\oc8051_golden_model_1.ABINPUT005 [1], ABINPUT006[1]);
  buf(\oc8051_golden_model_1.ABINPUT005 [2], ABINPUT006[2]);
  buf(\oc8051_golden_model_1.ABINPUT005 [3], ABINPUT006[3]);
  buf(\oc8051_golden_model_1.ABINPUT005 [4], ABINPUT006[4]);
  buf(\oc8051_golden_model_1.ABINPUT005 [5], ABINPUT006[5]);
  buf(\oc8051_golden_model_1.ABINPUT005 [6], ABINPUT006[6]);
  buf(\oc8051_golden_model_1.ABINPUT005 [7], ABINPUT006[7]);
  buf(\oc8051_golden_model_1.P0_next [0], ABINPUT004[0]);
  buf(\oc8051_golden_model_1.P0_next [1], ABINPUT004[1]);
  buf(\oc8051_golden_model_1.P0_next [2], ABINPUT004[2]);
  buf(\oc8051_golden_model_1.P0_next [3], ABINPUT004[3]);
  buf(\oc8051_golden_model_1.P0_next [4], ABINPUT004[4]);
  buf(\oc8051_golden_model_1.P0_next [5], ABINPUT004[5]);
  buf(\oc8051_golden_model_1.P0_next [6], ABINPUT004[6]);
  buf(\oc8051_golden_model_1.P0_next [7], ABINPUT004[7]);
  buf(\oc8051_golden_model_1.ABINPUT003 [0], ABINPUT004[0]);
  buf(\oc8051_golden_model_1.ABINPUT003 [1], ABINPUT004[1]);
  buf(\oc8051_golden_model_1.ABINPUT003 [2], ABINPUT004[2]);
  buf(\oc8051_golden_model_1.ABINPUT003 [3], ABINPUT004[3]);
  buf(\oc8051_golden_model_1.ABINPUT003 [4], ABINPUT004[4]);
  buf(\oc8051_golden_model_1.ABINPUT003 [5], ABINPUT004[5]);
  buf(\oc8051_golden_model_1.ABINPUT003 [6], ABINPUT004[6]);
  buf(\oc8051_golden_model_1.ABINPUT003 [7], ABINPUT004[7]);
  buf(\oc8051_golden_model_1.DPL_next [0], ABINPUT002[0]);
  buf(\oc8051_golden_model_1.DPL_next [1], ABINPUT002[1]);
  buf(\oc8051_golden_model_1.DPL_next [2], ABINPUT002[2]);
  buf(\oc8051_golden_model_1.DPL_next [3], ABINPUT002[3]);
  buf(\oc8051_golden_model_1.DPL_next [4], ABINPUT002[4]);
  buf(\oc8051_golden_model_1.DPL_next [5], ABINPUT002[5]);
  buf(\oc8051_golden_model_1.DPL_next [6], ABINPUT002[6]);
  buf(\oc8051_golden_model_1.DPL_next [7], ABINPUT002[7]);
  buf(\oc8051_golden_model_1.ABINPUT001 [0], ABINPUT002[0]);
  buf(\oc8051_golden_model_1.ABINPUT001 [1], ABINPUT002[1]);
  buf(\oc8051_golden_model_1.ABINPUT001 [2], ABINPUT002[2]);
  buf(\oc8051_golden_model_1.ABINPUT001 [3], ABINPUT002[3]);
  buf(\oc8051_golden_model_1.ABINPUT001 [4], ABINPUT002[4]);
  buf(\oc8051_golden_model_1.ABINPUT001 [5], ABINPUT002[5]);
  buf(\oc8051_golden_model_1.ABINPUT001 [6], ABINPUT002[6]);
  buf(\oc8051_golden_model_1.ABINPUT001 [7], ABINPUT002[7]);
  buf(\oc8051_golden_model_1.ACC_next [0], ABINPUT000[0]);
  buf(\oc8051_golden_model_1.ACC_next [1], ABINPUT000[1]);
  buf(\oc8051_golden_model_1.ACC_next [2], ABINPUT000[2]);
  buf(\oc8051_golden_model_1.ACC_next [3], ABINPUT000[3]);
  buf(\oc8051_golden_model_1.ACC_next [4], ABINPUT000[4]);
  buf(\oc8051_golden_model_1.ACC_next [5], ABINPUT000[5]);
  buf(\oc8051_golden_model_1.ACC_next [6], ABINPUT000[6]);
  buf(\oc8051_golden_model_1.ACC_next [7], ABINPUT000[7]);
  buf(\oc8051_golden_model_1.ABINPUT [0], ABINPUT000[0]);
  buf(\oc8051_golden_model_1.ABINPUT [1], ABINPUT000[1]);
  buf(\oc8051_golden_model_1.ABINPUT [2], ABINPUT000[2]);
  buf(\oc8051_golden_model_1.ABINPUT [3], ABINPUT000[3]);
  buf(\oc8051_golden_model_1.ABINPUT [4], ABINPUT000[4]);
  buf(\oc8051_golden_model_1.ABINPUT [5], ABINPUT000[5]);
  buf(\oc8051_golden_model_1.ABINPUT [6], ABINPUT000[6]);
  buf(\oc8051_golden_model_1.ABINPUT [7], ABINPUT000[7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e6 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.ACC_e6 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.ACC_e6 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.ACC_e6 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.ACC_e6 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.ACC_e6 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.ACC_e6 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.ACC_e6 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.ACC_e7 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.ACC_e7 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.ACC_e7 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.ACC_e7 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.ACC_e7 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.ACC_e7 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.ACC_e7 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.ACC_e7 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n2854 [0], \oc8051_golden_model_1.PSW_d4 [0]);
  buf(\oc8051_golden_model_1.n2854 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2854 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2854 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2854 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2854 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2854 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2854 [7], \oc8051_golden_model_1.n2838 [6]);
  buf(\oc8051_golden_model_1.n2858 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n2858 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n2858 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n2858 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n2858 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2858 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2858 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2858 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2859 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n2859 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n2859 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n2859 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n2860 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2860 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2860 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2860 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2860 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n2860 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n2860 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n2860 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n2861 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2862 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2863 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2864 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2865 , \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n2866 , \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n2441 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2867 , \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n2868 , \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.IRAM_full [0], ABINPUT009[0]);
  buf(\oc8051_golden_model_1.IRAM_full [1], ABINPUT009[1]);
  buf(\oc8051_golden_model_1.IRAM_full [2], ABINPUT009[2]);
  buf(\oc8051_golden_model_1.IRAM_full [3], ABINPUT009[3]);
  buf(\oc8051_golden_model_1.IRAM_full [4], ABINPUT009[4]);
  buf(\oc8051_golden_model_1.IRAM_full [5], ABINPUT009[5]);
  buf(\oc8051_golden_model_1.IRAM_full [6], ABINPUT009[6]);
  buf(\oc8051_golden_model_1.IRAM_full [7], ABINPUT009[7]);
  buf(\oc8051_golden_model_1.IRAM_full [8], ABINPUT009[8]);
  buf(\oc8051_golden_model_1.IRAM_full [9], ABINPUT009[9]);
  buf(\oc8051_golden_model_1.IRAM_full [10], ABINPUT009[10]);
  buf(\oc8051_golden_model_1.IRAM_full [11], ABINPUT009[11]);
  buf(\oc8051_golden_model_1.IRAM_full [12], ABINPUT009[12]);
  buf(\oc8051_golden_model_1.IRAM_full [13], ABINPUT009[13]);
  buf(\oc8051_golden_model_1.IRAM_full [14], ABINPUT009[14]);
  buf(\oc8051_golden_model_1.IRAM_full [15], ABINPUT009[15]);
  buf(\oc8051_golden_model_1.IRAM_full [16], ABINPUT009[16]);
  buf(\oc8051_golden_model_1.IRAM_full [17], ABINPUT009[17]);
  buf(\oc8051_golden_model_1.IRAM_full [18], ABINPUT009[18]);
  buf(\oc8051_golden_model_1.IRAM_full [19], ABINPUT009[19]);
  buf(\oc8051_golden_model_1.IRAM_full [20], ABINPUT009[20]);
  buf(\oc8051_golden_model_1.IRAM_full [21], ABINPUT009[21]);
  buf(\oc8051_golden_model_1.IRAM_full [22], ABINPUT009[22]);
  buf(\oc8051_golden_model_1.IRAM_full [23], ABINPUT009[23]);
  buf(\oc8051_golden_model_1.IRAM_full [24], ABINPUT009[24]);
  buf(\oc8051_golden_model_1.IRAM_full [25], ABINPUT009[25]);
  buf(\oc8051_golden_model_1.IRAM_full [26], ABINPUT009[26]);
  buf(\oc8051_golden_model_1.IRAM_full [27], ABINPUT009[27]);
  buf(\oc8051_golden_model_1.IRAM_full [28], ABINPUT009[28]);
  buf(\oc8051_golden_model_1.IRAM_full [29], ABINPUT009[29]);
  buf(\oc8051_golden_model_1.IRAM_full [30], ABINPUT009[30]);
  buf(\oc8051_golden_model_1.IRAM_full [31], ABINPUT009[31]);
  buf(\oc8051_golden_model_1.IRAM_full [32], ABINPUT009[32]);
  buf(\oc8051_golden_model_1.IRAM_full [33], ABINPUT009[33]);
  buf(\oc8051_golden_model_1.IRAM_full [34], ABINPUT009[34]);
  buf(\oc8051_golden_model_1.IRAM_full [35], ABINPUT009[35]);
  buf(\oc8051_golden_model_1.IRAM_full [36], ABINPUT009[36]);
  buf(\oc8051_golden_model_1.IRAM_full [37], ABINPUT009[37]);
  buf(\oc8051_golden_model_1.IRAM_full [38], ABINPUT009[38]);
  buf(\oc8051_golden_model_1.IRAM_full [39], ABINPUT009[39]);
  buf(\oc8051_golden_model_1.IRAM_full [40], ABINPUT009[40]);
  buf(\oc8051_golden_model_1.IRAM_full [41], ABINPUT009[41]);
  buf(\oc8051_golden_model_1.IRAM_full [42], ABINPUT009[42]);
  buf(\oc8051_golden_model_1.IRAM_full [43], ABINPUT009[43]);
  buf(\oc8051_golden_model_1.IRAM_full [44], ABINPUT009[44]);
  buf(\oc8051_golden_model_1.IRAM_full [45], ABINPUT009[45]);
  buf(\oc8051_golden_model_1.IRAM_full [46], ABINPUT009[46]);
  buf(\oc8051_golden_model_1.IRAM_full [47], ABINPUT009[47]);
  buf(\oc8051_golden_model_1.IRAM_full [48], ABINPUT009[48]);
  buf(\oc8051_golden_model_1.IRAM_full [49], ABINPUT009[49]);
  buf(\oc8051_golden_model_1.IRAM_full [50], ABINPUT009[50]);
  buf(\oc8051_golden_model_1.IRAM_full [51], ABINPUT009[51]);
  buf(\oc8051_golden_model_1.IRAM_full [52], ABINPUT009[52]);
  buf(\oc8051_golden_model_1.IRAM_full [53], ABINPUT009[53]);
  buf(\oc8051_golden_model_1.IRAM_full [54], ABINPUT009[54]);
  buf(\oc8051_golden_model_1.IRAM_full [55], ABINPUT009[55]);
  buf(\oc8051_golden_model_1.IRAM_full [56], ABINPUT009[56]);
  buf(\oc8051_golden_model_1.IRAM_full [57], ABINPUT009[57]);
  buf(\oc8051_golden_model_1.IRAM_full [58], ABINPUT009[58]);
  buf(\oc8051_golden_model_1.IRAM_full [59], ABINPUT009[59]);
  buf(\oc8051_golden_model_1.IRAM_full [60], ABINPUT009[60]);
  buf(\oc8051_golden_model_1.IRAM_full [61], ABINPUT009[61]);
  buf(\oc8051_golden_model_1.IRAM_full [62], ABINPUT009[62]);
  buf(\oc8051_golden_model_1.IRAM_full [63], ABINPUT009[63]);
  buf(\oc8051_golden_model_1.IRAM_full [64], ABINPUT009[64]);
  buf(\oc8051_golden_model_1.IRAM_full [65], ABINPUT009[65]);
  buf(\oc8051_golden_model_1.IRAM_full [66], ABINPUT009[66]);
  buf(\oc8051_golden_model_1.IRAM_full [67], ABINPUT009[67]);
  buf(\oc8051_golden_model_1.IRAM_full [68], ABINPUT009[68]);
  buf(\oc8051_golden_model_1.IRAM_full [69], ABINPUT009[69]);
  buf(\oc8051_golden_model_1.IRAM_full [70], ABINPUT009[70]);
  buf(\oc8051_golden_model_1.IRAM_full [71], ABINPUT009[71]);
  buf(\oc8051_golden_model_1.IRAM_full [72], ABINPUT009[72]);
  buf(\oc8051_golden_model_1.IRAM_full [73], ABINPUT009[73]);
  buf(\oc8051_golden_model_1.IRAM_full [74], ABINPUT009[74]);
  buf(\oc8051_golden_model_1.IRAM_full [75], ABINPUT009[75]);
  buf(\oc8051_golden_model_1.IRAM_full [76], ABINPUT009[76]);
  buf(\oc8051_golden_model_1.IRAM_full [77], ABINPUT009[77]);
  buf(\oc8051_golden_model_1.IRAM_full [78], ABINPUT009[78]);
  buf(\oc8051_golden_model_1.IRAM_full [79], ABINPUT009[79]);
  buf(\oc8051_golden_model_1.IRAM_full [80], ABINPUT009[80]);
  buf(\oc8051_golden_model_1.IRAM_full [81], ABINPUT009[81]);
  buf(\oc8051_golden_model_1.IRAM_full [82], ABINPUT009[82]);
  buf(\oc8051_golden_model_1.IRAM_full [83], ABINPUT009[83]);
  buf(\oc8051_golden_model_1.IRAM_full [84], ABINPUT009[84]);
  buf(\oc8051_golden_model_1.IRAM_full [85], ABINPUT009[85]);
  buf(\oc8051_golden_model_1.IRAM_full [86], ABINPUT009[86]);
  buf(\oc8051_golden_model_1.IRAM_full [87], ABINPUT009[87]);
  buf(\oc8051_golden_model_1.IRAM_full [88], ABINPUT009[88]);
  buf(\oc8051_golden_model_1.IRAM_full [89], ABINPUT009[89]);
  buf(\oc8051_golden_model_1.IRAM_full [90], ABINPUT009[90]);
  buf(\oc8051_golden_model_1.IRAM_full [91], ABINPUT009[91]);
  buf(\oc8051_golden_model_1.IRAM_full [92], ABINPUT009[92]);
  buf(\oc8051_golden_model_1.IRAM_full [93], ABINPUT009[93]);
  buf(\oc8051_golden_model_1.IRAM_full [94], ABINPUT009[94]);
  buf(\oc8051_golden_model_1.IRAM_full [95], ABINPUT009[95]);
  buf(\oc8051_golden_model_1.IRAM_full [96], ABINPUT009[96]);
  buf(\oc8051_golden_model_1.IRAM_full [97], ABINPUT009[97]);
  buf(\oc8051_golden_model_1.IRAM_full [98], ABINPUT009[98]);
  buf(\oc8051_golden_model_1.IRAM_full [99], ABINPUT009[99]);
  buf(\oc8051_golden_model_1.IRAM_full [100], ABINPUT009[100]);
  buf(\oc8051_golden_model_1.IRAM_full [101], ABINPUT009[101]);
  buf(\oc8051_golden_model_1.IRAM_full [102], ABINPUT009[102]);
  buf(\oc8051_golden_model_1.IRAM_full [103], ABINPUT009[103]);
  buf(\oc8051_golden_model_1.IRAM_full [104], ABINPUT009[104]);
  buf(\oc8051_golden_model_1.IRAM_full [105], ABINPUT009[105]);
  buf(\oc8051_golden_model_1.IRAM_full [106], ABINPUT009[106]);
  buf(\oc8051_golden_model_1.IRAM_full [107], ABINPUT009[107]);
  buf(\oc8051_golden_model_1.IRAM_full [108], ABINPUT009[108]);
  buf(\oc8051_golden_model_1.IRAM_full [109], ABINPUT009[109]);
  buf(\oc8051_golden_model_1.IRAM_full [110], ABINPUT009[110]);
  buf(\oc8051_golden_model_1.IRAM_full [111], ABINPUT009[111]);
  buf(\oc8051_golden_model_1.IRAM_full [112], ABINPUT009[112]);
  buf(\oc8051_golden_model_1.IRAM_full [113], ABINPUT009[113]);
  buf(\oc8051_golden_model_1.IRAM_full [114], ABINPUT009[114]);
  buf(\oc8051_golden_model_1.IRAM_full [115], ABINPUT009[115]);
  buf(\oc8051_golden_model_1.IRAM_full [116], ABINPUT009[116]);
  buf(\oc8051_golden_model_1.IRAM_full [117], ABINPUT009[117]);
  buf(\oc8051_golden_model_1.IRAM_full [118], ABINPUT009[118]);
  buf(\oc8051_golden_model_1.IRAM_full [119], ABINPUT009[119]);
  buf(\oc8051_golden_model_1.IRAM_full [120], ABINPUT009[120]);
  buf(\oc8051_golden_model_1.IRAM_full [121], ABINPUT009[121]);
  buf(\oc8051_golden_model_1.IRAM_full [122], ABINPUT009[122]);
  buf(\oc8051_golden_model_1.IRAM_full [123], ABINPUT009[123]);
  buf(\oc8051_golden_model_1.IRAM_full [124], ABINPUT009[124]);
  buf(\oc8051_golden_model_1.IRAM_full [125], ABINPUT009[125]);
  buf(\oc8051_golden_model_1.IRAM_full [126], ABINPUT009[126]);
  buf(\oc8051_golden_model_1.IRAM_full [127], ABINPUT009[127]);
  buf(\oc8051_golden_model_1.ABINPUT008 [0], ABINPUT009[0]);
  buf(\oc8051_golden_model_1.ABINPUT008 [1], ABINPUT009[1]);
  buf(\oc8051_golden_model_1.ABINPUT008 [2], ABINPUT009[2]);
  buf(\oc8051_golden_model_1.ABINPUT008 [3], ABINPUT009[3]);
  buf(\oc8051_golden_model_1.ABINPUT008 [4], ABINPUT009[4]);
  buf(\oc8051_golden_model_1.ABINPUT008 [5], ABINPUT009[5]);
  buf(\oc8051_golden_model_1.ABINPUT008 [6], ABINPUT009[6]);
  buf(\oc8051_golden_model_1.ABINPUT008 [7], ABINPUT009[7]);
  buf(\oc8051_golden_model_1.ABINPUT008 [8], ABINPUT009[8]);
  buf(\oc8051_golden_model_1.ABINPUT008 [9], ABINPUT009[9]);
  buf(\oc8051_golden_model_1.ABINPUT008 [10], ABINPUT009[10]);
  buf(\oc8051_golden_model_1.ABINPUT008 [11], ABINPUT009[11]);
  buf(\oc8051_golden_model_1.ABINPUT008 [12], ABINPUT009[12]);
  buf(\oc8051_golden_model_1.ABINPUT008 [13], ABINPUT009[13]);
  buf(\oc8051_golden_model_1.ABINPUT008 [14], ABINPUT009[14]);
  buf(\oc8051_golden_model_1.ABINPUT008 [15], ABINPUT009[15]);
  buf(\oc8051_golden_model_1.ABINPUT008 [16], ABINPUT009[16]);
  buf(\oc8051_golden_model_1.ABINPUT008 [17], ABINPUT009[17]);
  buf(\oc8051_golden_model_1.ABINPUT008 [18], ABINPUT009[18]);
  buf(\oc8051_golden_model_1.ABINPUT008 [19], ABINPUT009[19]);
  buf(\oc8051_golden_model_1.ABINPUT008 [20], ABINPUT009[20]);
  buf(\oc8051_golden_model_1.ABINPUT008 [21], ABINPUT009[21]);
  buf(\oc8051_golden_model_1.ABINPUT008 [22], ABINPUT009[22]);
  buf(\oc8051_golden_model_1.ABINPUT008 [23], ABINPUT009[23]);
  buf(\oc8051_golden_model_1.ABINPUT008 [24], ABINPUT009[24]);
  buf(\oc8051_golden_model_1.ABINPUT008 [25], ABINPUT009[25]);
  buf(\oc8051_golden_model_1.ABINPUT008 [26], ABINPUT009[26]);
  buf(\oc8051_golden_model_1.ABINPUT008 [27], ABINPUT009[27]);
  buf(\oc8051_golden_model_1.ABINPUT008 [28], ABINPUT009[28]);
  buf(\oc8051_golden_model_1.ABINPUT008 [29], ABINPUT009[29]);
  buf(\oc8051_golden_model_1.ABINPUT008 [30], ABINPUT009[30]);
  buf(\oc8051_golden_model_1.ABINPUT008 [31], ABINPUT009[31]);
  buf(\oc8051_golden_model_1.ABINPUT008 [32], ABINPUT009[32]);
  buf(\oc8051_golden_model_1.ABINPUT008 [33], ABINPUT009[33]);
  buf(\oc8051_golden_model_1.ABINPUT008 [34], ABINPUT009[34]);
  buf(\oc8051_golden_model_1.ABINPUT008 [35], ABINPUT009[35]);
  buf(\oc8051_golden_model_1.ABINPUT008 [36], ABINPUT009[36]);
  buf(\oc8051_golden_model_1.ABINPUT008 [37], ABINPUT009[37]);
  buf(\oc8051_golden_model_1.ABINPUT008 [38], ABINPUT009[38]);
  buf(\oc8051_golden_model_1.ABINPUT008 [39], ABINPUT009[39]);
  buf(\oc8051_golden_model_1.ABINPUT008 [40], ABINPUT009[40]);
  buf(\oc8051_golden_model_1.ABINPUT008 [41], ABINPUT009[41]);
  buf(\oc8051_golden_model_1.ABINPUT008 [42], ABINPUT009[42]);
  buf(\oc8051_golden_model_1.ABINPUT008 [43], ABINPUT009[43]);
  buf(\oc8051_golden_model_1.ABINPUT008 [44], ABINPUT009[44]);
  buf(\oc8051_golden_model_1.ABINPUT008 [45], ABINPUT009[45]);
  buf(\oc8051_golden_model_1.ABINPUT008 [46], ABINPUT009[46]);
  buf(\oc8051_golden_model_1.ABINPUT008 [47], ABINPUT009[47]);
  buf(\oc8051_golden_model_1.ABINPUT008 [48], ABINPUT009[48]);
  buf(\oc8051_golden_model_1.ABINPUT008 [49], ABINPUT009[49]);
  buf(\oc8051_golden_model_1.ABINPUT008 [50], ABINPUT009[50]);
  buf(\oc8051_golden_model_1.ABINPUT008 [51], ABINPUT009[51]);
  buf(\oc8051_golden_model_1.ABINPUT008 [52], ABINPUT009[52]);
  buf(\oc8051_golden_model_1.ABINPUT008 [53], ABINPUT009[53]);
  buf(\oc8051_golden_model_1.ABINPUT008 [54], ABINPUT009[54]);
  buf(\oc8051_golden_model_1.ABINPUT008 [55], ABINPUT009[55]);
  buf(\oc8051_golden_model_1.ABINPUT008 [56], ABINPUT009[56]);
  buf(\oc8051_golden_model_1.ABINPUT008 [57], ABINPUT009[57]);
  buf(\oc8051_golden_model_1.ABINPUT008 [58], ABINPUT009[58]);
  buf(\oc8051_golden_model_1.ABINPUT008 [59], ABINPUT009[59]);
  buf(\oc8051_golden_model_1.ABINPUT008 [60], ABINPUT009[60]);
  buf(\oc8051_golden_model_1.ABINPUT008 [61], ABINPUT009[61]);
  buf(\oc8051_golden_model_1.ABINPUT008 [62], ABINPUT009[62]);
  buf(\oc8051_golden_model_1.ABINPUT008 [63], ABINPUT009[63]);
  buf(\oc8051_golden_model_1.ABINPUT008 [64], ABINPUT009[64]);
  buf(\oc8051_golden_model_1.ABINPUT008 [65], ABINPUT009[65]);
  buf(\oc8051_golden_model_1.ABINPUT008 [66], ABINPUT009[66]);
  buf(\oc8051_golden_model_1.ABINPUT008 [67], ABINPUT009[67]);
  buf(\oc8051_golden_model_1.ABINPUT008 [68], ABINPUT009[68]);
  buf(\oc8051_golden_model_1.ABINPUT008 [69], ABINPUT009[69]);
  buf(\oc8051_golden_model_1.ABINPUT008 [70], ABINPUT009[70]);
  buf(\oc8051_golden_model_1.ABINPUT008 [71], ABINPUT009[71]);
  buf(\oc8051_golden_model_1.ABINPUT008 [72], ABINPUT009[72]);
  buf(\oc8051_golden_model_1.ABINPUT008 [73], ABINPUT009[73]);
  buf(\oc8051_golden_model_1.ABINPUT008 [74], ABINPUT009[74]);
  buf(\oc8051_golden_model_1.ABINPUT008 [75], ABINPUT009[75]);
  buf(\oc8051_golden_model_1.ABINPUT008 [76], ABINPUT009[76]);
  buf(\oc8051_golden_model_1.ABINPUT008 [77], ABINPUT009[77]);
  buf(\oc8051_golden_model_1.ABINPUT008 [78], ABINPUT009[78]);
  buf(\oc8051_golden_model_1.ABINPUT008 [79], ABINPUT009[79]);
  buf(\oc8051_golden_model_1.ABINPUT008 [80], ABINPUT009[80]);
  buf(\oc8051_golden_model_1.ABINPUT008 [81], ABINPUT009[81]);
  buf(\oc8051_golden_model_1.ABINPUT008 [82], ABINPUT009[82]);
  buf(\oc8051_golden_model_1.ABINPUT008 [83], ABINPUT009[83]);
  buf(\oc8051_golden_model_1.ABINPUT008 [84], ABINPUT009[84]);
  buf(\oc8051_golden_model_1.ABINPUT008 [85], ABINPUT009[85]);
  buf(\oc8051_golden_model_1.ABINPUT008 [86], ABINPUT009[86]);
  buf(\oc8051_golden_model_1.ABINPUT008 [87], ABINPUT009[87]);
  buf(\oc8051_golden_model_1.ABINPUT008 [88], ABINPUT009[88]);
  buf(\oc8051_golden_model_1.ABINPUT008 [89], ABINPUT009[89]);
  buf(\oc8051_golden_model_1.ABINPUT008 [90], ABINPUT009[90]);
  buf(\oc8051_golden_model_1.ABINPUT008 [91], ABINPUT009[91]);
  buf(\oc8051_golden_model_1.ABINPUT008 [92], ABINPUT009[92]);
  buf(\oc8051_golden_model_1.ABINPUT008 [93], ABINPUT009[93]);
  buf(\oc8051_golden_model_1.ABINPUT008 [94], ABINPUT009[94]);
  buf(\oc8051_golden_model_1.ABINPUT008 [95], ABINPUT009[95]);
  buf(\oc8051_golden_model_1.ABINPUT008 [96], ABINPUT009[96]);
  buf(\oc8051_golden_model_1.ABINPUT008 [97], ABINPUT009[97]);
  buf(\oc8051_golden_model_1.ABINPUT008 [98], ABINPUT009[98]);
  buf(\oc8051_golden_model_1.ABINPUT008 [99], ABINPUT009[99]);
  buf(\oc8051_golden_model_1.ABINPUT008 [100], ABINPUT009[100]);
  buf(\oc8051_golden_model_1.ABINPUT008 [101], ABINPUT009[101]);
  buf(\oc8051_golden_model_1.ABINPUT008 [102], ABINPUT009[102]);
  buf(\oc8051_golden_model_1.ABINPUT008 [103], ABINPUT009[103]);
  buf(\oc8051_golden_model_1.ABINPUT008 [104], ABINPUT009[104]);
  buf(\oc8051_golden_model_1.ABINPUT008 [105], ABINPUT009[105]);
  buf(\oc8051_golden_model_1.ABINPUT008 [106], ABINPUT009[106]);
  buf(\oc8051_golden_model_1.ABINPUT008 [107], ABINPUT009[107]);
  buf(\oc8051_golden_model_1.ABINPUT008 [108], ABINPUT009[108]);
  buf(\oc8051_golden_model_1.ABINPUT008 [109], ABINPUT009[109]);
  buf(\oc8051_golden_model_1.ABINPUT008 [110], ABINPUT009[110]);
  buf(\oc8051_golden_model_1.ABINPUT008 [111], ABINPUT009[111]);
  buf(\oc8051_golden_model_1.ABINPUT008 [112], ABINPUT009[112]);
  buf(\oc8051_golden_model_1.ABINPUT008 [113], ABINPUT009[113]);
  buf(\oc8051_golden_model_1.ABINPUT008 [114], ABINPUT009[114]);
  buf(\oc8051_golden_model_1.ABINPUT008 [115], ABINPUT009[115]);
  buf(\oc8051_golden_model_1.ABINPUT008 [116], ABINPUT009[116]);
  buf(\oc8051_golden_model_1.ABINPUT008 [117], ABINPUT009[117]);
  buf(\oc8051_golden_model_1.ABINPUT008 [118], ABINPUT009[118]);
  buf(\oc8051_golden_model_1.ABINPUT008 [119], ABINPUT009[119]);
  buf(\oc8051_golden_model_1.ABINPUT008 [120], ABINPUT009[120]);
  buf(\oc8051_golden_model_1.ABINPUT008 [121], ABINPUT009[121]);
  buf(\oc8051_golden_model_1.ABINPUT008 [122], ABINPUT009[122]);
  buf(\oc8051_golden_model_1.ABINPUT008 [123], ABINPUT009[123]);
  buf(\oc8051_golden_model_1.ABINPUT008 [124], ABINPUT009[124]);
  buf(\oc8051_golden_model_1.ABINPUT008 [125], ABINPUT009[125]);
  buf(\oc8051_golden_model_1.ABINPUT008 [126], ABINPUT009[126]);
  buf(\oc8051_golden_model_1.ABINPUT008 [127], ABINPUT009[127]);
  buf(\oc8051_golden_model_1.P3_next [0], ABINPUT007[0]);
  buf(\oc8051_golden_model_1.P3_next [1], ABINPUT007[1]);
  buf(\oc8051_golden_model_1.P3_next [2], ABINPUT007[2]);
  buf(\oc8051_golden_model_1.P3_next [3], ABINPUT007[3]);
  buf(\oc8051_golden_model_1.P3_next [4], ABINPUT007[4]);
  buf(\oc8051_golden_model_1.P3_next [5], ABINPUT007[5]);
  buf(\oc8051_golden_model_1.P3_next [6], ABINPUT007[6]);
  buf(\oc8051_golden_model_1.P3_next [7], ABINPUT007[7]);
  buf(\oc8051_golden_model_1.ABINPUT006 [0], ABINPUT007[0]);
  buf(\oc8051_golden_model_1.ABINPUT006 [1], ABINPUT007[1]);
  buf(\oc8051_golden_model_1.ABINPUT006 [2], ABINPUT007[2]);
  buf(\oc8051_golden_model_1.ABINPUT006 [3], ABINPUT007[3]);
  buf(\oc8051_golden_model_1.ABINPUT006 [4], ABINPUT007[4]);
  buf(\oc8051_golden_model_1.ABINPUT006 [5], ABINPUT007[5]);
  buf(\oc8051_golden_model_1.ABINPUT006 [6], ABINPUT007[6]);
  buf(\oc8051_golden_model_1.ABINPUT006 [7], ABINPUT007[7]);
  buf(\oc8051_golden_model_1.P1_next [0], ABINPUT005[0]);
  buf(\oc8051_golden_model_1.P1_next [1], ABINPUT005[1]);
  buf(\oc8051_golden_model_1.P1_next [2], ABINPUT005[2]);
  buf(\oc8051_golden_model_1.P1_next [3], ABINPUT005[3]);
  buf(\oc8051_golden_model_1.P1_next [4], ABINPUT005[4]);
  buf(\oc8051_golden_model_1.P1_next [5], ABINPUT005[5]);
  buf(\oc8051_golden_model_1.P1_next [6], ABINPUT005[6]);
  buf(\oc8051_golden_model_1.P1_next [7], ABINPUT005[7]);
  buf(\oc8051_golden_model_1.ABINPUT004 [0], ABINPUT005[0]);
  buf(\oc8051_golden_model_1.ABINPUT004 [1], ABINPUT005[1]);
  buf(\oc8051_golden_model_1.ABINPUT004 [2], ABINPUT005[2]);
  buf(\oc8051_golden_model_1.ABINPUT004 [3], ABINPUT005[3]);
  buf(\oc8051_golden_model_1.ABINPUT004 [4], ABINPUT005[4]);
  buf(\oc8051_golden_model_1.ABINPUT004 [5], ABINPUT005[5]);
  buf(\oc8051_golden_model_1.ABINPUT004 [6], ABINPUT005[6]);
  buf(\oc8051_golden_model_1.ABINPUT004 [7], ABINPUT005[7]);
  buf(\oc8051_golden_model_1.DPH_next [0], ABINPUT003[0]);
  buf(\oc8051_golden_model_1.DPH_next [1], ABINPUT003[1]);
  buf(\oc8051_golden_model_1.DPH_next [2], ABINPUT003[2]);
  buf(\oc8051_golden_model_1.DPH_next [3], ABINPUT003[3]);
  buf(\oc8051_golden_model_1.DPH_next [4], ABINPUT003[4]);
  buf(\oc8051_golden_model_1.DPH_next [5], ABINPUT003[5]);
  buf(\oc8051_golden_model_1.DPH_next [6], ABINPUT003[6]);
  buf(\oc8051_golden_model_1.DPH_next [7], ABINPUT003[7]);
  buf(\oc8051_golden_model_1.ABINPUT002 [0], ABINPUT003[0]);
  buf(\oc8051_golden_model_1.ABINPUT002 [1], ABINPUT003[1]);
  buf(\oc8051_golden_model_1.ABINPUT002 [2], ABINPUT003[2]);
  buf(\oc8051_golden_model_1.ABINPUT002 [3], ABINPUT003[3]);
  buf(\oc8051_golden_model_1.ABINPUT002 [4], ABINPUT003[4]);
  buf(\oc8051_golden_model_1.ABINPUT002 [5], ABINPUT003[5]);
  buf(\oc8051_golden_model_1.ABINPUT002 [6], ABINPUT003[6]);
  buf(\oc8051_golden_model_1.ABINPUT002 [7], ABINPUT003[7]);
  buf(\oc8051_golden_model_1.B_next [0], ABINPUT001[0]);
  buf(\oc8051_golden_model_1.B_next [1], ABINPUT001[1]);
  buf(\oc8051_golden_model_1.B_next [2], ABINPUT001[2]);
  buf(\oc8051_golden_model_1.B_next [3], ABINPUT001[3]);
  buf(\oc8051_golden_model_1.B_next [4], ABINPUT001[4]);
  buf(\oc8051_golden_model_1.B_next [5], ABINPUT001[5]);
  buf(\oc8051_golden_model_1.B_next [6], ABINPUT001[6]);
  buf(\oc8051_golden_model_1.B_next [7], ABINPUT001[7]);
  buf(\oc8051_golden_model_1.ABINPUT000 [0], ABINPUT001[0]);
  buf(\oc8051_golden_model_1.ABINPUT000 [1], ABINPUT001[1]);
  buf(\oc8051_golden_model_1.ABINPUT000 [2], ABINPUT001[2]);
  buf(\oc8051_golden_model_1.ABINPUT000 [3], ABINPUT001[3]);
  buf(\oc8051_golden_model_1.ABINPUT000 [4], ABINPUT001[4]);
  buf(\oc8051_golden_model_1.ABINPUT000 [5], ABINPUT001[5]);
  buf(\oc8051_golden_model_1.ABINPUT000 [6], ABINPUT001[6]);
  buf(\oc8051_golden_model_1.ABINPUT000 [7], ABINPUT001[7]);
  buf(\oc8051_golden_model_1.n2453 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2453 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2453 [2], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2453 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2453 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2453 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2453 [6], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2453 [7], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2454 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2454 [1], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2454 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2454 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2454 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2454 [5], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2454 [6], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2876 [0], \oc8051_golden_model_1.PSW_d6 [0]);
  buf(\oc8051_golden_model_1.n2876 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2876 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2876 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2876 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2876 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2876 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2876 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1368 );
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1457 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.PSW_27 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.PSW_27 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.PSW_28 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.PSW_28 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.PSW_28 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.PSW_28 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.PSW_28 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.PSW_28 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.PSW_28 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.PSW_28 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.PSW_28 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.PSW_28 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.PSW_28 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.PSW_28 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.PSW_28 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.PSW_28 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.PSW_28 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.PSW_28 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.PSW_28 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.PSW_37 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.PSW_37 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.PSW_37 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.PSW_37 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.PSW_38 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.PSW_38 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.PSW_38 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.PSW_38 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.PSW_38 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.PSW_38 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.PSW_38 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.PSW_38 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.PSW_38 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.PSW_38 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.PSW_38 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.PSW_38 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.PSW_38 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.PSW_38 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.PSW_38 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.PSW_38 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.PSW_38 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.PSW_38 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.PSW_38 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.PSW_38 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.PSW_38 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.PSW_38 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.PSW_38 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.PSW_38 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.PSW_38 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.PSW_38 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.PSW_38 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.PSW_38 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.PSW_47 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.PSW_56 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n2086 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2103 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2229 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2470 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2500 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2529 );
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2514 [1]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2514 [5]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2514 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2529 );
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2514 [1]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2514 [5]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2514 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n1214 );
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2596 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.PSW_b6 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.PSW_b9 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.PSW_b9 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.PSW_b9 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.PSW_b9 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.PSW_b9 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.PSW_b9 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.PSW_b9 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2714 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2838 [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.PSW_d6 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2895 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2913 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.PSW_c5 [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.PSW_c5 [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.PSW_c5 [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.PSW_c5 [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.PSW_c5 [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.PSW_c5 [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.PSW_c5 [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fa [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_fa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fb [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_fb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fc [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_fc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fd [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_fd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fe [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_fe [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fe [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fe [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fe [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fe [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fe [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fe [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ff [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.PSW_ff [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ff [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ff [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ff [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ff [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ff [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ff [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0573 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n0573 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n0573 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n0573 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n0573 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n0573 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n0573 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n0573 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n0606 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n0606 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n0606 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n0606 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n0606 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n0606 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n0606 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n0606 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n0713 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0713 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0713 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0713 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0713 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0713 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0713 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0713 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0713 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0745 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0745 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0745 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0745 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0745 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0745 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0745 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0745 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0745 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0745 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0745 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0745 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0745 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0745 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0745 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0745 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1004 [8], \oc8051_golden_model_1.P2 [0]);
  buf(\oc8051_golden_model_1.n1004 [9], \oc8051_golden_model_1.P2 [1]);
  buf(\oc8051_golden_model_1.n1004 [10], \oc8051_golden_model_1.P2 [2]);
  buf(\oc8051_golden_model_1.n1004 [11], \oc8051_golden_model_1.P2 [3]);
  buf(\oc8051_golden_model_1.n1004 [12], \oc8051_golden_model_1.P2 [4]);
  buf(\oc8051_golden_model_1.n1004 [13], \oc8051_golden_model_1.P2 [5]);
  buf(\oc8051_golden_model_1.n1004 [14], \oc8051_golden_model_1.P2 [6]);
  buf(\oc8051_golden_model_1.n1004 [15], \oc8051_golden_model_1.P2 [7]);
  buf(\oc8051_golden_model_1.n1008 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1008 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1008 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1008 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1008 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1008 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1008 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1009 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1010 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1023 , \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n1024 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n1024 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1024 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1024 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1024 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1024 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1024 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1024 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1031 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1031 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1031 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1031 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1031 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1031 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1031 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1031 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1032 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1033 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1034 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1035 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1036 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1037 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1038 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1039 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1047 [0], \oc8051_golden_model_1.PSW_03 [0]);
  buf(\oc8051_golden_model_1.n1047 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1047 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1047 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1047 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1047 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1047 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1047 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1064 [0], \oc8051_golden_model_1.PSW_04 [0]);
  buf(\oc8051_golden_model_1.n1064 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1064 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1064 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1064 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1064 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1064 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1064 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2469 , \oc8051_golden_model_1.n2470 [0]);
  buf(\oc8051_golden_model_1.n2470 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2470 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2470 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2470 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2474 , \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2476 , \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2482 , \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2483 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2483 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2483 [2], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2483 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2483 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2483 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2483 [6], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2483 [7], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2484 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2484 [1], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2484 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2484 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2484 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2484 [5], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2484 [6], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n1157 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1157 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1157 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1157 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1159 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1161 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1161 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1162 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1162 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1163 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1163 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1164 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1164 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1165 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1165 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1166 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1166 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1167 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2499 , \oc8051_golden_model_1.n2500 [0]);
  buf(\oc8051_golden_model_1.n2500 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2500 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2500 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2500 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2504 , \oc8051_golden_model_1.n2514 [6]);
  buf(\oc8051_golden_model_1.n2506 , \oc8051_golden_model_1.n2514 [5]);
  buf(\oc8051_golden_model_1.n2512 , \oc8051_golden_model_1.n2514 [1]);
  buf(\oc8051_golden_model_1.n2513 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2513 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2513 [2], \oc8051_golden_model_1.n2514 [1]);
  buf(\oc8051_golden_model_1.n2513 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2513 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2513 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2513 [6], \oc8051_golden_model_1.n2514 [5]);
  buf(\oc8051_golden_model_1.n2513 [7], \oc8051_golden_model_1.n2514 [6]);
  buf(\oc8051_golden_model_1.n2514 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2514 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2514 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2514 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1259 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1260 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1261 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1261 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1261 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1261 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1261 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1261 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1261 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1262 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1262 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1262 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1262 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1262 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1262 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1262 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1262 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1265 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1266 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1266 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1267 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1267 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1267 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1267 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1267 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1267 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1268 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1268 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1268 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1268 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1268 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1268 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1268 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1269 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1270 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1271 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1272 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1273 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1274 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1276 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1284 [0], \oc8051_golden_model_1.PSW_13 [0]);
  buf(\oc8051_golden_model_1.n1284 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1284 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1284 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1284 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1284 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1284 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1284 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2530 [0], \oc8051_golden_model_1.n2529 );
  buf(\oc8051_golden_model_1.n2530 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2530 [2], \oc8051_golden_model_1.n2514 [1]);
  buf(\oc8051_golden_model_1.n2530 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2530 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2530 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2530 [6], \oc8051_golden_model_1.n2514 [5]);
  buf(\oc8051_golden_model_1.n2530 [7], \oc8051_golden_model_1.n2514 [6]);
  buf(\oc8051_golden_model_1.n2534 , \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2536 , \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n1301 [0], \oc8051_golden_model_1.PSW_14 [0]);
  buf(\oc8051_golden_model_1.n1301 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1301 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1301 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1301 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1301 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1301 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1301 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2542 , \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2543 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2543 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2543 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2543 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2543 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2543 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2543 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2543 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2544 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2544 [1], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2544 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2544 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2544 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2544 [5], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2544 [6], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2559 , \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.n2560 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2560 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2560 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2560 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2562 , \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2563 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2563 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2563 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2563 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2563 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2563 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2563 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2563 [7], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2564 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2564 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2564 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2564 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2564 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2564 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2564 [6], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2565 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n2565 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2565 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2565 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2565 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2565 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2565 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1343 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1343 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1343 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1343 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1343 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1343 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1343 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1343 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1345 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1345 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1345 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1345 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1345 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1345 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1345 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1345 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1346 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1347 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1348 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1351 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1352 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1353 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2566 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2566 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2566 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2566 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2566 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2566 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2566 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [7], \oc8051_golden_model_1.n1214 );
  buf(\oc8051_golden_model_1.n2567 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2567 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2567 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2567 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2567 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2567 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2567 [6], \oc8051_golden_model_1.n1214 );
  buf(\oc8051_golden_model_1.n2568 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n2568 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2568 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2568 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2568 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2568 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2568 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2568 [7], \oc8051_golden_model_1.n1214 );
  buf(\oc8051_golden_model_1.n1360 , \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.n1361 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1361 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1361 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1361 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1361 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1361 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1361 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2572 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2572 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2572 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2572 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2572 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2572 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2572 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2572 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2572 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [15], 1'b0);
  buf(\oc8051_golden_model_1.n1363 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1363 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1363 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1363 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1363 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1363 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1363 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1363 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1363 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1367 [8], \oc8051_golden_model_1.n1368 );
  buf(\oc8051_golden_model_1.n1369 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1369 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1369 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1369 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1370 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1370 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1370 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1374 [4], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1375 , \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1376 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1376 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1376 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1376 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1376 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1376 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1376 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1376 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1376 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2578 , \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2579 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2579 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2579 [2], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2579 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2579 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2579 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2579 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2579 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2580 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2580 [1], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2580 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2580 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2580 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2580 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2580 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1384 , \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1385 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1385 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1385 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1385 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1385 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1385 [7], \oc8051_golden_model_1.n1368 );
  buf(\oc8051_golden_model_1.n1386 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1386 [1], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1386 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1386 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1386 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1386 [5], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1386 [6], \oc8051_golden_model_1.n1368 );
  buf(\oc8051_golden_model_1.n2595 , \oc8051_golden_model_1.n2596 [0]);
  buf(\oc8051_golden_model_1.n2596 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2596 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2596 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2596 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2596 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2596 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1401 , \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.n1402 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1402 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1402 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1402 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1402 [7], \oc8051_golden_model_1.n1368 );
  buf(\oc8051_golden_model_1.n1424 [8], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1425 , \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n2599 , \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2600 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2600 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2600 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2600 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2600 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2600 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2600 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2600 [7], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n1430 [4], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1431 , \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n2601 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2601 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2601 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2601 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2601 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2601 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2601 [6], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2602 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n2602 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2602 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2602 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2602 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2602 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2602 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1439 , \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1440 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1440 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1440 [2], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1440 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1440 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1440 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1440 [6], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1440 [7], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1441 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1441 [1], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1441 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1441 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1441 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1441 [5], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1441 [6], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1456 , \oc8051_golden_model_1.n1457 [0]);
  buf(\oc8051_golden_model_1.n1457 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1457 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1457 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1457 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1459 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n1459 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n1459 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n1459 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n1459 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1459 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1459 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1459 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1459 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1463 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n1463 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n1463 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n1463 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n1464 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n1464 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n1464 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n1464 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n1464 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1466 [4], \oc8051_golden_model_1.PSW_27 [6]);
  buf(\oc8051_golden_model_1.n1467 , \oc8051_golden_model_1.PSW_27 [6]);
  buf(\oc8051_golden_model_1.n1468 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n1468 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n1468 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n1468 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n1468 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1468 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1468 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1468 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1468 [8], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1476 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1476 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1476 [2], \oc8051_golden_model_1.PSW_26 [2]);
  buf(\oc8051_golden_model_1.n1476 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1476 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1476 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1476 [6], \oc8051_golden_model_1.PSW_27 [6]);
  buf(\oc8051_golden_model_1.n1476 [7], \oc8051_golden_model_1.PSW_26 [7]);
  buf(\oc8051_golden_model_1.n1477 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1477 [1], \oc8051_golden_model_1.PSW_26 [2]);
  buf(\oc8051_golden_model_1.n1477 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1477 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1477 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1477 [5], \oc8051_golden_model_1.PSW_27 [6]);
  buf(\oc8051_golden_model_1.n1477 [6], \oc8051_golden_model_1.PSW_26 [7]);
  buf(\oc8051_golden_model_1.n2634 , \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2635 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2635 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2635 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2635 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2635 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2635 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2635 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2635 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2636 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2636 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2636 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2636 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2636 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2636 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2636 [6], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2637 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n2637 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2637 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2637 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2637 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2637 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2637 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2643 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2643 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2643 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2643 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2643 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2643 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2643 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2643 [7], \oc8051_golden_model_1.PSW_b4 [7]);
  buf(\oc8051_golden_model_1.n1492 , \oc8051_golden_model_1.PSW_27 [0]);
  buf(\oc8051_golden_model_1.n1493 [0], \oc8051_golden_model_1.PSW_27 [0]);
  buf(\oc8051_golden_model_1.n1493 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1493 [2], \oc8051_golden_model_1.PSW_26 [2]);
  buf(\oc8051_golden_model_1.n1493 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1493 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1493 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1493 [6], \oc8051_golden_model_1.PSW_27 [6]);
  buf(\oc8051_golden_model_1.n1493 [7], \oc8051_golden_model_1.PSW_26 [7]);
  buf(\oc8051_golden_model_1.n2644 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2644 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2644 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2644 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2644 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2644 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2644 [6], \oc8051_golden_model_1.PSW_b4 [7]);
  buf(\oc8051_golden_model_1.n2645 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n2645 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2645 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2645 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2645 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2645 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2645 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2645 [7], \oc8051_golden_model_1.PSW_b4 [7]);
  buf(\oc8051_golden_model_1.n2651 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2651 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2651 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2651 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2651 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2651 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2651 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2651 [7], \oc8051_golden_model_1.PSW_b5 [7]);
  buf(\oc8051_golden_model_1.n1505 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1505 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1505 [2], \oc8051_golden_model_1.PSW_27 [2]);
  buf(\oc8051_golden_model_1.n1505 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1505 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1505 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1505 [6], \oc8051_golden_model_1.PSW_27 [6]);
  buf(\oc8051_golden_model_1.n1505 [7], \oc8051_golden_model_1.PSW_27 [7]);
  buf(\oc8051_golden_model_1.n1506 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1506 [1], \oc8051_golden_model_1.PSW_27 [2]);
  buf(\oc8051_golden_model_1.n1506 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1506 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1506 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1506 [5], \oc8051_golden_model_1.PSW_27 [6]);
  buf(\oc8051_golden_model_1.n1506 [6], \oc8051_golden_model_1.PSW_27 [7]);
  buf(\oc8051_golden_model_1.n1507 [0], \oc8051_golden_model_1.PSW_27 [0]);
  buf(\oc8051_golden_model_1.n1507 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1507 [2], \oc8051_golden_model_1.PSW_27 [2]);
  buf(\oc8051_golden_model_1.n1507 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1507 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1507 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1507 [6], \oc8051_golden_model_1.PSW_27 [6]);
  buf(\oc8051_golden_model_1.n1507 [7], \oc8051_golden_model_1.PSW_27 [7]);
  buf(\oc8051_golden_model_1.n2652 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2652 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2652 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2652 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2652 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2652 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2652 [6], \oc8051_golden_model_1.PSW_b5 [7]);
  buf(\oc8051_golden_model_1.n1509 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1509 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1509 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1509 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1509 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1509 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1509 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1509 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1509 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2653 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n2653 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2653 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2653 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2653 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2653 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2653 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2653 [7], \oc8051_golden_model_1.PSW_b5 [7]);
  buf(\oc8051_golden_model_1.n1511 [8], \oc8051_golden_model_1.PSW_28 [7]);
  buf(\oc8051_golden_model_1.n1512 , \oc8051_golden_model_1.PSW_28 [7]);
  buf(\oc8051_golden_model_1.n1513 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1513 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1513 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1513 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1513 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1515 [4], \oc8051_golden_model_1.PSW_28 [6]);
  buf(\oc8051_golden_model_1.n1516 , \oc8051_golden_model_1.PSW_28 [6]);
  buf(\oc8051_golden_model_1.n1517 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1517 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1517 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1517 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1517 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1517 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1517 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1517 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1517 [8], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n2658 , \oc8051_golden_model_1.PSW_b6 [7]);
  buf(\oc8051_golden_model_1.n2659 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2659 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2659 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2659 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2659 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2659 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2659 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2659 [7], \oc8051_golden_model_1.PSW_b6 [7]);
  buf(\oc8051_golden_model_1.n2660 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2660 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2660 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2660 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2660 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2660 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2660 [6], \oc8051_golden_model_1.PSW_b6 [7]);
  buf(\oc8051_golden_model_1.n1524 , \oc8051_golden_model_1.PSW_28 [2]);
  buf(\oc8051_golden_model_1.n1525 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1525 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1525 [2], \oc8051_golden_model_1.PSW_28 [2]);
  buf(\oc8051_golden_model_1.n1525 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1525 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1525 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1525 [6], \oc8051_golden_model_1.PSW_28 [6]);
  buf(\oc8051_golden_model_1.n1525 [7], \oc8051_golden_model_1.PSW_28 [7]);
  buf(\oc8051_golden_model_1.n1526 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1526 [1], \oc8051_golden_model_1.PSW_28 [2]);
  buf(\oc8051_golden_model_1.n1526 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1526 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1526 [5], \oc8051_golden_model_1.PSW_28 [6]);
  buf(\oc8051_golden_model_1.n1526 [6], \oc8051_golden_model_1.PSW_28 [7]);
  buf(\oc8051_golden_model_1.n2661 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n2661 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2661 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2661 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2661 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2661 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2661 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2661 [7], \oc8051_golden_model_1.PSW_b6 [7]);
  buf(\oc8051_golden_model_1.n2666 , \oc8051_golden_model_1.PSW_b9 [7]);
  buf(\oc8051_golden_model_1.n2667 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2667 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2667 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2667 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2667 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2667 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2667 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2667 [7], \oc8051_golden_model_1.PSW_b9 [7]);
  buf(\oc8051_golden_model_1.n2668 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2668 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2668 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2668 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2668 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2668 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2668 [6], \oc8051_golden_model_1.PSW_b9 [7]);
  buf(\oc8051_golden_model_1.n2669 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n2669 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2669 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2669 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2669 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2669 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2669 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2669 [7], \oc8051_golden_model_1.PSW_b9 [7]);
  buf(\oc8051_golden_model_1.n1541 , \oc8051_golden_model_1.PSW_28 [0]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.PSW_28 [0]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.PSW_28 [2]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.PSW_28 [6]);
  buf(\oc8051_golden_model_1.n1542 [7], \oc8051_golden_model_1.PSW_28 [7]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1545 , \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [2], \oc8051_golden_model_1.PSW_28 [2]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1546 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1546 [7], \oc8051_golden_model_1.PSW_28 [7]);
  buf(\oc8051_golden_model_1.n1547 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1547 [1], \oc8051_golden_model_1.PSW_28 [2]);
  buf(\oc8051_golden_model_1.n1547 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1547 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1547 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1547 [5], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1547 [6], \oc8051_golden_model_1.PSW_28 [7]);
  buf(\oc8051_golden_model_1.n1548 [0], \oc8051_golden_model_1.PSW_28 [0]);
  buf(\oc8051_golden_model_1.n1548 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1548 [2], \oc8051_golden_model_1.PSW_28 [2]);
  buf(\oc8051_golden_model_1.n1548 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1548 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1548 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1548 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1548 [7], \oc8051_golden_model_1.PSW_28 [7]);
  buf(\oc8051_golden_model_1.n1550 [8], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1551 , \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n2894 , \oc8051_golden_model_1.n2895 [0]);
  buf(\oc8051_golden_model_1.n2895 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2895 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2895 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2895 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2895 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2895 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2895 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2896 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2896 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2896 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2896 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2896 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2896 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2896 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1559 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1559 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1559 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1559 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1559 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1559 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1559 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1559 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1560 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1560 [1], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1560 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1560 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1560 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1560 [5], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1560 [6], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1561 [0], \oc8051_golden_model_1.PSW_28 [0]);
  buf(\oc8051_golden_model_1.n1561 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1561 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1561 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1561 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1561 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1561 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1562 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1562 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1562 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1562 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1562 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1562 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1562 [6], \oc8051_golden_model_1.PSW_28 [6]);
  buf(\oc8051_golden_model_1.n1562 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1563 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1563 [1], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1563 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1563 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1563 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1563 [5], \oc8051_golden_model_1.PSW_28 [6]);
  buf(\oc8051_golden_model_1.n1563 [6], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1564 [0], \oc8051_golden_model_1.PSW_28 [0]);
  buf(\oc8051_golden_model_1.n1564 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1564 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1564 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1564 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1564 [6], \oc8051_golden_model_1.PSW_28 [6]);
  buf(\oc8051_golden_model_1.n1567 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1567 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1567 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1567 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1567 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1567 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1567 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1567 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1567 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1568 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1568 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1568 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1568 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1568 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1568 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1568 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1569 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1569 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1569 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1569 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1569 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1569 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1569 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1569 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1570 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1570 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1570 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1570 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1570 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1570 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1570 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1570 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1571 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1571 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1571 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1571 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1571 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1571 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1571 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1572 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1573 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1574 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1575 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1576 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1577 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1578 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1579 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1587 [0], \oc8051_golden_model_1.PSW_33 [0]);
  buf(\oc8051_golden_model_1.n1587 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1587 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1587 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1587 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1587 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1587 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1587 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1588 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1588 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1591 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1595 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [4], 1'b0);
  buf(\oc8051_golden_model_1.n2694 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2694 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2694 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2694 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2694 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2694 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2694 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2695 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2695 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2695 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2695 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2695 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2695 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2695 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2696 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n2696 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2696 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2696 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2696 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2696 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2696 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2696 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2697 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2697 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2697 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2697 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2698 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2698 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2698 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2698 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2698 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2698 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2698 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2698 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1606 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1606 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1606 [2], \oc8051_golden_model_1.PSW_34 [2]);
  buf(\oc8051_golden_model_1.n1606 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1606 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1606 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1606 [6], \oc8051_golden_model_1.PSW_34 [6]);
  buf(\oc8051_golden_model_1.n1606 [7], \oc8051_golden_model_1.PSW_34 [7]);
  buf(\oc8051_golden_model_1.n1607 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1607 [1], \oc8051_golden_model_1.PSW_34 [2]);
  buf(\oc8051_golden_model_1.n1607 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1607 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1607 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1607 [5], \oc8051_golden_model_1.PSW_34 [6]);
  buf(\oc8051_golden_model_1.n1607 [6], \oc8051_golden_model_1.PSW_34 [7]);
  buf(\oc8051_golden_model_1.n2699 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2700 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2701 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2702 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2703 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2704 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2705 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2706 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2912 , \oc8051_golden_model_1.n2913 [0]);
  buf(\oc8051_golden_model_1.n2913 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2913 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2913 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2913 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2913 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2913 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2913 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1623 [0], \oc8051_golden_model_1.PSW_34 [0]);
  buf(\oc8051_golden_model_1.n1623 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1623 [2], \oc8051_golden_model_1.PSW_34 [2]);
  buf(\oc8051_golden_model_1.n1623 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1623 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1623 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1623 [6], \oc8051_golden_model_1.PSW_34 [6]);
  buf(\oc8051_golden_model_1.n1623 [7], \oc8051_golden_model_1.PSW_34 [7]);
  buf(\oc8051_golden_model_1.n2713 , \oc8051_golden_model_1.n2714 [0]);
  buf(\oc8051_golden_model_1.n2714 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2714 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2714 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2714 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2714 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2714 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2714 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1639 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1639 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1639 [2], \oc8051_golden_model_1.PSW_35 [2]);
  buf(\oc8051_golden_model_1.n1639 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1639 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1639 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1639 [6], \oc8051_golden_model_1.PSW_35 [6]);
  buf(\oc8051_golden_model_1.n1639 [7], \oc8051_golden_model_1.PSW_35 [7]);
  buf(\oc8051_golden_model_1.n1640 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1640 [1], \oc8051_golden_model_1.PSW_35 [2]);
  buf(\oc8051_golden_model_1.n1640 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1640 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1640 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1640 [5], \oc8051_golden_model_1.PSW_35 [6]);
  buf(\oc8051_golden_model_1.n1640 [6], \oc8051_golden_model_1.PSW_35 [7]);
  buf(\oc8051_golden_model_1.n1656 [0], \oc8051_golden_model_1.PSW_35 [0]);
  buf(\oc8051_golden_model_1.n1656 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1656 [2], \oc8051_golden_model_1.PSW_35 [2]);
  buf(\oc8051_golden_model_1.n1656 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1656 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1656 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1656 [6], \oc8051_golden_model_1.PSW_35 [6]);
  buf(\oc8051_golden_model_1.n1656 [7], \oc8051_golden_model_1.PSW_35 [7]);
  buf(\oc8051_golden_model_1.n1660 [8], \oc8051_golden_model_1.PSW_37 [7]);
  buf(\oc8051_golden_model_1.n1661 , \oc8051_golden_model_1.PSW_37 [7]);
  buf(\oc8051_golden_model_1.n1663 [4], \oc8051_golden_model_1.PSW_37 [6]);
  buf(\oc8051_golden_model_1.n1664 , \oc8051_golden_model_1.PSW_37 [6]);
  buf(\oc8051_golden_model_1.n1671 , \oc8051_golden_model_1.PSW_37 [2]);
  buf(\oc8051_golden_model_1.n1672 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1672 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1672 [2], \oc8051_golden_model_1.PSW_37 [2]);
  buf(\oc8051_golden_model_1.n1672 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1672 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1672 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1672 [6], \oc8051_golden_model_1.PSW_37 [6]);
  buf(\oc8051_golden_model_1.n1672 [7], \oc8051_golden_model_1.PSW_37 [7]);
  buf(\oc8051_golden_model_1.n1673 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1673 [1], \oc8051_golden_model_1.PSW_37 [2]);
  buf(\oc8051_golden_model_1.n1673 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1673 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1673 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1673 [5], \oc8051_golden_model_1.PSW_37 [6]);
  buf(\oc8051_golden_model_1.n1673 [6], \oc8051_golden_model_1.PSW_37 [7]);
  buf(\oc8051_golden_model_1.n1688 , \oc8051_golden_model_1.PSW_37 [0]);
  buf(\oc8051_golden_model_1.n1689 [0], \oc8051_golden_model_1.PSW_37 [0]);
  buf(\oc8051_golden_model_1.n1689 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1689 [2], \oc8051_golden_model_1.PSW_37 [2]);
  buf(\oc8051_golden_model_1.n1689 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1689 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1689 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1689 [6], \oc8051_golden_model_1.PSW_37 [6]);
  buf(\oc8051_golden_model_1.n1689 [7], \oc8051_golden_model_1.PSW_37 [7]);
  buf(\oc8051_golden_model_1.n1693 [8], \oc8051_golden_model_1.PSW_38 [7]);
  buf(\oc8051_golden_model_1.n1694 , \oc8051_golden_model_1.PSW_38 [7]);
  buf(\oc8051_golden_model_1.n1696 [4], \oc8051_golden_model_1.PSW_38 [6]);
  buf(\oc8051_golden_model_1.n1697 , \oc8051_golden_model_1.PSW_38 [6]);
  buf(\oc8051_golden_model_1.n1704 , \oc8051_golden_model_1.PSW_38 [2]);
  buf(\oc8051_golden_model_1.n1705 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1705 [2], \oc8051_golden_model_1.PSW_38 [2]);
  buf(\oc8051_golden_model_1.n1705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1705 [6], \oc8051_golden_model_1.PSW_38 [6]);
  buf(\oc8051_golden_model_1.n1705 [7], \oc8051_golden_model_1.PSW_38 [7]);
  buf(\oc8051_golden_model_1.n1706 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1706 [1], \oc8051_golden_model_1.PSW_38 [2]);
  buf(\oc8051_golden_model_1.n1706 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1706 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1706 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1706 [5], \oc8051_golden_model_1.PSW_38 [6]);
  buf(\oc8051_golden_model_1.n1706 [6], \oc8051_golden_model_1.PSW_38 [7]);
  buf(\oc8051_golden_model_1.n1721 , \oc8051_golden_model_1.PSW_38 [0]);
  buf(\oc8051_golden_model_1.n1722 [0], \oc8051_golden_model_1.PSW_38 [0]);
  buf(\oc8051_golden_model_1.n1722 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1722 [2], \oc8051_golden_model_1.PSW_38 [2]);
  buf(\oc8051_golden_model_1.n1722 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1722 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1722 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1722 [6], \oc8051_golden_model_1.PSW_38 [6]);
  buf(\oc8051_golden_model_1.n1722 [7], \oc8051_golden_model_1.PSW_38 [7]);
  buf(\oc8051_golden_model_1.n1749 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n1749 [1], \oc8051_golden_model_1.PSW_42 [1]);
  buf(\oc8051_golden_model_1.n1749 [2], \oc8051_golden_model_1.PSW_42 [2]);
  buf(\oc8051_golden_model_1.n1749 [3], \oc8051_golden_model_1.PSW_42 [3]);
  buf(\oc8051_golden_model_1.n1749 [4], \oc8051_golden_model_1.PSW_42 [4]);
  buf(\oc8051_golden_model_1.n1749 [5], \oc8051_golden_model_1.PSW_42 [5]);
  buf(\oc8051_golden_model_1.n1749 [6], \oc8051_golden_model_1.PSW_42 [6]);
  buf(\oc8051_golden_model_1.n1749 [7], \oc8051_golden_model_1.PSW_42 [7]);
  buf(\oc8051_golden_model_1.n1805 [0], \oc8051_golden_model_1.PSW_44 [0]);
  buf(\oc8051_golden_model_1.n1805 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1805 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1805 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1805 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1805 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1805 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1805 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1822 [0], \oc8051_golden_model_1.PSW_45 [0]);
  buf(\oc8051_golden_model_1.n1822 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1822 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1822 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1822 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1822 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1822 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1822 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1838 , \oc8051_golden_model_1.PSW_47 [0]);
  buf(\oc8051_golden_model_1.n1839 [0], \oc8051_golden_model_1.PSW_47 [0]);
  buf(\oc8051_golden_model_1.n1839 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1839 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1839 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1839 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1839 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1839 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1839 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1855 , \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.n1856 [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.n1856 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1856 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1856 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1856 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1856 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1856 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1856 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1881 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n1881 [1], \oc8051_golden_model_1.PSW_52 [1]);
  buf(\oc8051_golden_model_1.n1881 [2], \oc8051_golden_model_1.PSW_52 [2]);
  buf(\oc8051_golden_model_1.n1881 [3], \oc8051_golden_model_1.PSW_52 [3]);
  buf(\oc8051_golden_model_1.n1881 [4], \oc8051_golden_model_1.PSW_52 [4]);
  buf(\oc8051_golden_model_1.n1881 [5], \oc8051_golden_model_1.PSW_52 [5]);
  buf(\oc8051_golden_model_1.n1881 [6], \oc8051_golden_model_1.PSW_52 [6]);
  buf(\oc8051_golden_model_1.n1881 [7], \oc8051_golden_model_1.PSW_52 [7]);
  buf(\oc8051_golden_model_1.n2766 , \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.n2767 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2767 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2767 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2767 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2767 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2767 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2767 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2782 , \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.n2783 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2783 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2783 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2783 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2783 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2783 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2783 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1937 [0], \oc8051_golden_model_1.PSW_54 [0]);
  buf(\oc8051_golden_model_1.n1937 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1937 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1937 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1937 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1937 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1937 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1937 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1954 [0], \oc8051_golden_model_1.PSW_55 [0]);
  buf(\oc8051_golden_model_1.n1954 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1954 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1954 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1954 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1954 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1954 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1954 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1970 , \oc8051_golden_model_1.PSW_56 [0]);
  buf(\oc8051_golden_model_1.n1971 [0], \oc8051_golden_model_1.PSW_56 [0]);
  buf(\oc8051_golden_model_1.n1971 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1971 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1971 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1971 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1971 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1971 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1971 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2815 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2815 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2815 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2815 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2815 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2815 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2815 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2815 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2816 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2816 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2816 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2816 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2816 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2816 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2816 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2817 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n2817 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2817 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2817 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2817 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2817 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2817 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2817 [7], 1'b1);
  buf(\oc8051_golden_model_1.n1987 , \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.n1988 [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.n1988 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1988 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1988 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1988 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1988 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1988 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1988 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2836 , \oc8051_golden_model_1.n2838 [6]);
  buf(\oc8051_golden_model_1.n2837 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2837 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2837 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2837 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2837 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2837 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2837 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2837 [7], \oc8051_golden_model_1.n2838 [6]);
  buf(\oc8051_golden_model_1.n2838 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2838 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2838 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2838 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2838 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2838 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2085 , \oc8051_golden_model_1.n2086 [0]);
  buf(\oc8051_golden_model_1.n2086 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2086 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2086 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2086 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2086 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2086 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2086 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2102 , \oc8051_golden_model_1.n2103 [0]);
  buf(\oc8051_golden_model_1.n2103 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2103 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2103 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2103 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2103 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2103 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2103 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2119 , \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.n2120 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2120 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2120 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2120 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2120 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2120 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2120 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2136 , \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.n2137 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2137 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2137 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2137 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2137 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2137 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2137 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2141 , \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2142 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2142 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2142 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2142 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2142 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2142 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2142 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2143 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2143 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2143 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2143 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2143 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2143 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2143 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2143 [7], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2144 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2144 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2144 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2144 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2144 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2144 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2144 [6], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2145 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n2145 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2145 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2145 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2145 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2145 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2145 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2160 , \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.n2161 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2161 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2161 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2161 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2161 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2161 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2201 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2201 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2201 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2201 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2201 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2201 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2201 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2201 [7], \oc8051_golden_model_1.PSW_82 [7]);
  buf(\oc8051_golden_model_1.n2202 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2202 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2202 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2202 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2202 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2202 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2202 [6], \oc8051_golden_model_1.PSW_82 [7]);
  buf(\oc8051_golden_model_1.n2203 [0], \oc8051_golden_model_1.PSW_30 [0]);
  buf(\oc8051_golden_model_1.n2203 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2203 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2203 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2203 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2203 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2203 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2203 [7], \oc8051_golden_model_1.PSW_82 [7]);
  buf(\oc8051_golden_model_1.n2210 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2210 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2210 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2210 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2211 , \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2212 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2212 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2212 [2], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2212 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2212 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2212 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2212 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2212 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2213 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2213 [1], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2213 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2213 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2213 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2213 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2213 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2228 , \oc8051_golden_model_1.n2229 [0]);
  buf(\oc8051_golden_model_1.n2229 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2229 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2229 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2229 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2229 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2229 [7], 1'b0);
  buf(\oc8051_top_1.sub_result [0], ABINPUT[27]);
  buf(\oc8051_top_1.sub_result [1], ABINPUT[28]);
  buf(\oc8051_top_1.sub_result [2], ABINPUT[29]);
  buf(\oc8051_top_1.sub_result [3], ABINPUT[30]);
  buf(\oc8051_top_1.sub_result [4], ABINPUT[31]);
  buf(\oc8051_top_1.sub_result [5], ABINPUT[32]);
  buf(\oc8051_top_1.sub_result [6], ABINPUT[33]);
  buf(\oc8051_top_1.sub_result [7], ABINPUT[34]);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.ABINPUT [9], ABINPUT[9]);
  buf(\oc8051_top_1.ABINPUT [10], ABINPUT[10]);
  buf(\oc8051_top_1.ABINPUT [11], ABINPUT[11]);
  buf(\oc8051_top_1.ABINPUT [12], ABINPUT[12]);
  buf(\oc8051_top_1.ABINPUT [13], ABINPUT[13]);
  buf(\oc8051_top_1.ABINPUT [14], ABINPUT[14]);
  buf(\oc8051_top_1.ABINPUT [15], ABINPUT[15]);
  buf(\oc8051_top_1.ABINPUT [16], ABINPUT[16]);
  buf(\oc8051_top_1.ABINPUT [17], ABINPUT[17]);
  buf(\oc8051_top_1.ABINPUT [18], ABINPUT[18]);
  buf(\oc8051_top_1.ABINPUT [19], ABINPUT[19]);
  buf(\oc8051_top_1.ABINPUT [20], ABINPUT[20]);
  buf(\oc8051_top_1.ABINPUT [21], ABINPUT[21]);
  buf(\oc8051_top_1.ABINPUT [22], ABINPUT[22]);
  buf(\oc8051_top_1.ABINPUT [23], ABINPUT[23]);
  buf(\oc8051_top_1.ABINPUT [24], ABINPUT[24]);
  buf(\oc8051_top_1.ABINPUT [25], ABINPUT[25]);
  buf(\oc8051_top_1.ABINPUT [26], ABINPUT[26]);
  buf(\oc8051_top_1.ABINPUT [27], ABINPUT[27]);
  buf(\oc8051_top_1.ABINPUT [28], ABINPUT[28]);
  buf(\oc8051_top_1.ABINPUT [29], ABINPUT[29]);
  buf(\oc8051_top_1.ABINPUT [30], ABINPUT[30]);
  buf(\oc8051_top_1.ABINPUT [31], ABINPUT[31]);
  buf(\oc8051_top_1.ABINPUT [32], ABINPUT[32]);
  buf(\oc8051_top_1.ABINPUT [33], ABINPUT[33]);
  buf(\oc8051_top_1.ABINPUT [34], ABINPUT[34]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.desOv , ABINPUT[2]);
  buf(\oc8051_top_1.desAc , ABINPUT[1]);
  buf(\oc8051_top_1.desCy , ABINPUT[0]);
  buf(\oc8051_top_1.des2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.des2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.des2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.des2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.des2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.des2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.des2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.des2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.des1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.des1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.des1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.des1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.des1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.des1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.des1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.des1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.wr_dat [0], ABINPUT[3]);
  buf(\oc8051_top_1.wr_dat [1], ABINPUT[4]);
  buf(\oc8051_top_1.wr_dat [2], ABINPUT[5]);
  buf(\oc8051_top_1.wr_dat [3], ABINPUT[6]);
  buf(\oc8051_top_1.wr_dat [4], ABINPUT[7]);
  buf(\oc8051_top_1.wr_dat [5], ABINPUT[8]);
  buf(\oc8051_top_1.wr_dat [6], ABINPUT[9]);
  buf(\oc8051_top_1.wr_dat [7], ABINPUT[10]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(p12_equal, p1_valid_r);
  buf(IRAM_gm[0], ABINPUT009[0]);
  buf(IRAM_gm[1], ABINPUT009[1]);
  buf(IRAM_gm[2], ABINPUT009[2]);
  buf(IRAM_gm[3], ABINPUT009[3]);
  buf(IRAM_gm[4], ABINPUT009[4]);
  buf(IRAM_gm[5], ABINPUT009[5]);
  buf(IRAM_gm[6], ABINPUT009[6]);
  buf(IRAM_gm[7], ABINPUT009[7]);
  buf(IRAM_gm[8], ABINPUT009[8]);
  buf(IRAM_gm[9], ABINPUT009[9]);
  buf(IRAM_gm[10], ABINPUT009[10]);
  buf(IRAM_gm[11], ABINPUT009[11]);
  buf(IRAM_gm[12], ABINPUT009[12]);
  buf(IRAM_gm[13], ABINPUT009[13]);
  buf(IRAM_gm[14], ABINPUT009[14]);
  buf(IRAM_gm[15], ABINPUT009[15]);
  buf(IRAM_gm[16], ABINPUT009[16]);
  buf(IRAM_gm[17], ABINPUT009[17]);
  buf(IRAM_gm[18], ABINPUT009[18]);
  buf(IRAM_gm[19], ABINPUT009[19]);
  buf(IRAM_gm[20], ABINPUT009[20]);
  buf(IRAM_gm[21], ABINPUT009[21]);
  buf(IRAM_gm[22], ABINPUT009[22]);
  buf(IRAM_gm[23], ABINPUT009[23]);
  buf(IRAM_gm[24], ABINPUT009[24]);
  buf(IRAM_gm[25], ABINPUT009[25]);
  buf(IRAM_gm[26], ABINPUT009[26]);
  buf(IRAM_gm[27], ABINPUT009[27]);
  buf(IRAM_gm[28], ABINPUT009[28]);
  buf(IRAM_gm[29], ABINPUT009[29]);
  buf(IRAM_gm[30], ABINPUT009[30]);
  buf(IRAM_gm[31], ABINPUT009[31]);
  buf(IRAM_gm[32], ABINPUT009[32]);
  buf(IRAM_gm[33], ABINPUT009[33]);
  buf(IRAM_gm[34], ABINPUT009[34]);
  buf(IRAM_gm[35], ABINPUT009[35]);
  buf(IRAM_gm[36], ABINPUT009[36]);
  buf(IRAM_gm[37], ABINPUT009[37]);
  buf(IRAM_gm[38], ABINPUT009[38]);
  buf(IRAM_gm[39], ABINPUT009[39]);
  buf(IRAM_gm[40], ABINPUT009[40]);
  buf(IRAM_gm[41], ABINPUT009[41]);
  buf(IRAM_gm[42], ABINPUT009[42]);
  buf(IRAM_gm[43], ABINPUT009[43]);
  buf(IRAM_gm[44], ABINPUT009[44]);
  buf(IRAM_gm[45], ABINPUT009[45]);
  buf(IRAM_gm[46], ABINPUT009[46]);
  buf(IRAM_gm[47], ABINPUT009[47]);
  buf(IRAM_gm[48], ABINPUT009[48]);
  buf(IRAM_gm[49], ABINPUT009[49]);
  buf(IRAM_gm[50], ABINPUT009[50]);
  buf(IRAM_gm[51], ABINPUT009[51]);
  buf(IRAM_gm[52], ABINPUT009[52]);
  buf(IRAM_gm[53], ABINPUT009[53]);
  buf(IRAM_gm[54], ABINPUT009[54]);
  buf(IRAM_gm[55], ABINPUT009[55]);
  buf(IRAM_gm[56], ABINPUT009[56]);
  buf(IRAM_gm[57], ABINPUT009[57]);
  buf(IRAM_gm[58], ABINPUT009[58]);
  buf(IRAM_gm[59], ABINPUT009[59]);
  buf(IRAM_gm[60], ABINPUT009[60]);
  buf(IRAM_gm[61], ABINPUT009[61]);
  buf(IRAM_gm[62], ABINPUT009[62]);
  buf(IRAM_gm[63], ABINPUT009[63]);
  buf(IRAM_gm[64], ABINPUT009[64]);
  buf(IRAM_gm[65], ABINPUT009[65]);
  buf(IRAM_gm[66], ABINPUT009[66]);
  buf(IRAM_gm[67], ABINPUT009[67]);
  buf(IRAM_gm[68], ABINPUT009[68]);
  buf(IRAM_gm[69], ABINPUT009[69]);
  buf(IRAM_gm[70], ABINPUT009[70]);
  buf(IRAM_gm[71], ABINPUT009[71]);
  buf(IRAM_gm[72], ABINPUT009[72]);
  buf(IRAM_gm[73], ABINPUT009[73]);
  buf(IRAM_gm[74], ABINPUT009[74]);
  buf(IRAM_gm[75], ABINPUT009[75]);
  buf(IRAM_gm[76], ABINPUT009[76]);
  buf(IRAM_gm[77], ABINPUT009[77]);
  buf(IRAM_gm[78], ABINPUT009[78]);
  buf(IRAM_gm[79], ABINPUT009[79]);
  buf(IRAM_gm[80], ABINPUT009[80]);
  buf(IRAM_gm[81], ABINPUT009[81]);
  buf(IRAM_gm[82], ABINPUT009[82]);
  buf(IRAM_gm[83], ABINPUT009[83]);
  buf(IRAM_gm[84], ABINPUT009[84]);
  buf(IRAM_gm[85], ABINPUT009[85]);
  buf(IRAM_gm[86], ABINPUT009[86]);
  buf(IRAM_gm[87], ABINPUT009[87]);
  buf(IRAM_gm[88], ABINPUT009[88]);
  buf(IRAM_gm[89], ABINPUT009[89]);
  buf(IRAM_gm[90], ABINPUT009[90]);
  buf(IRAM_gm[91], ABINPUT009[91]);
  buf(IRAM_gm[92], ABINPUT009[92]);
  buf(IRAM_gm[93], ABINPUT009[93]);
  buf(IRAM_gm[94], ABINPUT009[94]);
  buf(IRAM_gm[95], ABINPUT009[95]);
  buf(IRAM_gm[96], ABINPUT009[96]);
  buf(IRAM_gm[97], ABINPUT009[97]);
  buf(IRAM_gm[98], ABINPUT009[98]);
  buf(IRAM_gm[99], ABINPUT009[99]);
  buf(IRAM_gm[100], ABINPUT009[100]);
  buf(IRAM_gm[101], ABINPUT009[101]);
  buf(IRAM_gm[102], ABINPUT009[102]);
  buf(IRAM_gm[103], ABINPUT009[103]);
  buf(IRAM_gm[104], ABINPUT009[104]);
  buf(IRAM_gm[105], ABINPUT009[105]);
  buf(IRAM_gm[106], ABINPUT009[106]);
  buf(IRAM_gm[107], ABINPUT009[107]);
  buf(IRAM_gm[108], ABINPUT009[108]);
  buf(IRAM_gm[109], ABINPUT009[109]);
  buf(IRAM_gm[110], ABINPUT009[110]);
  buf(IRAM_gm[111], ABINPUT009[111]);
  buf(IRAM_gm[112], ABINPUT009[112]);
  buf(IRAM_gm[113], ABINPUT009[113]);
  buf(IRAM_gm[114], ABINPUT009[114]);
  buf(IRAM_gm[115], ABINPUT009[115]);
  buf(IRAM_gm[116], ABINPUT009[116]);
  buf(IRAM_gm[117], ABINPUT009[117]);
  buf(IRAM_gm[118], ABINPUT009[118]);
  buf(IRAM_gm[119], ABINPUT009[119]);
  buf(IRAM_gm[120], ABINPUT009[120]);
  buf(IRAM_gm[121], ABINPUT009[121]);
  buf(IRAM_gm[122], ABINPUT009[122]);
  buf(IRAM_gm[123], ABINPUT009[123]);
  buf(IRAM_gm[124], ABINPUT009[124]);
  buf(IRAM_gm[125], ABINPUT009[125]);
  buf(IRAM_gm[126], ABINPUT009[126]);
  buf(IRAM_gm[127], ABINPUT009[127]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm_next[0], ABINPUT008[0]);
  buf(PSW_gm_next[1], ABINPUT008[1]);
  buf(PSW_gm_next[2], ABINPUT008[2]);
  buf(PSW_gm_next[3], ABINPUT008[3]);
  buf(PSW_gm_next[4], ABINPUT008[4]);
  buf(PSW_gm_next[5], ABINPUT008[5]);
  buf(PSW_gm_next[6], ABINPUT008[6]);
  buf(PSW_gm_next[7], ABINPUT008[7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
