
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire [15:0] _26842_;
  wire [7:0] _26843_;
  wire [7:0] _26844_;
  wire [7:0] _26845_;
  wire [7:0] _26846_;
  wire [7:0] _26847_;
  wire [7:0] _26848_;
  wire [7:0] _26849_;
  wire [7:0] _26850_;
  wire [7:0] _26851_;
  wire [7:0] _26852_;
  wire [7:0] _26853_;
  wire [7:0] _26854_;
  wire [7:0] _26855_;
  wire [7:0] _26856_;
  wire [7:0] _26857_;
  wire [7:0] _26858_;
  wire _26859_;
  wire [7:0] _26860_;
  wire [2:0] _26861_;
  wire [2:0] _26862_;
  wire [1:0] _26863_;
  wire [7:0] _26864_;
  wire _26865_;
  wire [1:0] _26866_;
  wire [1:0] _26867_;
  wire [2:0] _26868_;
  wire [2:0] _26869_;
  wire [1:0] _26870_;
  wire [3:0] _26871_;
  wire [1:0] _26872_;
  wire _26873_;
  wire [7:0] _26874_;
  wire [7:0] _26875_;
  wire [7:0] _26876_;
  wire [7:0] _26877_;
  wire [7:0] _26878_;
  wire [7:0] _26879_;
  wire [7:0] _26880_;
  wire [7:0] _26881_;
  wire [15:0] _26882_;
  wire [15:0] _26883_;
  wire _26884_;
  wire [4:0] _26885_;
  wire [7:0] _26886_;
  wire [7:0] _26887_;
  wire _26888_;
  wire _26889_;
  wire [15:0] _26890_;
  wire [15:0] _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire [7:0] _26895_;
  wire [2:0] _26896_;
  wire [7:0] _26897_;
  wire _26898_;
  wire [7:0] _26899_;
  wire _26900_;
  wire _26901_;
  wire [3:0] _26902_;
  wire [31:0] _26903_;
  wire [31:0] _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire [15:0] _26908_;
  wire _26909_;
  wire _26910_;
  wire [7:0] _26911_;
  wire _26912_;
  wire [2:0] _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire [3:0] _27304_;
  wire _27305_;
  wire _27306_;
  wire [7:0] _27307_;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not _27308_ (_22762_, rst);
  not _27309_ (_22763_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  nor _27310_ (_22764_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _27311_ (_22765_, _22764_, _22763_);
  not _27312_ (_22766_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _27313_ (_22767_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  and _27314_ (_22768_, _22767_, _22766_);
  and _27315_ (_22769_, _22768_, _22765_);
  and _27316_ (_22770_, _22769_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and _27317_ (_22771_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _27318_ (_22772_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _27319_ (_22773_, _22770_, _22772_);
  or _27320_ (_22775_, _22773_, _22771_);
  and _27321_ (_26882_[0], _22775_, _22762_);
  and _27322_ (_22777_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _27323_ (_22778_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _27324_ (_22780_, _22770_, _22778_);
  or _27325_ (_22781_, _22780_, _22777_);
  and _27326_ (_26882_[1], _22781_, _22762_);
  and _27327_ (_22782_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _27328_ (_22783_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _27329_ (_22784_, _22770_, _22783_);
  or _27330_ (_22785_, _22784_, _22782_);
  and _27331_ (_26882_[2], _22785_, _22762_);
  and _27332_ (_22786_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _27333_ (_22788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _27334_ (_22789_, _22770_, _22788_);
  or _27335_ (_22791_, _22789_, _22786_);
  and _27336_ (_26882_[3], _22791_, _22762_);
  and _27337_ (_22793_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not _27338_ (_22794_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _27339_ (_22795_, _22770_, _22794_);
  or _27340_ (_22796_, _22795_, _22793_);
  and _27341_ (_26882_[4], _22796_, _22762_);
  and _27342_ (_22797_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not _27343_ (_22798_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _27344_ (_22799_, _22770_, _22798_);
  or _27345_ (_22800_, _22799_, _22797_);
  and _27346_ (_26882_[5], _22800_, _22762_);
  and _27347_ (_22801_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not _27348_ (_22802_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _27349_ (_22803_, _22770_, _22802_);
  or _27350_ (_22804_, _22803_, _22801_);
  and _27351_ (_26882_[6], _22804_, _22762_);
  and _27352_ (_22805_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _27353_ (_22806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _27354_ (_22807_, _22770_, _22806_);
  or _27355_ (_22808_, _22807_, _22805_);
  and _27356_ (_26882_[7], _22808_, _22762_);
  and _27357_ (_22809_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not _27358_ (_22810_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _27359_ (_22811_, _22770_, _22810_);
  or _27360_ (_22812_, _22811_, _22809_);
  and _27361_ (_26882_[8], _22812_, _22762_);
  and _27362_ (_22813_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not _27363_ (_22814_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _27364_ (_22815_, _22770_, _22814_);
  or _27365_ (_22816_, _22815_, _22813_);
  and _27366_ (_26882_[9], _22816_, _22762_);
  and _27367_ (_22817_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not _27368_ (_22819_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _27369_ (_22820_, _22770_, _22819_);
  or _27370_ (_22821_, _22820_, _22817_);
  and _27371_ (_26882_[10], _22821_, _22762_);
  and _27372_ (_22822_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not _27373_ (_22823_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _27374_ (_22824_, _22770_, _22823_);
  or _27375_ (_22825_, _22824_, _22822_);
  and _27376_ (_26882_[11], _22825_, _22762_);
  and _27377_ (_22826_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not _27378_ (_22827_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor _27379_ (_22828_, _22770_, _22827_);
  or _27380_ (_22829_, _22828_, _22826_);
  and _27381_ (_26882_[12], _22829_, _22762_);
  and _27382_ (_22830_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not _27383_ (_22832_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _27384_ (_22833_, _22770_, _22832_);
  or _27385_ (_22834_, _22833_, _22830_);
  and _27386_ (_26882_[13], _22834_, _22762_);
  and _27387_ (_22836_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not _27388_ (_22837_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _27389_ (_22838_, _22770_, _22837_);
  or _27390_ (_22839_, _22838_, _22836_);
  and _27391_ (_26882_[14], _22839_, _22762_);
  and _27392_ (_22840_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _27393_ (_22841_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27394_ (_22842_, _22770_, _22841_);
  or _27395_ (_22843_, _22842_, _22840_);
  and _27396_ (_26883_[0], _22843_, _22762_);
  and _27397_ (_22844_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _27398_ (_22845_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _27399_ (_22846_, _22770_, _22845_);
  or _27400_ (_22847_, _22846_, _22844_);
  and _27401_ (_26883_[1], _22847_, _22762_);
  and _27402_ (_22848_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _27403_ (_22849_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _27404_ (_22850_, _22770_, _22849_);
  or _27405_ (_22852_, _22850_, _22848_);
  and _27406_ (_26883_[2], _22852_, _22762_);
  and _27407_ (_22853_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _27408_ (_22854_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _27409_ (_22855_, _22770_, _22854_);
  or _27410_ (_22857_, _22855_, _22853_);
  and _27411_ (_26883_[3], _22857_, _22762_);
  or _27412_ (_22859_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nand _27413_ (_22860_, _22770_, _22794_);
  and _27414_ (_22861_, _22860_, _22762_);
  and _27415_ (_26883_[4], _22861_, _22859_);
  and _27416_ (_22862_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not _27417_ (_22864_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _27418_ (_22865_, _22770_, _22864_);
  or _27419_ (_22867_, _22865_, _22862_);
  and _27420_ (_26883_[5], _22867_, _22762_);
  and _27421_ (_22868_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not _27422_ (_22869_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _27423_ (_22870_, _22770_, _22869_);
  or _27424_ (_22871_, _22870_, _22868_);
  and _27425_ (_26883_[6], _22871_, _22762_);
  and _27426_ (_22872_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not _27427_ (_22874_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _27428_ (_22875_, _22770_, _22874_);
  or _27429_ (_22876_, _22875_, _22872_);
  and _27430_ (_26883_[7], _22876_, _22762_);
  or _27431_ (_22877_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nand _27432_ (_22878_, _22770_, _22810_);
  and _27433_ (_22879_, _22878_, _22762_);
  and _27434_ (_26883_[8], _22879_, _22877_);
  and _27435_ (_22881_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  not _27436_ (_22882_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _27437_ (_22883_, _22770_, _22882_);
  or _27438_ (_22884_, _22883_, _22881_);
  and _27439_ (_26883_[9], _22884_, _22762_);
  and _27440_ (_22885_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  not _27441_ (_22886_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _27442_ (_22887_, _22770_, _22886_);
  or _27443_ (_22888_, _22887_, _22885_);
  and _27444_ (_26883_[10], _22888_, _22762_);
  and _27445_ (_22889_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not _27446_ (_22890_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _27447_ (_22891_, _22770_, _22890_);
  or _27448_ (_22892_, _22891_, _22889_);
  and _27449_ (_26883_[11], _22892_, _22762_);
  or _27450_ (_22893_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nand _27451_ (_22894_, _22770_, _22827_);
  and _27452_ (_22895_, _22894_, _22762_);
  and _27453_ (_26883_[12], _22895_, _22893_);
  and _27454_ (_22896_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not _27455_ (_22897_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _27456_ (_22899_, _22770_, _22897_);
  or _27457_ (_22900_, _22899_, _22896_);
  and _27458_ (_26883_[13], _22900_, _22762_);
  or _27459_ (_22901_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nand _27460_ (_22903_, _22770_, _22837_);
  and _27461_ (_22904_, _22903_, _22762_);
  and _27462_ (_26883_[14], _22904_, _22901_);
  and _27463_ (_22905_, \oc8051_top_1.oc8051_decoder1.wr , _22766_);
  not _27464_ (_22906_, _22905_);
  not _27465_ (_22907_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _27466_ (_22908_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _22766_);
  and _27467_ (_22909_, _22908_, _22907_);
  and _27468_ (_22910_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and _27469_ (_22912_, _22910_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _27470_ (_22913_, _22912_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _27471_ (_22914_, _22913_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _27472_ (_22915_, _22914_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _27473_ (_22917_, _22915_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and _27474_ (_22918_, _22917_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  not _27475_ (_22919_, _22918_);
  and _27476_ (_22920_, _22909_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  or _27477_ (_22921_, _22917_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and _27478_ (_22922_, _22921_, _22920_);
  and _27479_ (_22923_, _22922_, _22919_);
  not _27480_ (_22924_, _22923_);
  and _27481_ (_22926_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _27482_ (_22927_, _22926_, _22908_);
  not _27483_ (_22928_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _27484_ (_22929_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _22766_);
  and _27485_ (_22930_, _22929_, _22928_);
  and _27486_ (_22931_, _22930_, _22907_);
  and _27487_ (_22932_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor _27488_ (_22934_, _22932_, _22927_);
  nor _27489_ (_22935_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _27490_ (_22937_, _22935_, _22908_);
  and _27491_ (_22938_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and _27492_ (_22939_, _22930_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _27493_ (_22940_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor _27494_ (_22941_, _22940_, _22938_);
  and _27495_ (_22942_, _22941_, _22934_);
  nand _27496_ (_22943_, _22942_, _22924_);
  not _27497_ (_22944_, _22943_);
  nor _27498_ (_22945_, _22944_, _22909_);
  nor _27499_ (_22946_, _22945_, _22906_);
  not _27500_ (_22947_, _22946_);
  not _27501_ (_22948_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _27502_ (_22949_, _22943_, _22948_);
  nor _27503_ (_22950_, _22913_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not _27504_ (_22951_, _22950_);
  not _27505_ (_22952_, _22920_);
  nor _27506_ (_22953_, _22952_, _22914_);
  and _27507_ (_22954_, _22953_, _22951_);
  not _27508_ (_22956_, _22954_);
  and _27509_ (_22957_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor _27510_ (_22958_, _22957_, _22927_);
  and _27511_ (_22960_, _22935_, _22928_);
  or _27512_ (_22961_, _22960_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _27513_ (_22962_, _22961_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and _27514_ (_22963_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _27515_ (_22964_, _22963_, _22962_);
  and _27516_ (_22966_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not _27517_ (_22967_, _22966_);
  and _27518_ (_22968_, _22967_, _22964_);
  and _27519_ (_22969_, _22968_, _22958_);
  and _27520_ (_22970_, _22969_, _22956_);
  not _27521_ (_22971_, _22970_);
  and _27522_ (_22972_, _22971_, _22949_);
  nor _27523_ (_22973_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _27524_ (_22974_, _22973_, _22910_);
  and _27525_ (_22975_, _22974_, _22920_);
  and _27526_ (_22976_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor _27527_ (_22977_, _22976_, _22975_);
  and _27528_ (_22978_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and _27529_ (_22979_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and _27530_ (_22980_, _22961_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or _27531_ (_22981_, _22980_, _22979_);
  nor _27532_ (_22982_, _22981_, _22978_);
  and _27533_ (_22983_, _22982_, _22977_);
  nor _27534_ (_22984_, _22983_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _27535_ (_22985_, _22984_, _22972_);
  nor _27536_ (_22986_, _22985_, _22947_);
  nor _27537_ (_22987_, _22912_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _27538_ (_22989_, _22987_, _22913_);
  and _27539_ (_22990_, _22989_, _22920_);
  not _27540_ (_22991_, _22990_);
  and _27541_ (_22992_, _22961_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and _27542_ (_22994_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _27543_ (_22995_, _22994_, _22992_);
  and _27544_ (_22996_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and _27545_ (_22997_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor _27546_ (_22999_, _22997_, _22996_);
  and _27547_ (_23000_, _22999_, _22995_);
  and _27548_ (_23002_, _23000_, _22991_);
  not _27549_ (_23003_, _23002_);
  and _27550_ (_23004_, _23003_, _22949_);
  and _27551_ (_23005_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and _27552_ (_23006_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor _27553_ (_23008_, _23006_, _23005_);
  and _27554_ (_23009_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  not _27555_ (_23011_, _23009_);
  not _27556_ (_23012_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _27557_ (_23014_, _22920_, _23012_);
  and _27558_ (_23015_, _22961_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _27559_ (_23016_, _23015_, _23014_);
  and _27560_ (_23017_, _23016_, _23011_);
  and _27561_ (_23018_, _23017_, _23008_);
  nor _27562_ (_23019_, _23018_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _27563_ (_23020_, _23019_, _23004_);
  and _27564_ (_23021_, _23020_, _22986_);
  nor _27565_ (_23022_, _22915_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _27566_ (_23023_, _23022_);
  nor _27567_ (_23024_, _22952_, _22917_);
  and _27568_ (_23025_, _23024_, _23023_);
  not _27569_ (_23026_, _23025_);
  and _27570_ (_23027_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor _27571_ (_23028_, _23027_, _22927_);
  and _27572_ (_23029_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _27573_ (_23030_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor _27574_ (_23031_, _23030_, _23029_);
  and _27575_ (_23033_, _23031_, _23028_);
  and _27576_ (_23034_, _23033_, _23026_);
  not _27577_ (_23035_, _23034_);
  and _27578_ (_23036_, _23035_, _22949_);
  nor _27579_ (_23038_, _23002_, _22949_);
  nor _27580_ (_23039_, _23038_, _23036_);
  nor _27581_ (_23040_, _23039_, _22947_);
  nor _27582_ (_23041_, _22914_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _27583_ (_23042_, _23041_);
  nor _27584_ (_23043_, _22952_, _22915_);
  and _27585_ (_23044_, _23043_, _23042_);
  not _27586_ (_23045_, _23044_);
  and _27587_ (_23046_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor _27588_ (_23047_, _23046_, _22927_);
  and _27589_ (_23048_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _27590_ (_23049_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nor _27591_ (_23050_, _23049_, _23048_);
  and _27592_ (_23051_, _23050_, _23047_);
  and _27593_ (_23052_, _23051_, _23045_);
  not _27594_ (_23053_, _23052_);
  and _27595_ (_23054_, _23053_, _22949_);
  nor _27596_ (_23055_, _22910_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _27597_ (_23056_, _23055_, _22912_);
  and _27598_ (_23057_, _23056_, _22920_);
  and _27599_ (_23058_, _22937_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _27600_ (_23059_, _23058_, _23057_);
  and _27601_ (_23060_, _22939_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and _27602_ (_23061_, _22931_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and _27603_ (_23062_, _22961_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _27604_ (_23063_, _23062_, _23061_);
  nor _27605_ (_23064_, _23063_, _23060_);
  and _27606_ (_23065_, _23064_, _23059_);
  nor _27607_ (_23066_, _23065_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _27608_ (_23067_, _23066_, _23054_);
  and _27609_ (_23068_, _23067_, _23040_);
  and _27610_ (_23069_, _23068_, _23021_);
  nor _27611_ (_23070_, _22970_, _22949_);
  and _27612_ (_23071_, _23070_, _22946_);
  and _27613_ (_23072_, _23071_, _23053_);
  nor _27614_ (_23073_, _23035_, _22943_);
  nor _27615_ (_23074_, _23073_, _22949_);
  not _27616_ (_23075_, _23074_);
  and _27617_ (_23076_, _23075_, _23072_);
  and _27618_ (_23077_, _23076_, _23069_);
  nor _27619_ (_23078_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _27620_ (_23079_, \oc8051_top_1.oc8051_ram_top1.bit_select [2], \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand _27621_ (_23080_, _23079_, _23078_);
  and _27622_ (_23081_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _22766_);
  and _27623_ (_23082_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _22766_);
  nor _27624_ (_23083_, _23082_, _23081_);
  not _27625_ (_23084_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _27626_ (_23085_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _22766_);
  and _27627_ (_23086_, _23085_, _23084_);
  and _27628_ (_23087_, _23086_, _23083_);
  not _27629_ (_23088_, _23087_);
  not _27630_ (_23089_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _27631_ (_23090_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not _27632_ (_23091_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand _27633_ (_23092_, _23091_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _27634_ (_23093_, _23092_, _23090_);
  or _27635_ (_23094_, _23093_, _23089_);
  not _27636_ (_23095_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _27637_ (_23096_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand _27638_ (_23097_, _23096_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _27639_ (_23098_, _23097_, _23095_);
  and _27640_ (_23099_, _23098_, _23094_);
  not _27641_ (_23100_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  or _27642_ (_23101_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _27643_ (_23102_, _23101_, _23091_);
  or _27644_ (_23103_, _23102_, _23100_);
  not _27645_ (_23104_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  or _27646_ (_23105_, _23092_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _27647_ (_23106_, _23105_, _23104_);
  and _27648_ (_23107_, _23106_, _23103_);
  and _27649_ (_23108_, _23107_, _23099_);
  or _27650_ (_23109_, _23101_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  not _27651_ (_23110_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _27652_ (_23111_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _23110_);
  or _27653_ (_23112_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not _27654_ (_23113_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or _27655_ (_23114_, _23113_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and _27656_ (_23115_, _23114_, _23112_);
  or _27657_ (_23116_, _23115_, _23111_);
  nand _27658_ (_23117_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _23110_);
  or _27659_ (_23118_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand _27660_ (_23120_, _23118_, _23116_);
  or _27661_ (_23121_, _23120_, _23109_);
  and _27662_ (_23122_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _27663_ (_23123_, _23122_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _27664_ (_23124_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  not _27665_ (_23126_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nand _27666_ (_23127_, _23122_, _23090_);
  or _27667_ (_23128_, _23127_, _23126_);
  and _27668_ (_23129_, _23128_, _23124_);
  and _27669_ (_23130_, _23129_, _23121_);
  and _27670_ (_23131_, _23130_, _23108_);
  or _27671_ (_23132_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _27672_ (_23133_, _23132_, _23120_);
  and _27673_ (_23134_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _27674_ (_23135_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not _27675_ (_23137_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand _27676_ (_23138_, _23137_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nor _27677_ (_23139_, _23138_, _23126_);
  nor _27678_ (_23140_, _23139_, _23135_);
  and _27679_ (_23141_, _23140_, _23133_);
  not _27680_ (_23142_, _23141_);
  and _27681_ (_23143_, _23142_, _23131_);
  nor _27682_ (_23144_, _23141_, _23131_);
  and _27683_ (_23145_, _23141_, _23131_);
  nor _27684_ (_23146_, _23145_, _23144_);
  not _27685_ (_23147_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _27686_ (_23148_, _23093_, _23147_);
  not _27687_ (_23149_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _27688_ (_23150_, _23097_, _23149_);
  and _27689_ (_23151_, _23150_, _23148_);
  not _27690_ (_23152_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  or _27691_ (_23153_, _23102_, _23152_);
  not _27692_ (_23154_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or _27693_ (_23155_, _23105_, _23154_);
  and _27694_ (_23156_, _23155_, _23153_);
  and _27695_ (_23157_, _23156_, _23151_);
  or _27696_ (_23158_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  or _27697_ (_23159_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _23113_);
  and _27698_ (_23160_, _23159_, _23158_);
  or _27699_ (_23161_, _23160_, _23111_);
  or _27700_ (_23163_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _27701_ (_23164_, _23163_, _23161_);
  or _27702_ (_23165_, _23164_, _23109_);
  not _27703_ (_23166_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _27704_ (_23167_, _23127_, _23166_);
  nand _27705_ (_23168_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and _27706_ (_23169_, _23168_, _23167_);
  and _27707_ (_23170_, _23169_, _23165_);
  and _27708_ (_23171_, _23170_, _23157_);
  or _27709_ (_23172_, _23164_, _23132_);
  nand _27710_ (_23173_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or _27711_ (_23174_, _23138_, _23166_);
  and _27712_ (_23175_, _23174_, _23173_);
  nand _27713_ (_23177_, _23175_, _23172_);
  nor _27714_ (_23178_, _23177_, _23171_);
  not _27715_ (_23179_, _23177_);
  nor _27716_ (_23180_, _23179_, _23171_);
  and _27717_ (_23181_, _23179_, _23171_);
  nor _27718_ (_23182_, _23181_, _23180_);
  not _27719_ (_23183_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or _27720_ (_23184_, _23093_, _23183_);
  not _27721_ (_23185_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _27722_ (_23186_, _23097_, _23185_);
  and _27723_ (_23187_, _23186_, _23184_);
  not _27724_ (_23188_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  or _27725_ (_23190_, _23102_, _23188_);
  not _27726_ (_23191_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or _27727_ (_23192_, _23105_, _23191_);
  and _27728_ (_23193_, _23192_, _23190_);
  and _27729_ (_23194_, _23193_, _23187_);
  or _27730_ (_23195_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  or _27731_ (_23196_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _23113_);
  and _27732_ (_23197_, _23196_, _23195_);
  or _27733_ (_23198_, _23197_, _23111_);
  or _27734_ (_23199_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _27735_ (_23200_, _23199_, _23198_);
  or _27736_ (_23201_, _23200_, _23109_);
  not _27737_ (_23202_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _27738_ (_23203_, _23127_, _23202_);
  nand _27739_ (_23204_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and _27740_ (_23205_, _23204_, _23203_);
  and _27741_ (_23206_, _23205_, _23201_);
  nand _27742_ (_23208_, _23206_, _23194_);
  or _27743_ (_23209_, _23200_, _23132_);
  nand _27744_ (_23211_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or _27745_ (_23212_, _23138_, _23202_);
  and _27746_ (_23213_, _23212_, _23211_);
  and _27747_ (_23214_, _23213_, _23209_);
  and _27748_ (_23215_, _23214_, _23208_);
  nand _27749_ (_23216_, _23213_, _23209_);
  and _27750_ (_23217_, _23216_, _23208_);
  nor _27751_ (_23218_, _23216_, _23208_);
  nor _27752_ (_23219_, _23218_, _23217_);
  not _27753_ (_23220_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or _27754_ (_23221_, _23093_, _23220_);
  not _27755_ (_23222_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _27756_ (_23223_, _23097_, _23222_);
  and _27757_ (_23224_, _23223_, _23221_);
  not _27758_ (_23225_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  or _27759_ (_23226_, _23102_, _23225_);
  not _27760_ (_23227_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or _27761_ (_23228_, _23105_, _23227_);
  and _27762_ (_23229_, _23228_, _23226_);
  and _27763_ (_23230_, _23229_, _23224_);
  or _27764_ (_23231_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or _27765_ (_23232_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _23113_);
  and _27766_ (_23233_, _23232_, _23231_);
  or _27767_ (_23235_, _23233_, _23111_);
  or _27768_ (_23236_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _27769_ (_23237_, _23236_, _23235_);
  or _27770_ (_23238_, _23237_, _23109_);
  not _27771_ (_23239_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _27772_ (_23240_, _23127_, _23239_);
  nand _27773_ (_23241_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and _27774_ (_23242_, _23241_, _23240_);
  and _27775_ (_23243_, _23242_, _23238_);
  and _27776_ (_23244_, _23243_, _23230_);
  or _27777_ (_23245_, _23237_, _23132_);
  nand _27778_ (_23246_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or _27779_ (_23247_, _23138_, _23239_);
  and _27780_ (_23249_, _23247_, _23246_);
  nand _27781_ (_23250_, _23249_, _23245_);
  and _27782_ (_23251_, _23250_, _23244_);
  nor _27783_ (_23252_, _23251_, _23219_);
  nor _27784_ (_23253_, _23252_, _23215_);
  nor _27785_ (_23254_, _23253_, _23182_);
  nor _27786_ (_23256_, _23254_, _23178_);
  and _27787_ (_23257_, _23253_, _23182_);
  nor _27788_ (_23258_, _23257_, _23254_);
  not _27789_ (_23259_, _23258_);
  and _27790_ (_23260_, _23251_, _23219_);
  nor _27791_ (_23261_, _23260_, _23252_);
  not _27792_ (_23262_, _23261_);
  and _27793_ (_23263_, _23249_, _23245_);
  nor _27794_ (_23264_, _23263_, _23244_);
  and _27795_ (_23265_, _23263_, _23244_);
  nor _27796_ (_23266_, _23265_, _23264_);
  not _27797_ (_23267_, _23266_);
  not _27798_ (_23268_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _27799_ (_23269_, _23093_, _23268_);
  not _27800_ (_23270_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _27801_ (_23271_, _23097_, _23270_);
  and _27802_ (_23272_, _23271_, _23269_);
  not _27803_ (_23273_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  or _27804_ (_23274_, _23102_, _23273_);
  not _27805_ (_23275_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or _27806_ (_23276_, _23105_, _23275_);
  and _27807_ (_23277_, _23276_, _23274_);
  and _27808_ (_23278_, _23277_, _23272_);
  or _27809_ (_23279_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or _27810_ (_23280_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _23113_);
  and _27811_ (_23281_, _23280_, _23279_);
  or _27812_ (_23282_, _23281_, _23111_);
  or _27813_ (_23283_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _27814_ (_23284_, _23283_, _23282_);
  or _27815_ (_23285_, _23284_, _23109_);
  nand _27816_ (_23286_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  not _27817_ (_23287_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _27818_ (_23288_, _23127_, _23287_);
  and _27819_ (_23289_, _23288_, _23286_);
  and _27820_ (_23290_, _23289_, _23285_);
  and _27821_ (_23291_, _23290_, _23278_);
  or _27822_ (_23292_, _23284_, _23132_);
  nand _27823_ (_23293_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or _27824_ (_23294_, _23138_, _23287_);
  and _27825_ (_23295_, _23294_, _23293_);
  and _27826_ (_23296_, _23295_, _23292_);
  and _27827_ (_23298_, _23296_, _23291_);
  nor _27828_ (_23299_, _23296_, _23291_);
  nor _27829_ (_23301_, _23299_, _23298_);
  not _27830_ (_23302_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  or _27831_ (_23303_, _23102_, _23302_);
  not _27832_ (_23304_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _27833_ (_23305_, _23127_, _23304_);
  and _27834_ (_23306_, _23305_, _23303_);
  not _27835_ (_23307_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _27836_ (_23308_, _23093_, _23307_);
  not _27837_ (_23309_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _27838_ (_23310_, _23097_, _23309_);
  and _27839_ (_23311_, _23310_, _23308_);
  and _27840_ (_23312_, _23311_, _23306_);
  or _27841_ (_23313_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  or _27842_ (_23314_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _23113_);
  and _27843_ (_23315_, _23314_, _23313_);
  or _27844_ (_23316_, _23315_, _23111_);
  or _27845_ (_23317_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _27846_ (_23318_, _23317_, _23316_);
  or _27847_ (_23320_, _23318_, _23109_);
  nand _27848_ (_23321_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  not _27849_ (_23322_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or _27850_ (_23323_, _23105_, _23322_);
  and _27851_ (_23324_, _23323_, _23321_);
  and _27852_ (_23325_, _23324_, _23320_);
  nand _27853_ (_23326_, _23325_, _23312_);
  or _27854_ (_23327_, _23318_, _23132_);
  nand _27855_ (_23329_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or _27856_ (_23330_, _23138_, _23304_);
  and _27857_ (_23331_, _23330_, _23329_);
  nand _27858_ (_23332_, _23331_, _23327_);
  and _27859_ (_23333_, _23332_, _23326_);
  nor _27860_ (_23334_, _23332_, _23326_);
  nor _27861_ (_23335_, _23334_, _23333_);
  not _27862_ (_23336_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _27863_ (_23337_, _23093_, _23336_);
  not _27864_ (_23338_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _27865_ (_23339_, _23097_, _23338_);
  and _27866_ (_23340_, _23339_, _23337_);
  not _27867_ (_23341_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  or _27868_ (_23342_, _23102_, _23341_);
  not _27869_ (_23343_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or _27870_ (_23344_, _23105_, _23343_);
  and _27871_ (_23345_, _23344_, _23342_);
  and _27872_ (_23346_, _23345_, _23340_);
  or _27873_ (_23347_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or _27874_ (_23348_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _23113_);
  and _27875_ (_23349_, _23348_, _23347_);
  or _27876_ (_23350_, _23349_, _23111_);
  or _27877_ (_23351_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _27878_ (_23352_, _23351_, _23350_);
  or _27879_ (_23353_, _23352_, _23109_);
  nand _27880_ (_23354_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  not _27881_ (_23355_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _27882_ (_23356_, _23127_, _23355_);
  and _27883_ (_23357_, _23356_, _23354_);
  and _27884_ (_23358_, _23357_, _23353_);
  nand _27885_ (_23359_, _23358_, _23346_);
  or _27886_ (_23360_, _23352_, _23132_);
  nand _27887_ (_23361_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or _27888_ (_23362_, _23138_, _23355_);
  and _27889_ (_23363_, _23362_, _23361_);
  nand _27890_ (_23364_, _23363_, _23360_);
  and _27891_ (_23365_, _23364_, _23359_);
  nor _27892_ (_23366_, _23364_, _23359_);
  nor _27893_ (_23367_, _23366_, _23365_);
  not _27894_ (_23368_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _27895_ (_23369_, _23093_, _23368_);
  not _27896_ (_23370_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _27897_ (_23371_, _23097_, _23370_);
  nor _27898_ (_23372_, _23371_, _23369_);
  not _27899_ (_23373_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor _27900_ (_23374_, _23102_, _23373_);
  not _27901_ (_23375_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor _27902_ (_23376_, _23105_, _23375_);
  nor _27903_ (_23377_, _23376_, _23374_);
  and _27904_ (_23378_, _23377_, _23372_);
  or _27905_ (_23379_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or _27906_ (_23380_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _23113_);
  and _27907_ (_23381_, _23380_, _23379_);
  or _27908_ (_23382_, _23381_, _23111_);
  or _27909_ (_23383_, _23117_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _27910_ (_23384_, _23383_, _23382_);
  or _27911_ (_23385_, _23384_, _23109_);
  and _27912_ (_23386_, _23123_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  not _27913_ (_23387_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _27914_ (_23389_, _23127_, _23387_);
  nor _27915_ (_23390_, _23389_, _23386_);
  and _27916_ (_23391_, _23390_, _23385_);
  and _27917_ (_23392_, _23391_, _23378_);
  or _27918_ (_23393_, _23384_, _23132_);
  nand _27919_ (_23394_, _23134_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  or _27920_ (_23395_, _23138_, _23387_);
  and _27921_ (_23396_, _23395_, _23394_);
  nand _27922_ (_23397_, _23396_, _23393_);
  and _27923_ (_23398_, _23397_, _23392_);
  nor _27924_ (_23399_, _23398_, _23367_);
  and _27925_ (_23400_, _23363_, _23360_);
  and _27926_ (_23401_, _23400_, _23359_);
  nor _27927_ (_23402_, _23401_, _23399_);
  nor _27928_ (_23403_, _23402_, _23335_);
  and _27929_ (_23404_, _23331_, _23327_);
  and _27930_ (_23405_, _23404_, _23326_);
  nor _27931_ (_23407_, _23405_, _23403_);
  nor _27932_ (_23408_, _23407_, _23301_);
  and _27933_ (_23409_, _23407_, _23301_);
  nor _27934_ (_23411_, _23409_, _23408_);
  and _27935_ (_23412_, _23402_, _23335_);
  nor _27936_ (_23413_, _23412_, _23403_);
  not _27937_ (_23414_, _23413_);
  and _27938_ (_23415_, _23398_, _23367_);
  nor _27939_ (_23416_, _23415_, _23399_);
  not _27940_ (_23417_, _23416_);
  and _27941_ (_23418_, _23396_, _23393_);
  nor _27942_ (_23419_, _23418_, _23392_);
  and _27943_ (_23420_, _23418_, _23392_);
  nor _27944_ (_23421_, _23420_, _23419_);
  not _27945_ (_23422_, _23421_);
  nor _27946_ (_23423_, _23117_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not _27947_ (_23424_, _23423_);
  not _27948_ (_23425_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and _27949_ (_23427_, _23425_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _27950_ (_23428_, _23427_, _23160_);
  and _27951_ (_23429_, _23428_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _27952_ (_23430_, _23233_, _23078_);
  and _27953_ (_23431_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _27954_ (_23432_, _23431_, _23115_);
  not _27955_ (_23433_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _27956_ (_23434_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _23433_);
  nand _27957_ (_23435_, _23434_, _23197_);
  and _27958_ (_23436_, _23435_, _23432_);
  and _27959_ (_23437_, _23436_, _23430_);
  nand _27960_ (_23438_, _23437_, _23429_);
  not _27961_ (_23439_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _27962_ (_23440_, _23427_, _23315_);
  and _27963_ (_23441_, _23440_, _23439_);
  nand _27964_ (_23442_, _23434_, _23349_);
  nand _27965_ (_23443_, _23431_, _23281_);
  nand _27966_ (_23444_, _23381_, _23078_);
  and _27967_ (_23445_, _23444_, _23443_);
  and _27968_ (_23446_, _23445_, _23442_);
  nand _27969_ (_23447_, _23446_, _23441_);
  nand _27970_ (_23448_, _23447_, _23438_);
  nand _27971_ (_23449_, _23448_, _23117_);
  and _27972_ (_23450_, _23449_, _23424_);
  and _27973_ (_23451_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _27974_ (_23452_, _23451_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _27975_ (_23453_, _23452_);
  and _27976_ (_23454_, _23453_, _23450_);
  and _27977_ (_23455_, _23453_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _27978_ (_23456_, _23455_, _23454_);
  and _27979_ (_23457_, _23456_, _23422_);
  and _27980_ (_23458_, _23457_, _23417_);
  and _27981_ (_23459_, _23458_, _23414_);
  not _27982_ (_23460_, _23459_);
  nor _27983_ (_23461_, _23460_, _23411_);
  nand _27984_ (_23462_, _23295_, _23292_);
  or _27985_ (_23463_, _23462_, _23291_);
  and _27986_ (_23464_, _23462_, _23291_);
  or _27987_ (_23465_, _23407_, _23464_);
  and _27988_ (_23466_, _23465_, _23463_);
  or _27989_ (_23467_, _23466_, _23461_);
  and _27990_ (_23468_, _23467_, _23267_);
  and _27991_ (_23469_, _23468_, _23262_);
  and _27992_ (_23470_, _23469_, _23259_);
  nor _27993_ (_23471_, _23470_, _23256_);
  nor _27994_ (_23472_, _23471_, _23146_);
  nor _27995_ (_23473_, _23472_, _23143_);
  nor _27996_ (_23474_, _23473_, _23088_);
  not _27997_ (_23475_, _23474_);
  not _27998_ (_23476_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _27999_ (_23478_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _22766_);
  and _28000_ (_23479_, _23478_, _23476_);
  and _28001_ (_23480_, _23479_, _23083_);
  not _28002_ (_23481_, _23480_);
  not _28003_ (_23482_, _23144_);
  not _28004_ (_23483_, _23146_);
  not _28005_ (_23484_, _23335_);
  and _28006_ (_23485_, _23419_, _23367_);
  nor _28007_ (_23486_, _23485_, _23365_);
  nor _28008_ (_23487_, _23486_, _23484_);
  nor _28009_ (_23488_, _23487_, _23333_);
  nor _28010_ (_23489_, _23488_, _23301_);
  and _28011_ (_23490_, _23488_, _23301_);
  nor _28012_ (_23491_, _23490_, _23489_);
  and _28013_ (_23492_, _23456_, _23421_);
  and _28014_ (_23493_, _23492_, _23367_);
  and _28015_ (_23494_, _23486_, _23484_);
  nor _28016_ (_23495_, _23494_, _23487_);
  and _28017_ (_23496_, _23495_, _23493_);
  not _28018_ (_23497_, _23496_);
  nor _28019_ (_23498_, _23497_, _23491_);
  nor _28020_ (_23499_, _23488_, _23298_);
  or _28021_ (_23500_, _23499_, _23299_);
  or _28022_ (_23501_, _23500_, _23498_);
  and _28023_ (_23502_, _23501_, _23266_);
  and _28024_ (_23503_, _23502_, _23219_);
  not _28025_ (_23505_, _23182_);
  and _28026_ (_23506_, _23264_, _23219_);
  nor _28027_ (_23508_, _23506_, _23217_);
  nor _28028_ (_23509_, _23508_, _23505_);
  and _28029_ (_23510_, _23508_, _23505_);
  nor _28030_ (_23511_, _23510_, _23509_);
  and _28031_ (_23512_, _23511_, _23503_);
  not _28032_ (_23514_, _23512_);
  nor _28033_ (_23515_, _23509_, _23180_);
  and _28034_ (_23516_, _23515_, _23514_);
  or _28035_ (_23518_, _23516_, _23483_);
  and _28036_ (_23519_, _23518_, _23482_);
  nor _28037_ (_23520_, _23519_, _23481_);
  nor _28038_ (_23521_, _23455_, _23454_);
  not _28039_ (_23522_, _23208_);
  and _28040_ (_23523_, _23522_, _23171_);
  not _28041_ (_23524_, _23523_);
  not _28042_ (_23525_, _23244_);
  not _28043_ (_23526_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _28044_ (_23527_, _23082_, _23526_);
  and _28045_ (_23528_, _23527_, _23479_);
  nor _28046_ (_23529_, _23359_, _23326_);
  nor _28047_ (_23530_, _23529_, _23291_);
  and _28048_ (_23531_, _23530_, _23528_);
  and _28049_ (_23532_, _23531_, _23525_);
  nor _28050_ (_23533_, _23532_, _23524_);
  nand _28051_ (_23534_, _23533_, _23521_);
  not _28052_ (_23535_, _23533_);
  not _28053_ (_23536_, _23131_);
  and _28054_ (_23537_, _23456_, _23536_);
  and _28055_ (_23538_, _23537_, _23535_);
  not _28056_ (_23539_, _23528_);
  and _28057_ (_23540_, _23521_, _23131_);
  or _28058_ (_23541_, _23540_, _23539_);
  nor _28059_ (_23542_, _23541_, _23538_);
  and _28060_ (_23543_, _23542_, _23534_);
  not _28061_ (_23544_, _23543_);
  nor _28062_ (_23545_, _23455_, _23450_);
  not _28063_ (_23546_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _28064_ (_23547_, _23081_, _23546_);
  and _28065_ (_23548_, _23547_, _23479_);
  nor _28066_ (_23549_, _23478_, _23085_);
  and _28067_ (_23550_, _23549_, _23547_);
  not _28068_ (_23551_, _23550_);
  nor _28069_ (_23552_, _23551_, _23454_);
  nor _28070_ (_23553_, _23552_, _23548_);
  nor _28071_ (_23555_, _23553_, _23545_);
  not _28072_ (_23556_, _23555_);
  and _28073_ (_23557_, _23527_, _23086_);
  and _28074_ (_23558_, _23557_, _23521_);
  not _28075_ (_23559_, _23558_);
  not _28076_ (_23560_, _23531_);
  not _28077_ (_23561_, _23450_);
  and _28078_ (_23562_, _23081_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _28079_ (_23563_, _23562_, _23549_);
  and _28080_ (_23564_, _23563_, _23455_);
  and _28081_ (_23565_, _23564_, _23561_);
  not _28082_ (_23567_, _23392_);
  and _28083_ (_23568_, _23562_, _23479_);
  and _28084_ (_23569_, _23568_, _23567_);
  and _28085_ (_23570_, _23085_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _28086_ (_23571_, _23570_, _23547_);
  and _28087_ (_23572_, _23571_, _23536_);
  nor _28088_ (_23574_, _23572_, _23569_);
  not _28089_ (_23575_, _23574_);
  nor _28090_ (_23576_, _23575_, _23565_);
  and _28091_ (_23577_, _23576_, _23560_);
  and _28092_ (_23578_, _23577_, _23559_);
  and _28093_ (_23579_, _23549_, _23083_);
  and _28094_ (_23580_, _23579_, _23456_);
  and _28095_ (_23581_, _23452_, _23450_);
  and _28096_ (_23582_, _23547_, _23086_);
  and _28097_ (_23583_, _23570_, _23527_);
  and _28098_ (_23584_, _23583_, _23450_);
  nor _28099_ (_23585_, _23584_, _23582_);
  nor _28100_ (_23587_, _23585_, _23581_);
  nor _28101_ (_23588_, _23587_, _23580_);
  and _28102_ (_23589_, _23588_, _23578_);
  and _28103_ (_23590_, _23589_, _23556_);
  and _28104_ (_23591_, _23590_, _23544_);
  not _28105_ (_23592_, _23591_);
  nor _28106_ (_23593_, _23592_, _23520_);
  and _28107_ (_23594_, _23593_, _23475_);
  nor _28108_ (_23595_, _23594_, _23080_);
  and _28109_ (_23596_, _23570_, _23083_);
  not _28110_ (_23597_, _23596_);
  and _28111_ (_23598_, _23479_, _23526_);
  and _28112_ (_23599_, _23549_, _23527_);
  nor _28113_ (_23600_, _23599_, _23598_);
  and _28114_ (_23601_, _23600_, _23597_);
  and _28115_ (_23602_, _23562_, _23476_);
  not _28116_ (_23603_, _23602_);
  and _28117_ (_23604_, _23547_, _23085_);
  nor _28118_ (_23605_, _23604_, _23579_);
  and _28119_ (_23606_, _23605_, _23603_);
  and _28120_ (_23607_, _23606_, _23601_);
  nor _28121_ (_23608_, _23607_, _23244_);
  and _28122_ (_23609_, _23562_, _23086_);
  not _28123_ (_23610_, _23326_);
  and _28124_ (_23611_, _23610_, _23291_);
  not _28125_ (_23612_, _23359_);
  and _28126_ (_23613_, _23392_, _23612_);
  and _28127_ (_23614_, _23613_, _23611_);
  or _28128_ (_23615_, _23614_, _23521_);
  not _28129_ (_23616_, _23291_);
  and _28130_ (_23617_, _23567_, _23359_);
  and _28131_ (_23618_, _23617_, _23326_);
  and _28132_ (_23619_, _23618_, _23616_);
  or _28133_ (_23621_, _23619_, _23456_);
  and _28134_ (_23622_, _23621_, _23615_);
  or _28135_ (_23623_, _23622_, _23525_);
  nand _28136_ (_23624_, _23622_, _23525_);
  and _28137_ (_23625_, _23624_, _23623_);
  and _28138_ (_23626_, _23625_, _23609_);
  and _28139_ (_23627_, _23570_, _23562_);
  or _28140_ (_23628_, _23521_, _23263_);
  or _28141_ (_23629_, _23456_, _23244_);
  nand _28142_ (_23630_, _23629_, _23628_);
  nand _28143_ (_23631_, _23630_, _23627_);
  and _28144_ (_23632_, _23550_, _23266_);
  and _28145_ (_23633_, _23583_, _23264_);
  not _28146_ (_23634_, _23548_);
  nor _28147_ (_23635_, _23634_, _23265_);
  and _28148_ (_23636_, _23557_, _23244_);
  or _28149_ (_23637_, _23636_, _23635_);
  or _28150_ (_23638_, _23637_, _23633_);
  nor _28151_ (_23639_, _23638_, _23632_);
  nand _28152_ (_23640_, _23639_, _23631_);
  or _28153_ (_23641_, _23640_, _23626_);
  or _28154_ (_23642_, _23641_, _23608_);
  and _28155_ (_23643_, _23642_, _22948_);
  and _28156_ (_23644_, _23078_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _28157_ (_23645_, _23233_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor _28158_ (_23646_, _23645_, _23644_);
  or _28159_ (_23647_, _23646_, _23643_);
  or _28160_ (_23648_, _23647_, _23595_);
  and _28161_ (_23649_, _23648_, _22946_);
  and _28162_ (_23651_, _23649_, _23077_);
  not _28163_ (_23652_, _23077_);
  and _28164_ (_23653_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  or _28165_ (_02714_, _23653_, _23651_);
  nor _28166_ (_23654_, _23067_, _22947_);
  and _28167_ (_23655_, _23654_, _23039_);
  and _28168_ (_23656_, _23655_, _23021_);
  nor _28169_ (_23657_, _23053_, _22949_);
  not _28170_ (_23658_, _23657_);
  and _28171_ (_23660_, _23658_, _22946_);
  nor _28172_ (_23661_, _23660_, _23071_);
  and _28173_ (_23662_, _23035_, _22943_);
  and _28174_ (_23663_, _23662_, _22946_);
  and _28175_ (_23664_, _23663_, _23661_);
  and _28176_ (_23665_, _23664_, _23656_);
  nand _28177_ (_23666_, _23431_, _23079_);
  nor _28178_ (_23667_, _23666_, _23594_);
  nand _28179_ (_23668_, _23431_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _28180_ (_23669_, _23115_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _28181_ (_23670_, _23669_, _23668_);
  nor _28182_ (_23671_, _23607_, _23131_);
  not _28183_ (_23672_, _23671_);
  and _28184_ (_23673_, _23614_, _23244_);
  and _28185_ (_23674_, _23673_, _23523_);
  nor _28186_ (_23675_, _23674_, _23521_);
  nand _28187_ (_23676_, _23619_, _23525_);
  or _28188_ (_23677_, _23676_, _23522_);
  or _28189_ (_23678_, _23677_, _23171_);
  and _28190_ (_23679_, _23678_, _23521_);
  nor _28191_ (_23680_, _23679_, _23675_);
  or _28192_ (_23681_, _23680_, _23131_);
  nand _28193_ (_23682_, _23680_, _23131_);
  nand _28194_ (_23683_, _23682_, _23681_);
  nand _28195_ (_23684_, _23683_, _23609_);
  and _28196_ (_23686_, _23456_, _23141_);
  not _28197_ (_23687_, _23686_);
  not _28198_ (_23688_, _23627_);
  nor _28199_ (_23689_, _23688_, _23540_);
  and _28200_ (_23690_, _23689_, _23687_);
  and _28201_ (_23691_, _23550_, _23146_);
  and _28202_ (_23692_, _23583_, _23144_);
  nor _28203_ (_23693_, _23634_, _23145_);
  and _28204_ (_23694_, _23557_, _23131_);
  or _28205_ (_23695_, _23694_, _23693_);
  or _28206_ (_23696_, _23695_, _23692_);
  nor _28207_ (_23697_, _23696_, _23691_);
  not _28208_ (_23699_, _23697_);
  nor _28209_ (_23700_, _23699_, _23690_);
  and _28210_ (_23701_, _23700_, _23684_);
  and _28211_ (_23702_, _23701_, _23672_);
  nor _28212_ (_23704_, _23702_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  or _28213_ (_23705_, _23704_, _23670_);
  or _28214_ (_23706_, _23705_, _23667_);
  and _28215_ (_23707_, _23706_, _22946_);
  and _28216_ (_23708_, _23707_, _23665_);
  not _28217_ (_23709_, _23665_);
  and _28218_ (_23710_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  or _28219_ (_27079_, _23710_, _23708_);
  not _28220_ (_23711_, _23594_);
  and _28221_ (_23712_, _23439_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _28222_ (_23713_, _23712_, _23431_);
  and _28223_ (_23714_, _23713_, _23711_);
  and _28224_ (_23715_, _23627_, _23462_);
  nor _28225_ (_23716_, _23618_, _23616_);
  or _28226_ (_23717_, _23716_, _23621_);
  nand _28227_ (_23718_, _23529_, _23392_);
  and _28228_ (_23719_, _23718_, _23616_);
  or _28229_ (_23720_, _23719_, _23614_);
  nand _28230_ (_23721_, _23720_, _23456_);
  nand _28231_ (_23722_, _23721_, _23717_);
  and _28232_ (_23724_, _23722_, _23609_);
  nor _28233_ (_23725_, _23724_, _23715_);
  nor _28234_ (_23726_, _23607_, _23291_);
  not _28235_ (_23727_, _23726_);
  and _28236_ (_23728_, _23550_, _23301_);
  not _28237_ (_23729_, _23728_);
  nor _28238_ (_23730_, _23634_, _23298_);
  not _28239_ (_23731_, _23730_);
  and _28240_ (_23732_, _23583_, _23299_);
  and _28241_ (_23733_, _23557_, _23291_);
  nor _28242_ (_23734_, _23733_, _23732_);
  and _28243_ (_23735_, _23734_, _23731_);
  and _28244_ (_23736_, _23735_, _23729_);
  and _28245_ (_23737_, _23736_, _23727_);
  nand _28246_ (_23738_, _23737_, _23725_);
  and _28247_ (_23739_, _23738_, _22948_);
  and _28248_ (_23740_, _23712_, _23425_);
  and _28249_ (_23741_, _23712_, _23433_);
  or _28250_ (_23742_, _23741_, _23079_);
  or _28251_ (_23743_, _23742_, _23740_);
  and _28252_ (_23744_, _23743_, _23281_);
  or _28253_ (_23745_, _23744_, _23739_);
  or _28254_ (_23746_, _23745_, _23714_);
  and _28255_ (_23747_, _23746_, _22946_);
  and _28256_ (_23748_, _23747_, _23077_);
  and _28257_ (_23749_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  or _28258_ (_09923_, _23749_, _23748_);
  nor _28259_ (_23750_, _23020_, _22947_);
  and _28260_ (_23751_, _23750_, _22986_);
  and _28261_ (_23752_, _23751_, _23655_);
  and _28262_ (_23753_, _23034_, _22943_);
  and _28263_ (_23754_, _23753_, _23072_);
  and _28264_ (_23755_, _23754_, _23752_);
  and _28265_ (_23756_, _23712_, _23078_);
  nand _28266_ (_23757_, _23756_, _23594_);
  nor _28267_ (_23758_, _23551_, _23419_);
  nor _28268_ (_23759_, _23758_, _23548_);
  or _28269_ (_23760_, _23759_, _23420_);
  and _28270_ (_23761_, _23583_, _23419_);
  and _28271_ (_23762_, _23557_, _23392_);
  nor _28272_ (_23764_, _23762_, _23761_);
  and _28273_ (_23765_, _23627_, _23397_);
  and _28274_ (_23766_, _23609_, _23392_);
  nor _28275_ (_23767_, _23766_, _23765_);
  nor _28276_ (_23768_, _23607_, _23392_);
  not _28277_ (_23769_, _23768_);
  and _28278_ (_23770_, _23769_, _23767_);
  and _28279_ (_23771_, _23770_, _23764_);
  and _28280_ (_23772_, _23771_, _23760_);
  nand _28281_ (_23773_, _23772_, _22948_);
  or _28282_ (_23774_, _23381_, _22948_);
  and _28283_ (_23775_, _23774_, _23773_);
  or _28284_ (_23776_, _23775_, _23756_);
  and _28285_ (_23777_, _23776_, _23757_);
  and _28286_ (_23778_, _23777_, _22946_);
  and _28287_ (_23779_, _23778_, _23755_);
  not _28288_ (_23780_, _23755_);
  and _28289_ (_23781_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  or _28290_ (_13798_, _23781_, _23779_);
  nor _28291_ (_23782_, _23750_, _22986_);
  nor _28292_ (_23783_, _23654_, _23040_);
  and _28293_ (_23784_, _23783_, _23782_);
  and _28294_ (_23785_, _23071_, _23052_);
  nor _28295_ (_23786_, _23034_, _22949_);
  and _28296_ (_23787_, _23786_, _22946_);
  and _28297_ (_23788_, _23787_, _22944_);
  and _28298_ (_23789_, _23788_, _23785_);
  and _28299_ (_23790_, _23789_, _23784_);
  nand _28300_ (_23791_, _23712_, _23427_);
  nor _28301_ (_23792_, _23791_, _23594_);
  and _28302_ (_23793_, _23627_, _23332_);
  not _28303_ (_23794_, _23613_);
  or _28304_ (_23795_, _23794_, _23521_);
  not _28305_ (_23796_, _23617_);
  or _28306_ (_23797_, _23796_, _23456_);
  and _28307_ (_23798_, _23797_, _23795_);
  nand _28308_ (_23799_, _23798_, _23610_);
  or _28309_ (_23800_, _23798_, _23610_);
  and _28310_ (_23801_, _23800_, _23609_);
  and _28311_ (_23802_, _23801_, _23799_);
  nor _28312_ (_23803_, _23802_, _23793_);
  and _28313_ (_23804_, _23550_, _23335_);
  nor _28314_ (_23805_, _23634_, _23334_);
  or _28315_ (_23806_, _23805_, _23804_);
  not _28316_ (_23807_, _23806_);
  and _28317_ (_23808_, _23583_, _23333_);
  and _28318_ (_23809_, _23557_, _23610_);
  nor _28319_ (_23810_, _23809_, _23808_);
  and _28320_ (_23811_, _23810_, _23807_);
  nor _28321_ (_23812_, _23607_, _23610_);
  not _28322_ (_23813_, _23812_);
  and _28323_ (_23814_, _23813_, _23811_);
  nand _28324_ (_23816_, _23814_, _23803_);
  and _28325_ (_23817_, _23816_, _22948_);
  or _28326_ (_23818_, _23713_, _23079_);
  or _28327_ (_23820_, _23818_, _23741_);
  and _28328_ (_23821_, _23820_, _23315_);
  or _28329_ (_23822_, _23821_, _23817_);
  or _28330_ (_23823_, _23822_, _23792_);
  and _28331_ (_23824_, _23823_, _22946_);
  and _28332_ (_23825_, _23824_, _23790_);
  not _28333_ (_23827_, _23790_);
  and _28334_ (_23828_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  or _28335_ (_16236_, _23828_, _23825_);
  and _28336_ (_23829_, _23790_, _23649_);
  and _28337_ (_23830_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  or _28338_ (_16455_, _23830_, _23829_);
  and _28339_ (_23831_, _23790_, _23747_);
  and _28340_ (_23832_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  or _28341_ (_22627_, _23832_, _23831_);
  and _28342_ (_23833_, _23754_, _23656_);
  and _28343_ (_23834_, _23833_, _23824_);
  not _28344_ (_23835_, _23833_);
  and _28345_ (_23836_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or _28346_ (_22643_, _23836_, _23834_);
  not _28347_ (_23837_, _22767_);
  not _28348_ (_23838_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _28349_ (_23839_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _28350_ (_23840_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _28351_ (_23841_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _28352_ (_23842_, _23841_, _23840_);
  and _28353_ (_23843_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _28354_ (_23844_, _23841_, _23840_);
  and _28355_ (_23845_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _28356_ (_23846_, _23841_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _28357_ (_23847_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _28358_ (_23848_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _28359_ (_23849_, _23848_, _23840_);
  and _28360_ (_23850_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _28361_ (_23851_, _23850_, _23847_);
  nor _28362_ (_23852_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _28363_ (_23853_, _23852_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _28364_ (_23854_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  not _28365_ (_23855_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _28366_ (_23856_, _23855_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _28367_ (_23857_, _23856_, _23840_);
  and _28368_ (_23858_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _28369_ (_23859_, _23858_, _23854_);
  nand _28370_ (_23860_, _23859_, _23851_);
  or _28371_ (_23861_, _23860_, _23845_);
  nor _28372_ (_23862_, _23861_, _23843_);
  and _28373_ (_23863_, _23862_, _23839_);
  and _28374_ (_23864_, _23863_, _23838_);
  nor _28375_ (_23865_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _23838_);
  nor _28376_ (_23866_, _23865_, _23864_);
  or _28377_ (_23867_, _23866_, _23837_);
  or _28378_ (_23868_, _22767_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _28379_ (_23869_, _23868_, _22762_);
  and _28380_ (_26864_[1], _23869_, _23867_);
  nand _28381_ (_23870_, _23712_, _23434_);
  nor _28382_ (_23871_, _23870_, _23594_);
  and _28383_ (_23872_, _23627_, _23364_);
  nor _28384_ (_23873_, _23617_, _23613_);
  nand _28385_ (_23874_, _23873_, _23456_);
  or _28386_ (_23875_, _23873_, _23456_);
  and _28387_ (_23876_, _23875_, _23609_);
  and _28388_ (_23877_, _23876_, _23874_);
  nor _28389_ (_23878_, _23877_, _23872_);
  nor _28390_ (_23879_, _23607_, _23612_);
  not _28391_ (_23880_, _23879_);
  and _28392_ (_23881_, _23550_, _23367_);
  not _28393_ (_23882_, _23881_);
  nor _28394_ (_23883_, _23634_, _23366_);
  not _28395_ (_23884_, _23883_);
  and _28396_ (_23885_, _23583_, _23365_);
  and _28397_ (_23886_, _23557_, _23612_);
  nor _28398_ (_23887_, _23886_, _23885_);
  and _28399_ (_23888_, _23887_, _23884_);
  and _28400_ (_23889_, _23888_, _23882_);
  and _28401_ (_23890_, _23889_, _23880_);
  nand _28402_ (_23892_, _23890_, _23878_);
  and _28403_ (_23893_, _23892_, _22948_);
  or _28404_ (_23894_, _23740_, _23818_);
  and _28405_ (_23895_, _23894_, _23349_);
  or _28406_ (_23896_, _23895_, _23893_);
  or _28407_ (_23897_, _23896_, _23871_);
  and _28408_ (_23898_, _23897_, _22946_);
  and _28409_ (_23899_, _23898_, _23833_);
  and _28410_ (_23900_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or _28411_ (_22722_, _23900_, _23899_);
  and _28412_ (_23901_, _23750_, _22985_);
  and _28413_ (_23902_, _23654_, _23040_);
  and _28414_ (_23903_, _23902_, _23901_);
  not _28415_ (_23904_, _23070_);
  and _28416_ (_23905_, _23660_, _23904_);
  and _28417_ (_23906_, _23905_, _23788_);
  and _28418_ (_23907_, _23906_, _23903_);
  and _28419_ (_23908_, _23907_, _23747_);
  not _28420_ (_23909_, _23907_);
  and _28421_ (_23910_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or _28422_ (_22746_, _23910_, _23908_);
  and _28423_ (_23911_, _23783_, _23751_);
  and _28424_ (_23912_, _23911_, _23789_);
  nand _28425_ (_23913_, _23434_, _23079_);
  nor _28426_ (_23914_, _23913_, _23594_);
  and _28427_ (_23915_, _23521_, _23522_);
  and _28428_ (_23916_, _23456_, _23214_);
  or _28429_ (_23917_, _23916_, _23688_);
  nor _28430_ (_23918_, _23917_, _23915_);
  or _28431_ (_23919_, _23676_, _23456_);
  nand _28432_ (_23920_, _23673_, _23456_);
  and _28433_ (_23921_, _23920_, _23919_);
  and _28434_ (_23922_, _23921_, _23522_);
  or _28435_ (_23923_, _23921_, _23522_);
  nand _28436_ (_23924_, _23923_, _23609_);
  nor _28437_ (_23925_, _23924_, _23922_);
  nor _28438_ (_23926_, _23925_, _23918_);
  and _28439_ (_23927_, _23550_, _23219_);
  and _28440_ (_23929_, _23583_, _23217_);
  nor _28441_ (_23930_, _23634_, _23218_);
  and _28442_ (_23932_, _23557_, _23522_);
  or _28443_ (_23933_, _23932_, _23930_);
  or _28444_ (_23934_, _23933_, _23929_);
  nor _28445_ (_23935_, _23934_, _23927_);
  nor _28446_ (_23936_, _23607_, _23522_);
  not _28447_ (_23937_, _23936_);
  and _28448_ (_23938_, _23937_, _23935_);
  nand _28449_ (_23939_, _23938_, _23926_);
  and _28450_ (_23940_, _23939_, _22948_);
  nand _28451_ (_23941_, _23434_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _28452_ (_23942_, _23197_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _28453_ (_23943_, _23942_, _23941_);
  or _28454_ (_23944_, _23943_, _23940_);
  or _28455_ (_23945_, _23944_, _23914_);
  and _28456_ (_23946_, _23945_, _22946_);
  and _28457_ (_23947_, _23946_, _23912_);
  not _28458_ (_23948_, _23912_);
  and _28459_ (_23949_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  or _28460_ (_22757_, _23949_, _23947_);
  not _28461_ (_23950_, _22768_);
  nor _28462_ (_23951_, _23848_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _28463_ (_23952_, _23951_, _23950_);
  nor _28464_ (_23953_, _23952_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _28465_ (_23954_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  not _28466_ (_23955_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor _28467_ (_23956_, _23953_, _23955_);
  or _28468_ (_23957_, _23956_, _23954_);
  and _28469_ (_26904_[31], _23957_, _22762_);
  and _28470_ (_23958_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _28471_ (_23959_, _23958_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  or _28472_ (_23960_, _23959_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _28473_ (_26902_[3], _23960_, _22762_);
  or _28474_ (_23961_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  nand _28475_ (_23962_, _23953_, _23955_);
  and _28476_ (_23963_, _23962_, _22762_);
  and _28477_ (_26903_[31], _23963_, _23961_);
  and _28478_ (_26900_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _22762_);
  not _28479_ (_23964_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _28480_ (_23965_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor _28481_ (_23966_, _23965_, _23964_);
  and _28482_ (_23967_, _23965_, _23964_);
  nor _28483_ (_23968_, _23967_, _23966_);
  not _28484_ (_23969_, _23968_);
  and _28485_ (_23970_, _23969_, _26902_[3]);
  nor _28486_ (_23971_, _23966_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _28487_ (_23972_, _23966_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _28488_ (_23973_, _23972_, _23971_);
  nor _28489_ (_23974_, _23958_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _28490_ (_23975_, _23974_, _23959_);
  or _28491_ (_23976_, _23975_, _23965_);
  and _28492_ (_23977_, _23976_, _23973_);
  and _28493_ (_26901_, _23977_, _23970_);
  not _28494_ (_23978_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and _28495_ (_23979_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _23978_);
  and _28496_ (_23980_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _28497_ (_23981_, _23980_, _23979_);
  and _28498_ (_26899_[7], _23981_, _22762_);
  and _28499_ (_23982_, _23907_, _23898_);
  and _28500_ (_23983_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or _28501_ (_24175_, _23983_, _23982_);
  and _28502_ (_23984_, _23755_, _23649_);
  and _28503_ (_23985_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  or _28504_ (_24247_, _23985_, _23984_);
  and _28505_ (_23986_, _23751_, _23068_);
  and _28506_ (_23987_, _23986_, _23906_);
  and _28507_ (_23988_, _23987_, _23747_);
  not _28508_ (_23989_, _23987_);
  and _28509_ (_23990_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  or _28510_ (_24383_, _23990_, _23988_);
  and _28511_ (_23991_, _23902_, _23021_);
  and _28512_ (_23992_, _23991_, _23906_);
  and _28513_ (_23993_, _23992_, _23778_);
  not _28514_ (_23994_, _23992_);
  and _28515_ (_23995_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or _28516_ (_26943_, _23995_, _23993_);
  and _28517_ (_23997_, _23946_, _23907_);
  and _28518_ (_23998_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or _28519_ (_26940_, _23998_, _23997_);
  and _28520_ (_24000_, _23907_, _23707_);
  and _28521_ (_24001_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or _28522_ (_26941_, _24001_, _24000_);
  and _28523_ (_24003_, _23907_, _23649_);
  and _28524_ (_24004_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or _28525_ (_26939_, _24004_, _24003_);
  and _28526_ (_24005_, _23902_, _23782_);
  and _28527_ (_24006_, _24005_, _23906_);
  and _28528_ (_24007_, _24006_, _23707_);
  not _28529_ (_24008_, _24006_);
  and _28530_ (_24009_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or _28531_ (_26938_, _24009_, _24007_);
  and _28532_ (_24010_, _23783_, _23021_);
  and _28533_ (_24011_, _24010_, _23789_);
  and _28534_ (_24012_, _24011_, _23707_);
  not _28535_ (_24013_, _24011_);
  and _28536_ (_24014_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or _28537_ (_27264_, _24014_, _24012_);
  nand _28538_ (_24015_, _23427_, _23079_);
  nor _28539_ (_24016_, _24015_, _23594_);
  nor _28540_ (_24017_, _23607_, _23171_);
  and _28541_ (_24018_, _23677_, _23171_);
  not _28542_ (_24019_, _24018_);
  and _28543_ (_24020_, _24019_, _23679_);
  and _28544_ (_24021_, _23673_, _23522_);
  nor _28545_ (_24022_, _24021_, _23171_);
  nor _28546_ (_24023_, _24022_, _23674_);
  nor _28547_ (_24024_, _24023_, _23521_);
  or _28548_ (_24025_, _24024_, _24020_);
  nand _28549_ (_24026_, _24025_, _23609_);
  and _28550_ (_24027_, _23456_, _23177_);
  not _28551_ (_24028_, _23171_);
  and _28552_ (_24029_, _23521_, _24028_);
  nor _28553_ (_24030_, _24029_, _24027_);
  nor _28554_ (_24031_, _24030_, _23688_);
  not _28555_ (_24032_, _24031_);
  and _28556_ (_24033_, _23550_, _23182_);
  nor _28557_ (_24034_, _23634_, _23181_);
  or _28558_ (_24035_, _24034_, _24033_);
  not _28559_ (_24036_, _24035_);
  and _28560_ (_24037_, _23583_, _23180_);
  and _28561_ (_24038_, _23557_, _23171_);
  nor _28562_ (_24039_, _24038_, _24037_);
  and _28563_ (_24040_, _24039_, _24036_);
  and _28564_ (_24041_, _24040_, _24032_);
  nand _28565_ (_24042_, _24041_, _24026_);
  or _28566_ (_24043_, _24042_, _24017_);
  and _28567_ (_24044_, _24043_, _22948_);
  nand _28568_ (_24045_, _23427_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _28569_ (_24046_, _23160_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _28570_ (_24047_, _24046_, _24045_);
  or _28571_ (_24048_, _24047_, _24044_);
  or _28572_ (_24049_, _24048_, _24016_);
  and _28573_ (_24050_, _24049_, _22946_);
  and _28574_ (_24051_, _24050_, _24011_);
  and _28575_ (_24052_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or _28576_ (_27263_, _24052_, _24051_);
  and _28577_ (_24053_, _23833_, _23649_);
  and _28578_ (_24054_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or _28579_ (_27064_, _24054_, _24053_);
  and _28580_ (_24055_, _23833_, _23747_);
  and _28581_ (_24056_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or _28582_ (_27063_, _24056_, _24055_);
  and _28583_ (_24057_, _23912_, _23747_);
  and _28584_ (_24058_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  or _28585_ (_27267_, _24058_, _24057_);
  and _28586_ (_24059_, _23912_, _23824_);
  and _28587_ (_24060_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  or _28588_ (_27266_, _24060_, _24059_);
  and _28589_ (_24061_, _23912_, _23898_);
  and _28590_ (_24062_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  or _28591_ (_27265_, _24062_, _24061_);
  and _28592_ (_24063_, _23052_, _22970_);
  and _28593_ (_24064_, _24063_, _23753_);
  not _28594_ (_24065_, _23018_);
  and _28595_ (_24066_, _23065_, _22983_);
  and _28596_ (_24067_, _24066_, _24065_);
  nor _28597_ (_24068_, _22909_, _22906_);
  and _28598_ (_24069_, _24068_, _22948_);
  not _28599_ (_24070_, _24069_);
  nor _28600_ (_24071_, _24070_, _23002_);
  and _28601_ (_24072_, _24071_, _24067_);
  and _28602_ (_24073_, _24072_, _24064_);
  or _28603_ (_24074_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _28604_ (_24075_, _24074_, _22762_);
  and _28605_ (_24076_, _24067_, _23003_);
  and _28606_ (_24077_, _24064_, _24069_);
  and _28607_ (_24078_, _24077_, _24076_);
  not _28608_ (_24079_, _24078_);
  or _28609_ (_24080_, _24079_, _23738_);
  and _28610_ (_26382_, _24080_, _24075_);
  and _28611_ (_24081_, _24010_, _23754_);
  and _28612_ (_24082_, _24081_, _23824_);
  not _28613_ (_24083_, _24081_);
  and _28614_ (_24084_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or _28615_ (_27052_, _24084_, _24082_);
  and _28616_ (_24085_, _23901_, _23783_);
  and _28617_ (_24086_, _24085_, _23789_);
  and _28618_ (_24087_, _24086_, _23707_);
  not _28619_ (_24088_, _24086_);
  and _28620_ (_24089_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or _28621_ (_27257_, _24089_, _24087_);
  and _28622_ (_24090_, _24011_, _23898_);
  and _28623_ (_24092_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or _28624_ (_27259_, _24092_, _24090_);
  and _28625_ (_24093_, _24081_, _23898_);
  and _28626_ (_24094_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or _28627_ (_27051_, _24094_, _24093_);
  nor _28628_ (_24095_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _28629_ (_24096_, _24095_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _28630_ (_26907_, _24096_, _22762_);
  and _28631_ (_24098_, _26900_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _28632_ (_26906_, _24098_, _26907_);
  and _28633_ (_24100_, _24011_, _23778_);
  and _28634_ (_24101_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or _28635_ (_27258_, _24101_, _24100_);
  and _28636_ (_24102_, _24081_, _23778_);
  and _28637_ (_24103_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or _28638_ (_27050_, _24103_, _24102_);
  not _28639_ (_24104_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _28640_ (_24105_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , _24104_);
  and _28641_ (_26905_, _24105_, _22762_);
  and _28642_ (_24107_, _24011_, _23649_);
  and _28643_ (_24108_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or _28644_ (_27262_, _24108_, _24107_);
  and _28645_ (_24109_, _24011_, _23747_);
  and _28646_ (_24110_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or _28647_ (_27261_, _24110_, _24109_);
  and _28648_ (_24111_, _24011_, _23824_);
  and _28649_ (_24112_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or _28650_ (_27260_, _24112_, _24111_);
  and _28651_ (_24113_, _24081_, _23946_);
  and _28652_ (_24114_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or _28653_ (_27055_, _24114_, _24113_);
  and _28654_ (_24115_, _24081_, _23649_);
  and _28655_ (_24116_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or _28656_ (_27054_, _24116_, _24115_);
  nor _28657_ (_24117_, _23018_, _22983_);
  and _28658_ (_24118_, _24117_, _23065_);
  and _28659_ (_24119_, _24118_, _24071_);
  and _28660_ (_24120_, _24119_, _24064_);
  and _28661_ (_24121_, _24120_, _22762_);
  and _28662_ (_24122_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not _28663_ (_24123_, _23065_);
  and _28664_ (_24124_, _24065_, _22983_);
  and _28665_ (_24125_, _24124_, _24123_);
  and _28666_ (_24126_, _24125_, _24071_);
  and _28667_ (_24127_, _24126_, _24064_);
  not _28668_ (_24128_, _24127_);
  or _28669_ (_24129_, _24128_, _23892_);
  not _28670_ (_24130_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not _28671_ (_24131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _28672_ (_24132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _24131_);
  not _28673_ (_24134_, _24132_);
  not _28674_ (_24135_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not _28675_ (_24136_, t1_i);
  and _28676_ (_24137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _24136_);
  nor _28677_ (_24138_, _24137_, _24135_);
  not _28678_ (_24139_, _24138_);
  not _28679_ (_24140_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _28680_ (_24141_, _24140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  nor _28681_ (_24142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _28682_ (_24143_, _24142_);
  and _28683_ (_24144_, _24143_, _24141_);
  and _28684_ (_24145_, _24144_, _24139_);
  not _28685_ (_24146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand _28686_ (_24147_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand _28687_ (_24148_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _28688_ (_24149_, _24148_, _24147_);
  nor _28689_ (_24150_, _24149_, _24146_);
  and _28690_ (_24151_, _24150_, _24145_);
  and _28691_ (_24152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _28692_ (_24153_, _24152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _28693_ (_24154_, _24153_, _24151_);
  nor _28694_ (_24155_, _24154_, _24134_);
  not _28695_ (_24156_, _24155_);
  not _28696_ (_24157_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _28697_ (_24158_, _24151_, _24131_);
  nor _28698_ (_24159_, _24158_, _24132_);
  nor _28699_ (_24160_, _24159_, _24157_);
  and _28700_ (_24161_, _24160_, _24156_);
  nor _28701_ (_24162_, _24161_, _24130_);
  and _28702_ (_24163_, _24161_, _24130_);
  or _28703_ (_24164_, _24163_, _24162_);
  or _28704_ (_24165_, _24164_, _24127_);
  nor _28705_ (_24166_, _24120_, rst);
  and _28706_ (_24167_, _24166_, _24165_);
  and _28707_ (_24168_, _24167_, _24129_);
  or _28708_ (_00740_, _24168_, _24122_);
  and _28709_ (_24169_, _24081_, _23747_);
  and _28710_ (_24170_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or _28711_ (_27053_, _24170_, _24169_);
  not _28712_ (_24171_, _24120_);
  or _28713_ (_24172_, _24171_, _23642_);
  and _28714_ (_24173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _28715_ (_24174_, _24173_, _24127_);
  nor _28716_ (_24176_, _24174_, _24146_);
  not _28717_ (_24177_, _24145_);
  nor _28718_ (_24178_, _24149_, _24177_);
  or _28719_ (_24179_, _24178_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _28720_ (_24180_, _24173_, _24151_);
  and _28721_ (_24181_, _24180_, _24179_);
  not _28722_ (_24182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _28723_ (_24184_, _24182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _28724_ (_24185_, _24184_, _24154_);
  and _28725_ (_24186_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _28726_ (_24187_, _24186_, _24181_);
  nor _28727_ (_24188_, _24187_, _24127_);
  or _28728_ (_24189_, _24188_, _24176_);
  or _28729_ (_24190_, _24189_, _24120_);
  and _28730_ (_24191_, _24190_, _22762_);
  and _28731_ (_00832_, _24191_, _24172_);
  and _28732_ (_24192_, _24086_, _23946_);
  and _28733_ (_24193_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or _28734_ (_27255_, _24193_, _24192_);
  and _28735_ (_24194_, _24085_, _23754_);
  and _28736_ (_24195_, _24194_, _23747_);
  not _28737_ (_24196_, _24194_);
  and _28738_ (_24197_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or _28739_ (_27048_, _24197_, _24195_);
  and _28740_ (_24198_, _24194_, _23649_);
  and _28741_ (_24199_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or _28742_ (_27049_, _24199_, _24198_);
  and _28743_ (_24201_, _23788_, _23661_);
  and _28744_ (_24203_, _24201_, _23991_);
  not _28745_ (_24204_, _24203_);
  and _28746_ (_24206_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  and _28747_ (_24207_, _24203_, _23747_);
  or _28748_ (_27248_, _24207_, _24206_);
  and _28749_ (_01412_, t1_i, _22762_);
  and _28750_ (_24208_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  and _28751_ (_24209_, _24203_, _23824_);
  or _28752_ (_27247_, _24209_, _24208_);
  and _28753_ (_24210_, _23824_, _23077_);
  and _28754_ (_24211_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  or _28755_ (_27214_, _24211_, _24210_);
  and _28756_ (_24212_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  and _28757_ (_24213_, _24203_, _23707_);
  or _28758_ (_01716_, _24213_, _24212_);
  and _28759_ (_24214_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  and _28760_ (_24215_, _24203_, _24050_);
  or _28761_ (_27250_, _24215_, _24214_);
  and _28762_ (_24216_, _24194_, _23707_);
  and _28763_ (_24217_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or _28764_ (_01953_, _24217_, _24216_);
  and _28765_ (_24218_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  and _28766_ (_24219_, _24203_, _23946_);
  or _28767_ (_27249_, _24219_, _24218_);
  and _28768_ (_24220_, _24194_, _24050_);
  and _28769_ (_24221_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or _28770_ (_02060_, _24221_, _24220_);
  and _28771_ (_24222_, _24201_, _23903_);
  not _28772_ (_24223_, _24222_);
  and _28773_ (_24224_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  and _28774_ (_24225_, _24222_, _23946_);
  or _28775_ (_02437_, _24225_, _24224_);
  and _28776_ (_24226_, _23784_, _23754_);
  and _28777_ (_24228_, _24226_, _23707_);
  not _28778_ (_24229_, _24226_);
  and _28779_ (_24230_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  or _28780_ (_02582_, _24230_, _24228_);
  and _28781_ (_24231_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _28782_ (_24232_, _24127_, _23702_);
  and _28783_ (_24234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _28784_ (_24235_, _24234_, _24150_);
  and _28785_ (_24236_, _24235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _28786_ (_24237_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _28787_ (_24238_, _24237_, _24236_);
  and _28788_ (_24239_, _24238_, _24153_);
  and _28789_ (_24240_, _24145_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _28790_ (_24241_, _24240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _28791_ (_24242_, _24241_, _24239_);
  and _28792_ (_24243_, _24242_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _28793_ (_24244_, _24242_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _28794_ (_24245_, _24244_, _24132_);
  nor _28795_ (_24246_, _24245_, _24243_);
  and _28796_ (_24248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _28797_ (_24249_, _24236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _28798_ (_24250_, _24249_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _28799_ (_24251_, _24250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _28800_ (_24252_, _24251_, _24145_);
  and _28801_ (_24253_, _24252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _28802_ (_24254_, _24253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _28803_ (_24255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _28804_ (_24256_, _24255_);
  and _28805_ (_24257_, _24253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _28806_ (_24258_, _24257_, _24256_);
  and _28807_ (_24259_, _24258_, _24254_);
  or _28808_ (_24260_, _24259_, _24248_);
  or _28809_ (_24261_, _24260_, _24246_);
  or _28810_ (_24262_, _24261_, _24127_);
  and _28811_ (_24263_, _24262_, _24166_);
  and _28812_ (_24264_, _24263_, _24232_);
  or _28813_ (_02663_, _24264_, _24231_);
  and _28814_ (_24265_, _24226_, _24050_);
  and _28815_ (_24266_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  or _28816_ (_02867_, _24266_, _24265_);
  and _28817_ (_24267_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  and _28818_ (_24268_, _24203_, _23778_);
  or _28819_ (_02903_, _24268_, _24267_);
  and _28820_ (_24269_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  and _28821_ (_24270_, _24222_, _23707_);
  or _28822_ (_03083_, _24270_, _24269_);
  and _28823_ (_24271_, _24194_, _23778_);
  and _28824_ (_24272_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or _28825_ (_03542_, _24272_, _24271_);
  and _28826_ (_24273_, _24194_, _23898_);
  and _28827_ (_24274_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or _28828_ (_27046_, _24274_, _24273_);
  and _28829_ (_24275_, _23902_, _23751_);
  and _28830_ (_24276_, _24275_, _24201_);
  not _28831_ (_24277_, _24276_);
  and _28832_ (_24279_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  and _28833_ (_24280_, _24276_, _23824_);
  or _28834_ (_03788_, _24280_, _24279_);
  and _28835_ (_24282_, _23782_, _23655_);
  and _28836_ (_24283_, _24282_, _23076_);
  and _28837_ (_24284_, _24283_, _23824_);
  not _28838_ (_24285_, _24283_);
  and _28839_ (_24286_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  or _28840_ (_03822_, _24286_, _24284_);
  and _28841_ (_24287_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  and _28842_ (_24288_, _24276_, _23898_);
  or _28843_ (_03855_, _24288_, _24287_);
  not _28844_ (_24289_, _22983_);
  and _28845_ (_24290_, _23018_, _24289_);
  and _28846_ (_24291_, _24290_, _23065_);
  and _28847_ (_24292_, _24291_, _24071_);
  and _28848_ (_24293_, _24292_, _24064_);
  not _28849_ (_24294_, _24293_);
  and _28850_ (_24295_, _23018_, _22983_);
  and _28851_ (_24296_, _24295_, _24123_);
  and _28852_ (_24297_, _24296_, _24071_);
  and _28853_ (_24299_, _24297_, _24064_);
  and _28854_ (_24300_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  or _28855_ (_24301_, _24300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and _28856_ (_24302_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _28857_ (_24303_, _24302_, _22762_);
  and _28858_ (_24304_, _24303_, _24301_);
  not _28859_ (_24305_, _24300_);
  and _28860_ (_24307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _28861_ (_24308_, _24307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _28862_ (_24309_, _24308_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _28863_ (_24310_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _28864_ (_24312_, _24310_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _28865_ (_24313_, _24312_, _24309_);
  and _28866_ (_24315_, _24313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _28867_ (_24316_, _24315_, _24305_);
  nand _28868_ (_24317_, _24316_, _24304_);
  nor _28869_ (_24318_, _24317_, _24299_);
  and _28870_ (_04338_, _24318_, _24294_);
  and _28871_ (_24319_, _24226_, _23778_);
  and _28872_ (_24320_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  or _28873_ (_04361_, _24320_, _24319_);
  and _28874_ (_24322_, _24226_, _23898_);
  and _28875_ (_24323_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  or _28876_ (_04416_, _24323_, _24322_);
  and _28877_ (_24324_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and _28878_ (_24325_, _24276_, _23946_);
  or _28879_ (_04519_, _24325_, _24324_);
  and _28880_ (_24326_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and _28881_ (_24328_, _24276_, _23649_);
  or _28882_ (_04742_, _24328_, _24326_);
  and _28883_ (_24329_, _23782_, _23068_);
  and _28884_ (_24331_, _24329_, _23754_);
  and _28885_ (_24332_, _24331_, _23778_);
  not _28886_ (_24333_, _24331_);
  and _28887_ (_24334_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or _28888_ (_04802_, _24334_, _24332_);
  and _28889_ (_24335_, _23898_, _23077_);
  and _28890_ (_24336_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  or _28891_ (_04851_, _24336_, _24335_);
  and _28892_ (_24337_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  not _28893_ (_24338_, _24337_);
  nand _28894_ (_24339_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _28895_ (_24340_, _24339_, _24338_);
  nand _28896_ (_24341_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand _28897_ (_24342_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _28898_ (_24343_, _24342_, _24341_);
  nand _28899_ (_24344_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand _28900_ (_24345_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and _28901_ (_24346_, _24345_, _24344_);
  and _28902_ (_24347_, _24346_, _24343_);
  and _28903_ (_24348_, _24347_, _24340_);
  or _28904_ (_24349_, _24348_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _28905_ (_24350_, _24349_, _23838_);
  nor _28906_ (_24351_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _23838_);
  or _28907_ (_24352_, _24351_, _24350_);
  nor _28908_ (_26860_[3], _24352_, rst);
  and _28909_ (_24353_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and _28910_ (_24354_, _24276_, _23707_);
  or _28911_ (_05258_, _24354_, _24353_);
  and _28912_ (_24356_, _23785_, _23075_);
  and _28913_ (_24358_, _24356_, _24282_);
  and _28914_ (_24359_, _24358_, _23824_);
  not _28915_ (_24360_, _24358_);
  and _28916_ (_24361_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  or _28917_ (_05587_, _24361_, _24359_);
  and _28918_ (_24362_, _24226_, _23747_);
  and _28919_ (_24363_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  or _28920_ (_27045_, _24363_, _24362_);
  and _28921_ (_24364_, _24358_, _23898_);
  and _28922_ (_24365_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  or _28923_ (_05673_, _24365_, _24364_);
  and _28924_ (_24366_, _24226_, _23649_);
  and _28925_ (_24367_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  or _28926_ (_05825_, _24367_, _24366_);
  and _28927_ (_24368_, _24358_, _23778_);
  and _28928_ (_24369_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  or _28929_ (_05902_, _24369_, _24368_);
  and _28930_ (_24370_, _23905_, _23075_);
  and _28931_ (_24371_, _24370_, _23991_);
  and _28932_ (_24372_, _24371_, _23707_);
  not _28933_ (_24373_, _24371_);
  and _28934_ (_24374_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or _28935_ (_06170_, _24374_, _24372_);
  and _28936_ (_24375_, _24370_, _23784_);
  and _28937_ (_24376_, _24375_, _23778_);
  not _28938_ (_24377_, _24375_);
  and _28939_ (_24378_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or _28940_ (_06542_, _24378_, _24376_);
  and _28941_ (_24379_, _24375_, _23824_);
  and _28942_ (_24380_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or _28943_ (_06585_, _24380_, _24379_);
  and _28944_ (_24381_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _28945_ (_24382_, _22767_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _28946_ (_24384_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _28947_ (_24385_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and _28948_ (_24386_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _28949_ (_24388_, _24386_, _24385_);
  and _28950_ (_24389_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _28951_ (_24391_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _28952_ (_24392_, _24391_, _24389_);
  and _28953_ (_24393_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and _28954_ (_24394_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _28955_ (_24396_, _24394_, _24393_);
  and _28956_ (_24397_, _24396_, _24392_);
  and _28957_ (_24399_, _24397_, _24388_);
  nor _28958_ (_24400_, _24399_, _24384_);
  and _28959_ (_24401_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  nor _28960_ (_24402_, _24401_, _24400_);
  and _28961_ (_24403_, _24402_, _22769_);
  not _28962_ (_24404_, _24403_);
  not _28963_ (_24405_, _22765_);
  nor _28964_ (_24406_, _22768_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _28965_ (_24407_, _24406_, _24405_);
  and _28966_ (_24408_, _24407_, _24404_);
  not _28967_ (_24409_, _22769_);
  nor _28968_ (_24411_, _23866_, _24409_);
  not _28969_ (_24412_, _24411_);
  nor _28970_ (_24414_, _22768_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _28971_ (_24415_, _24414_, _24405_);
  and _28972_ (_24417_, _24415_, _24412_);
  and _28973_ (_24418_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _28974_ (_24420_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _28975_ (_24421_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or _28976_ (_24422_, _24421_, _24420_);
  and _28977_ (_24424_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _28978_ (_24425_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and _28979_ (_24426_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _28980_ (_24427_, _24426_, _24425_);
  or _28981_ (_24428_, _24427_, _24424_);
  or _28982_ (_24429_, _24428_, _24422_);
  or _28983_ (_24430_, _24429_, _24418_);
  nand _28984_ (_24431_, _24430_, _23839_);
  nand _28985_ (_24432_, _24431_, _23838_);
  nor _28986_ (_24434_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _23838_);
  not _28987_ (_24435_, _24434_);
  and _28988_ (_24436_, _24435_, _24432_);
  or _28989_ (_24437_, _24436_, _24409_);
  nor _28990_ (_24438_, _22768_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _28991_ (_24439_, _24438_, _24405_);
  and _28992_ (_24440_, _24439_, _24437_);
  and _28993_ (_24441_, _24352_, _22769_);
  not _28994_ (_24442_, _24441_);
  nor _28995_ (_24443_, _22768_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _28996_ (_24444_, _24443_, _24405_);
  and _28997_ (_24445_, _24444_, _24442_);
  nor _28998_ (_24446_, _24445_, _24440_);
  and _28999_ (_24447_, _24446_, _24417_);
  and _29000_ (_24448_, _24447_, _24408_);
  and _29001_ (_24450_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _29002_ (_24451_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and _29003_ (_24452_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _29004_ (_24453_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _29005_ (_24454_, _24453_, _24452_);
  and _29006_ (_24455_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and _29007_ (_24456_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _29008_ (_24457_, _24456_, _24455_);
  nand _29009_ (_24458_, _24457_, _24454_);
  or _29010_ (_24459_, _24458_, _24451_);
  nor _29011_ (_24460_, _24459_, _24450_);
  and _29012_ (_24461_, _24460_, _23839_);
  and _29013_ (_24462_, _24461_, _23838_);
  nor _29014_ (_24463_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _23838_);
  nor _29015_ (_24464_, _24463_, _24462_);
  nor _29016_ (_24466_, _24464_, _24409_);
  not _29017_ (_24467_, _24466_);
  nor _29018_ (_24469_, _22768_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _29019_ (_24470_, _24469_, _24405_);
  nand _29020_ (_24471_, _24470_, _24467_);
  nand _29021_ (_24472_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand _29022_ (_24473_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _29023_ (_24474_, _24473_, _24472_);
  nand _29024_ (_24475_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nand _29025_ (_24476_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and _29026_ (_24477_, _24476_, _24475_);
  and _29027_ (_24478_, _24477_, _24474_);
  and _29028_ (_24479_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _29029_ (_24480_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor _29030_ (_24481_, _24480_, _24479_);
  and _29031_ (_24482_, _24481_, _24478_);
  or _29032_ (_24483_, _24482_, _24384_);
  and _29033_ (_24484_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _29034_ (_24485_, _24484_);
  and _29035_ (_24486_, _24485_, _24483_);
  nand _29036_ (_24487_, _24486_, _22769_);
  nor _29037_ (_24488_, _22768_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _29038_ (_24489_, _24488_, _24405_);
  and _29039_ (_24490_, _24489_, _24487_);
  and _29040_ (_24491_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _29041_ (_24492_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _29042_ (_24493_, _24492_, _24491_);
  nand _29043_ (_24494_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nand _29044_ (_24495_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and _29045_ (_24497_, _24495_, _24494_);
  nand _29046_ (_24498_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand _29047_ (_24500_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _29048_ (_24501_, _24500_, _24498_);
  and _29049_ (_24503_, _24501_, _24497_);
  and _29050_ (_24504_, _24503_, _24493_);
  or _29051_ (_24505_, _24504_, _24384_);
  and _29052_ (_24506_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _29053_ (_24507_, _24506_);
  and _29054_ (_24508_, _24507_, _24505_);
  nand _29055_ (_24509_, _24508_, _22769_);
  nor _29056_ (_24510_, _22768_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _29057_ (_24511_, _24510_, _24405_);
  and _29058_ (_24512_, _24511_, _24509_);
  not _29059_ (_24513_, _24512_);
  nor _29060_ (_24514_, _24513_, _24490_);
  nor _29061_ (_24515_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _29062_ (_24516_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _29063_ (_24517_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _29064_ (_24518_, _24517_, _24516_);
  and _29065_ (_24519_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and _29066_ (_24520_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _29067_ (_24521_, _24520_, _24519_);
  and _29068_ (_24522_, _24521_, _24518_);
  and _29069_ (_24523_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _29070_ (_24524_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor _29071_ (_24525_, _24524_, _24523_);
  nand _29072_ (_24526_, _24525_, _24522_);
  nand _29073_ (_24527_, _24526_, _24515_);
  and _29074_ (_24528_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _29075_ (_24529_, _24528_);
  and _29076_ (_24530_, _24529_, _24527_);
  nand _29077_ (_24531_, _24530_, _22769_);
  nor _29078_ (_24532_, _22768_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _29079_ (_24533_, _24532_, _24405_);
  and _29080_ (_24534_, _24533_, _24531_);
  and _29081_ (_24535_, _24534_, _24514_);
  and _29082_ (_24536_, _24535_, _24471_);
  and _29083_ (_24537_, _24536_, _24448_);
  and _29084_ (_24538_, _24470_, _24467_);
  and _29085_ (_24539_, _24513_, _24490_);
  and _29086_ (_24540_, _24539_, _24534_);
  and _29087_ (_24541_, _24540_, _24538_);
  and _29088_ (_24542_, _24541_, _24448_);
  nor _29089_ (_24543_, _24542_, _24537_);
  not _29090_ (_24544_, _24534_);
  and _29091_ (_24545_, _24544_, _24514_);
  and _29092_ (_24546_, _24545_, _24538_);
  and _29093_ (_24548_, _24546_, _24448_);
  not _29094_ (_24549_, _24548_);
  and _29095_ (_24550_, _24549_, _24543_);
  and _29096_ (_24552_, _24545_, _24471_);
  not _29097_ (_24553_, _24445_);
  and _29098_ (_24554_, _24553_, _24440_);
  nor _29099_ (_24555_, _24417_, _24408_);
  and _29100_ (_24556_, _24555_, _24554_);
  and _29101_ (_24558_, _24556_, _24552_);
  and _29102_ (_24559_, _24556_, _24536_);
  nor _29103_ (_24560_, _24559_, _24558_);
  and _29104_ (_24561_, _24560_, _24550_);
  nor _29105_ (_24562_, _24561_, _24382_);
  not _29106_ (_24563_, _24562_);
  not _29107_ (_24564_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _29108_ (_24565_, \oc8051_top_1.oc8051_decoder1.state [1], _22766_);
  and _29109_ (_24566_, _24565_, _24564_);
  and _29110_ (_24567_, _24555_, _24446_);
  and _29111_ (_24568_, _24567_, _24539_);
  and _29112_ (_24569_, _24568_, _24566_);
  nor _29113_ (_24570_, _24560_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _29114_ (_24572_, _24570_, _23837_);
  nor _29115_ (_24573_, _24572_, _24569_);
  and _29116_ (_24574_, _24573_, _24563_);
  nor _29117_ (_24575_, _24574_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _29118_ (_24576_, _24575_, _24381_);
  not _29119_ (_24577_, _24576_);
  and _29120_ (_24578_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _29121_ (_24579_, _24578_);
  and _29122_ (_24581_, _24554_, _24417_);
  and _29123_ (_24582_, _24544_, _24490_);
  and _29124_ (_24584_, _24582_, _24512_);
  and _29125_ (_24585_, _24584_, _24581_);
  and _29126_ (_24586_, _24581_, _24546_);
  or _29127_ (_24587_, _24586_, _24585_);
  and _29128_ (_24588_, _24539_, _24544_);
  and _29129_ (_24589_, _24588_, _24538_);
  and _29130_ (_24591_, _24581_, _24589_);
  nor _29131_ (_24592_, _24512_, _24490_);
  and _29132_ (_24593_, _24592_, _24534_);
  and _29133_ (_24594_, _24593_, _24581_);
  or _29134_ (_24595_, _24594_, _24591_);
  and _29135_ (_24596_, _24581_, _24471_);
  and _29136_ (_24597_, _24534_, _24490_);
  and _29137_ (_24598_, _24597_, _24512_);
  or _29138_ (_24599_, _24598_, _24588_);
  and _29139_ (_24600_, _24599_, _24596_);
  or _29140_ (_24601_, _24600_, _24595_);
  nor _29141_ (_24602_, _24601_, _24587_);
  and _29142_ (_24604_, _24540_, _24471_);
  and _29143_ (_24605_, _24581_, _24604_);
  and _29144_ (_24606_, _24535_, _24538_);
  and _29145_ (_24607_, _24606_, _24581_);
  and _29146_ (_24608_, _24581_, _24552_);
  or _29147_ (_24610_, _24608_, _24607_);
  nor _29148_ (_24611_, _24610_, _24605_);
  not _29149_ (_24612_, _24408_);
  and _29150_ (_24613_, _24447_, _24612_);
  and _29151_ (_24614_, _24613_, _24593_);
  not _29152_ (_24615_, _24614_);
  and _29153_ (_24616_, _24592_, _24544_);
  and _29154_ (_24617_, _24616_, _24581_);
  and _29155_ (_24618_, _24584_, _24538_);
  and _29156_ (_24619_, _24618_, _24567_);
  nor _29157_ (_24620_, _24619_, _24617_);
  and _29158_ (_24621_, _24620_, _24615_);
  and _29159_ (_24622_, _24621_, _24611_);
  and _29160_ (_24623_, _24622_, _24602_);
  and _29161_ (_24624_, _24623_, _24550_);
  nor _29162_ (_24625_, _24624_, _24382_);
  and _29163_ (_24626_, \oc8051_top_1.oc8051_decoder1.state [0], _22766_);
  and _29164_ (_24627_, _24626_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _29165_ (_24628_, _24614_, _24627_);
  and _29166_ (_24629_, _24566_, _24540_);
  and _29167_ (_24630_, _24629_, _24567_);
  or _29168_ (_24631_, _24630_, _24628_);
  or _29169_ (_24632_, _24631_, _24625_);
  nand _29170_ (_24633_, _24632_, _22766_);
  and _29171_ (_24634_, _24633_, _24579_);
  nor _29172_ (_24635_, _24634_, _24577_);
  and _29173_ (_26909_, _24635_, _22762_);
  and _29174_ (_24636_, _24375_, _23747_);
  and _29175_ (_24637_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or _29176_ (_27175_, _24637_, _24636_);
  and _29177_ (_24639_, _24356_, _24005_);
  and _29178_ (_24640_, _24639_, _24050_);
  not _29179_ (_24641_, _24639_);
  and _29180_ (_24642_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or _29181_ (_27170_, _24642_, _24640_);
  and _29182_ (_24643_, _23053_, _23034_);
  nor _29183_ (_24644_, _23002_, _22970_);
  and _29184_ (_24645_, _24068_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _29185_ (_24646_, _24645_, _22943_);
  and _29186_ (_24647_, _24646_, _24644_);
  and _29187_ (_24648_, _24647_, _24643_);
  and _29188_ (_24649_, _24648_, _24118_);
  nand _29189_ (_24650_, _24649_, _23594_);
  or _29190_ (_24651_, _24649_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _29191_ (_24652_, _24069_, _23002_);
  nor _29192_ (_24653_, _23065_, _22983_);
  and _29193_ (_24654_, _24653_, _24065_);
  and _29194_ (_24655_, _24654_, _24652_);
  nor _29195_ (_24656_, _23052_, _22970_);
  and _29196_ (_24657_, _24656_, _23753_);
  and _29197_ (_24658_, _24657_, _24655_);
  not _29198_ (_24659_, _24658_);
  and _29199_ (_24660_, _24659_, _24651_);
  and _29200_ (_24661_, _24660_, _24650_);
  and _29201_ (_24662_, _24658_, _23738_);
  or _29202_ (_24663_, _24662_, _24661_);
  and _29203_ (_06844_, _24663_, _22762_);
  and _29204_ (_24664_, _24648_, _24291_);
  nand _29205_ (_24665_, _24664_, _23594_);
  or _29206_ (_24666_, _24664_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _29207_ (_24667_, _24666_, _24659_);
  and _29208_ (_24668_, _24667_, _24665_);
  and _29209_ (_24669_, _24658_, _23816_);
  or _29210_ (_24670_, _24669_, _24668_);
  and _29211_ (_06893_, _24670_, _22762_);
  and _29212_ (_24671_, _24648_, _24067_);
  nand _29213_ (_24672_, _24671_, _23594_);
  or _29214_ (_24673_, _24671_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _29215_ (_24674_, _24673_, _24659_);
  and _29216_ (_24675_, _24674_, _24672_);
  and _29217_ (_24676_, _24658_, _23892_);
  or _29218_ (_24677_, _24676_, _24675_);
  and _29219_ (_06909_, _24677_, _22762_);
  and _29220_ (_24678_, _24066_, _23018_);
  and _29221_ (_24679_, _24678_, _24648_);
  nand _29222_ (_24680_, _24679_, _23594_);
  or _29223_ (_24682_, _24679_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _29224_ (_24683_, _24682_, _24659_);
  and _29225_ (_24684_, _24683_, _24680_);
  not _29226_ (_24685_, _23772_);
  and _29227_ (_24686_, _24658_, _24685_);
  or _29228_ (_24687_, _24686_, _24684_);
  and _29229_ (_06934_, _24687_, _22762_);
  and _29230_ (_24688_, _24356_, _23903_);
  and _29231_ (_24689_, _24688_, _23898_);
  not _29232_ (_24690_, _24688_);
  and _29233_ (_24691_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  or _29234_ (_06977_, _24691_, _24689_);
  and _29235_ (_24692_, _24201_, _23656_);
  not _29236_ (_24693_, _24692_);
  and _29237_ (_24694_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  and _29238_ (_24695_, _24692_, _23898_);
  or _29239_ (_07011_, _24695_, _24694_);
  and _29240_ (_24696_, _24688_, _23747_);
  and _29241_ (_24698_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  or _29242_ (_07034_, _24698_, _24696_);
  and _29243_ (_24699_, _24370_, _24329_);
  and _29244_ (_24700_, _24699_, _23824_);
  not _29245_ (_24701_, _24699_);
  and _29246_ (_24702_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  or _29247_ (_07185_, _24702_, _24700_);
  and _29248_ (_24703_, _24688_, _23946_);
  and _29249_ (_24704_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  or _29250_ (_07208_, _24704_, _24703_);
  and _29251_ (_24705_, _24653_, _23018_);
  and _29252_ (_24706_, _24705_, _24648_);
  nand _29253_ (_24707_, _24706_, _23594_);
  or _29254_ (_24708_, _24706_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _29255_ (_24709_, _24708_, _24659_);
  and _29256_ (_24710_, _24709_, _24707_);
  and _29257_ (_24711_, _24658_, _24043_);
  or _29258_ (_24712_, _24711_, _24710_);
  and _29259_ (_07234_, _24712_, _22762_);
  and _29260_ (_24713_, _24688_, _23707_);
  and _29261_ (_24714_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  or _29262_ (_27171_, _24714_, _24713_);
  and _29263_ (_24715_, _24648_, _24125_);
  nand _29264_ (_24716_, _24715_, _23594_);
  or _29265_ (_24717_, _24715_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _29266_ (_24718_, _24717_, _24659_);
  and _29267_ (_24719_, _24718_, _24716_);
  and _29268_ (_24720_, _24658_, _23939_);
  or _29269_ (_24721_, _24720_, _24719_);
  and _29270_ (_07281_, _24721_, _22762_);
  and _29271_ (_24722_, _24356_, _23991_);
  and _29272_ (_24723_, _24722_, _23778_);
  not _29273_ (_24724_, _24722_);
  and _29274_ (_24725_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  or _29275_ (_27173_, _24725_, _24723_);
  and _29276_ (_24726_, _24722_, _23898_);
  and _29277_ (_24727_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  or _29278_ (_07490_, _24727_, _24726_);
  and _29279_ (_24728_, _23003_, _22970_);
  and _29280_ (_24729_, _24728_, _24646_);
  and _29281_ (_24730_, _24729_, _24643_);
  and _29282_ (_24731_, _24730_, _24067_);
  nand _29283_ (_24732_, _24731_, _23594_);
  and _29284_ (_24733_, _23053_, _22970_);
  and _29285_ (_24734_, _24733_, _23753_);
  and _29286_ (_24735_, _24678_, _24071_);
  and _29287_ (_24736_, _24735_, _24734_);
  not _29288_ (_24737_, _24736_);
  or _29289_ (_24738_, _24731_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _29290_ (_24739_, _24738_, _24737_);
  and _29291_ (_24740_, _24739_, _24732_);
  and _29292_ (_24741_, _24736_, _23892_);
  or _29293_ (_24742_, _24741_, _24740_);
  and _29294_ (_07512_, _24742_, _22762_);
  and _29295_ (_24743_, _24722_, _23649_);
  and _29296_ (_24744_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  or _29297_ (_07528_, _24744_, _24743_);
  and _29298_ (_24745_, _24296_, _23711_);
  nor _29299_ (_24746_, _24295_, _24123_);
  and _29300_ (_24747_, _24746_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _29301_ (_24748_, _24747_, _24745_);
  and _29302_ (_24749_, _24748_, _24730_);
  not _29303_ (_24750_, _24730_);
  nor _29304_ (_24751_, _24295_, _23065_);
  or _29305_ (_24752_, _24751_, _24678_);
  or _29306_ (_24753_, _24752_, _24750_);
  and _29307_ (_24754_, _24753_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _29308_ (_24755_, _24754_, _24736_);
  or _29309_ (_24756_, _24755_, _24749_);
  or _29310_ (_24757_, _24737_, _23642_);
  and _29311_ (_24758_, _24757_, _22762_);
  and _29312_ (_07548_, _24758_, _24756_);
  and _29313_ (_24759_, _24730_, _24118_);
  nand _29314_ (_24760_, _24759_, _23594_);
  or _29315_ (_24761_, _24759_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _29316_ (_24762_, _24761_, _24737_);
  and _29317_ (_24763_, _24762_, _24760_);
  and _29318_ (_24764_, _24736_, _23738_);
  or _29319_ (_24765_, _24764_, _24763_);
  and _29320_ (_07595_, _24765_, _22762_);
  and _29321_ (_24766_, _23905_, _23753_);
  and _29322_ (_24767_, _24766_, _24275_);
  not _29323_ (_24768_, _24767_);
  and _29324_ (_24769_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and _29325_ (_24770_, _24767_, _23747_);
  or _29326_ (_07629_, _24770_, _24769_);
  and _29327_ (_24771_, _24730_, _24291_);
  nand _29328_ (_24772_, _24771_, _23594_);
  or _29329_ (_24773_, _24771_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _29330_ (_24774_, _24773_, _24737_);
  and _29331_ (_24775_, _24774_, _24772_);
  and _29332_ (_24776_, _24736_, _23816_);
  or _29333_ (_24777_, _24776_, _24775_);
  and _29334_ (_07661_, _24777_, _22762_);
  and _29335_ (_24778_, _24730_, _24678_);
  nand _29336_ (_24779_, _24778_, _23594_);
  or _29337_ (_24780_, _24778_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _29338_ (_24781_, _24780_, _24737_);
  and _29339_ (_24782_, _24781_, _24779_);
  and _29340_ (_24783_, _24736_, _24685_);
  or _29341_ (_24784_, _24783_, _24782_);
  and _29342_ (_07683_, _24784_, _22762_);
  and _29343_ (_24785_, _24722_, _23946_);
  and _29344_ (_24786_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  or _29345_ (_07737_, _24786_, _24785_);
  and _29346_ (_24787_, _24722_, _23707_);
  and _29347_ (_24788_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  or _29348_ (_07894_, _24788_, _24787_);
  and _29349_ (_24789_, _24356_, _24275_);
  and _29350_ (_24790_, _24789_, _23778_);
  not _29351_ (_24791_, _24789_);
  and _29352_ (_24792_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or _29353_ (_07925_, _24792_, _24790_);
  and _29354_ (_24793_, _24789_, _23747_);
  and _29355_ (_24794_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or _29356_ (_07944_, _24794_, _24793_);
  and _29357_ (_24795_, _24730_, _24705_);
  nand _29358_ (_24796_, _24795_, _23594_);
  or _29359_ (_24797_, _24795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _29360_ (_24798_, _24797_, _24737_);
  and _29361_ (_24799_, _24798_, _24796_);
  and _29362_ (_24800_, _24736_, _24043_);
  or _29363_ (_24801_, _24800_, _24799_);
  and _29364_ (_07995_, _24801_, _22762_);
  and _29365_ (_24802_, _24789_, _23649_);
  and _29366_ (_24803_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or _29367_ (_08032_, _24803_, _24802_);
  and _29368_ (_24804_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and _29369_ (_24805_, _24767_, _23824_);
  or _29370_ (_08049_, _24805_, _24804_);
  and _29371_ (_24806_, _24789_, _24050_);
  and _29372_ (_24807_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or _29373_ (_08086_, _24807_, _24806_);
  and _29374_ (_24808_, _24789_, _23707_);
  and _29375_ (_24809_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or _29376_ (_08131_, _24809_, _24808_);
  and _29377_ (_24810_, _24375_, _24050_);
  and _29378_ (_24811_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or _29379_ (_08161_, _24811_, _24810_);
  and _29380_ (_24812_, _23052_, _23034_);
  and _29381_ (_24813_, _24812_, _24729_);
  and _29382_ (_24814_, _24813_, _24296_);
  or _29383_ (_24815_, _24814_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _29384_ (_24816_, _24735_, _24064_);
  not _29385_ (_24817_, _24816_);
  and _29386_ (_24818_, _24817_, _24815_);
  nand _29387_ (_24819_, _24814_, _23594_);
  and _29388_ (_24820_, _24819_, _24818_);
  and _29389_ (_24821_, _24816_, _23642_);
  or _29390_ (_24822_, _24821_, _24820_);
  and _29391_ (_08221_, _24822_, _22762_);
  and _29392_ (_24823_, _24813_, _24291_);
  nand _29393_ (_24824_, _24823_, _23594_);
  or _29394_ (_24825_, _24823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _29395_ (_24826_, _24825_, _24817_);
  and _29396_ (_24827_, _24826_, _24824_);
  and _29397_ (_24828_, _24816_, _23816_);
  or _29398_ (_24829_, _24828_, _24827_);
  and _29399_ (_08240_, _24829_, _22762_);
  and _29400_ (_24830_, _24813_, _24678_);
  or _29401_ (_24831_, _24830_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _29402_ (_24832_, _24831_, _24817_);
  nand _29403_ (_24833_, _24830_, _23594_);
  and _29404_ (_24834_, _24833_, _24832_);
  and _29405_ (_24835_, _24816_, _24685_);
  or _29406_ (_24836_, _24835_, _24834_);
  and _29407_ (_08258_, _24836_, _22762_);
  and _29408_ (_24837_, _24375_, _23707_);
  and _29409_ (_24838_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or _29410_ (_27176_, _24838_, _24837_);
  and _29411_ (_24839_, _24370_, _24085_);
  and _29412_ (_24840_, _24839_, _23898_);
  not _29413_ (_24841_, _24839_);
  and _29414_ (_24842_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  or _29415_ (_08365_, _24842_, _24840_);
  and _29416_ (_24843_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and _29417_ (_24844_, _24767_, _23898_);
  or _29418_ (_08380_, _24844_, _24843_);
  or _29419_ (_24845_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _29420_ (_24846_, _24845_, _22762_);
  or _29421_ (_24847_, _24079_, _23642_);
  and _29422_ (_08395_, _24847_, _24846_);
  and _29423_ (_24848_, _24839_, _23824_);
  and _29424_ (_24849_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  or _29425_ (_08416_, _24849_, _24848_);
  and _29426_ (_24850_, _24839_, _23946_);
  and _29427_ (_24851_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  or _29428_ (_08466_, _24851_, _24850_);
  and _29429_ (_24852_, _23911_, _23076_);
  and _29430_ (_24853_, _24852_, _23649_);
  not _29431_ (_24854_, _24852_);
  and _29432_ (_24855_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  or _29433_ (_08496_, _24855_, _24853_);
  and _29434_ (_24856_, _24839_, _24050_);
  and _29435_ (_24857_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  or _29436_ (_08544_, _24857_, _24856_);
  and _29437_ (_24858_, _24370_, _24010_);
  and _29438_ (_24859_, _24858_, _23778_);
  not _29439_ (_24860_, _24858_);
  and _29440_ (_24861_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  or _29441_ (_08572_, _24861_, _24859_);
  and _29442_ (_24862_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _29443_ (_24863_, _24862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _29444_ (_24864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _29445_ (_24865_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _29446_ (_24866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _24865_);
  and _29447_ (_24867_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _29448_ (_24868_, _24867_, _24866_);
  and _29449_ (_24869_, _24868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor _29450_ (_24870_, _24869_, _24864_);
  not _29451_ (_24871_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _29452_ (_24872_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _29453_ (_24873_, _24872_, _24871_);
  nand _29454_ (_24874_, _24873_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not _29455_ (_24875_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _29456_ (_24876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor _29457_ (_24877_, _24876_, _24875_);
  and _29458_ (_24878_, _24877_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _29459_ (_24879_, _24878_);
  and _29460_ (_24880_, _24879_, _24874_);
  and _29461_ (_24881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _29462_ (_24882_, _24881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _29463_ (_24883_, _24882_);
  and _29464_ (_24884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _29465_ (_24885_, _24884_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _29466_ (_24886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _29467_ (_24887_, _24886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _29468_ (_24888_, _24887_, _24885_);
  and _29469_ (_24889_, _24888_, _24883_);
  and _29470_ (_24890_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _29471_ (_24891_, _24890_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _29472_ (_24892_, _24891_);
  and _29473_ (_24893_, _24892_, _24889_);
  and _29474_ (_24894_, _24893_, _24880_);
  nor _29475_ (_24895_, _24894_, _24870_);
  and _29476_ (_24896_, _24864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  not _29477_ (_24897_, _24896_);
  not _29478_ (_24898_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _29479_ (_24899_, _24873_, _24898_);
  not _29480_ (_24900_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _29481_ (_24901_, _24877_, _24900_);
  nor _29482_ (_24902_, _24901_, _24899_);
  not _29483_ (_24903_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _29484_ (_24904_, _24890_, _24903_);
  not _29485_ (_24905_, _24904_);
  not _29486_ (_24906_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _29487_ (_24907_, _24881_, _24906_);
  not _29488_ (_24908_, _24907_);
  not _29489_ (_24909_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _29490_ (_24910_, _24884_, _24909_);
  not _29491_ (_24911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _29492_ (_24912_, _24886_, _24911_);
  nor _29493_ (_24913_, _24912_, _24910_);
  and _29494_ (_24914_, _24913_, _24908_);
  and _29495_ (_24915_, _24914_, _24905_);
  and _29496_ (_24916_, _24915_, _24902_);
  or _29497_ (_24917_, _24916_, _24897_);
  nor _29498_ (_24918_, _24917_, _24895_);
  nand _29499_ (_24919_, _24918_, _24863_);
  and _29500_ (_24920_, _24895_, _24863_);
  or _29501_ (_24921_, _24920_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and _29502_ (_24922_, _24921_, _22762_);
  and _29503_ (_08672_, _24922_, _24919_);
  and _29504_ (_24923_, _24858_, _23898_);
  and _29505_ (_24924_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  or _29506_ (_27177_, _24924_, _24923_);
  and _29507_ (_24925_, _24858_, _23649_);
  and _29508_ (_24926_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  or _29509_ (_27178_, _24926_, _24925_);
  and _29510_ (_24927_, _24858_, _24050_);
  and _29511_ (_24928_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  or _29512_ (_08777_, _24928_, _24927_);
  nand _29513_ (_24929_, _24530_, _22767_);
  or _29514_ (_24930_, _22767_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _29515_ (_24931_, _24930_, _22762_);
  and _29516_ (_26864_[5], _24931_, _24929_);
  and _29517_ (_24932_, _24370_, _23911_);
  and _29518_ (_24933_, _24932_, _23898_);
  not _29519_ (_24934_, _24932_);
  and _29520_ (_24935_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or _29521_ (_08852_, _24935_, _24933_);
  and _29522_ (_24936_, _24932_, _23747_);
  and _29523_ (_24937_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or _29524_ (_08908_, _24937_, _24936_);
  nor _29525_ (_24938_, _24862_, _24865_);
  nand _29526_ (_24939_, _24938_, _24918_);
  and _29527_ (_24940_, _24938_, _24895_);
  or _29528_ (_24941_, _24940_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and _29529_ (_24942_, _24941_, _22762_);
  and _29530_ (_08926_, _24942_, _24939_);
  and _29531_ (_24943_, _24932_, _23946_);
  and _29532_ (_24944_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or _29533_ (_09009_, _24944_, _24943_);
  and _29534_ (_24945_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and _29535_ (_24946_, _24767_, _23946_);
  or _29536_ (_09056_, _24946_, _24945_);
  and _29537_ (_24947_, _24932_, _23707_);
  and _29538_ (_24948_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or _29539_ (_09081_, _24948_, _24947_);
  not _29540_ (_24949_, _24917_);
  nor _29541_ (_24950_, _24949_, _24895_);
  nor _29542_ (_24951_, _24950_, _24862_);
  not _29543_ (_24952_, _24951_);
  and _29544_ (_24953_, _24952_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _29545_ (_24954_, _24862_);
  nor _29546_ (_24955_, _24874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _29547_ (_24956_, _24955_, _24891_);
  not _29548_ (_24957_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _29549_ (_24958_, _24878_, _24865_);
  or _29550_ (_24959_, _24958_, _24957_);
  nand _29551_ (_24960_, _24959_, _24956_);
  and _29552_ (_24961_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _29553_ (_24962_, _24961_, _24892_);
  and _29554_ (_24963_, _24962_, _24960_);
  or _29555_ (_24964_, _24963_, _24887_);
  not _29556_ (_24965_, _24885_);
  not _29557_ (_24966_, _24887_);
  or _29558_ (_24967_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _24865_);
  or _29559_ (_24968_, _24967_, _24966_);
  and _29560_ (_24969_, _24968_, _24965_);
  and _29561_ (_24970_, _24969_, _24964_);
  and _29562_ (_24971_, _24961_, _24885_);
  or _29563_ (_24972_, _24971_, _24882_);
  or _29564_ (_24973_, _24972_, _24970_);
  or _29565_ (_24974_, _24967_, _24883_);
  and _29566_ (_24975_, _24974_, _24895_);
  and _29567_ (_24976_, _24975_, _24973_);
  or _29568_ (_24977_, _24967_, _24908_);
  and _29569_ (_24978_, _24899_, _24865_);
  nor _29570_ (_24979_, _24978_, _24904_);
  and _29571_ (_24980_, _24901_, _24865_);
  or _29572_ (_24981_, _24980_, _24957_);
  nand _29573_ (_24982_, _24981_, _24979_);
  or _29574_ (_24983_, _24961_, _24905_);
  and _29575_ (_24984_, _24983_, _24982_);
  or _29576_ (_24985_, _24984_, _24912_);
  not _29577_ (_24986_, _24910_);
  not _29578_ (_24987_, _24912_);
  or _29579_ (_24988_, _24967_, _24987_);
  and _29580_ (_24989_, _24988_, _24986_);
  and _29581_ (_24990_, _24989_, _24985_);
  and _29582_ (_24991_, _24961_, _24910_);
  or _29583_ (_24992_, _24991_, _24907_);
  or _29584_ (_24993_, _24992_, _24990_);
  and _29585_ (_24994_, _24993_, _24918_);
  and _29586_ (_24995_, _24994_, _24977_);
  or _29587_ (_24996_, _24995_, _24976_);
  and _29588_ (_24997_, _24996_, _24954_);
  or _29589_ (_24998_, _24997_, _24953_);
  and _29590_ (_09127_, _24998_, _22762_);
  and _29591_ (_24999_, _24370_, _24282_);
  and _29592_ (_25000_, _24999_, _23778_);
  not _29593_ (_25001_, _24999_);
  and _29594_ (_25002_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or _29595_ (_09156_, _25002_, _25000_);
  nand _29596_ (_25003_, _24950_, _24863_);
  nor _29597_ (_25004_, _24895_, _24862_);
  or _29598_ (_25005_, _25004_, _24865_);
  and _29599_ (_25006_, _25005_, _22762_);
  and _29600_ (_09190_, _25006_, _25003_);
  and _29601_ (_25007_, _24999_, _23747_);
  and _29602_ (_25008_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or _29603_ (_27183_, _25008_, _25007_);
  and _29604_ (_25009_, _24999_, _23946_);
  and _29605_ (_25010_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or _29606_ (_09277_, _25010_, _25009_);
  and _29607_ (_25011_, _24999_, _23707_);
  and _29608_ (_25012_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or _29609_ (_09338_, _25012_, _25011_);
  and _29610_ (_25013_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _29611_ (_25014_, _24236_, _24145_);
  nand _29612_ (_25015_, _25014_, _24153_);
  and _29613_ (_25016_, _25015_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  not _29614_ (_25017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _29615_ (_25018_, _25014_, _24256_);
  or _29616_ (_25019_, _25018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _29617_ (_25020_, _25019_, _25017_);
  or _29618_ (_25021_, _25020_, _25016_);
  nor _29619_ (_25022_, _24153_, _24182_);
  or _29620_ (_25023_, _25022_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _29621_ (_25024_, _25023_);
  and _29622_ (_25025_, _24235_, _24145_);
  and _29623_ (_25026_, _25025_, _25024_);
  or _29624_ (_25027_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _29625_ (_25028_, _25027_, _25021_);
  nor _29626_ (_25029_, _25028_, _24127_);
  and _29627_ (_25030_, _24127_, _23816_);
  or _29628_ (_25031_, _25030_, _25029_);
  and _29629_ (_25032_, _25031_, _24166_);
  or _29630_ (_09365_, _25032_, _25013_);
  and _29631_ (_25033_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and _29632_ (_25034_, _24767_, _24050_);
  or _29633_ (_09393_, _25034_, _25033_);
  not _29634_ (_25035_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor _29635_ (_25036_, _24951_, _25035_);
  or _29636_ (_25037_, _24892_, _24887_);
  and _29637_ (_25038_, _25037_, _24965_);
  and _29638_ (_25039_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _24865_);
  or _29639_ (_25040_, _25039_, _25038_);
  and _29640_ (_25041_, _24878_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _29641_ (_25042_, _25041_, _25035_);
  nor _29642_ (_25043_, _24874_, _24865_);
  nor _29643_ (_25044_, _25043_, _24891_);
  nand _29644_ (_25045_, _25044_, _24888_);
  or _29645_ (_25046_, _25045_, _25042_);
  and _29646_ (_25047_, _25046_, _25040_);
  or _29647_ (_25048_, _25047_, _24882_);
  or _29648_ (_25049_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _29649_ (_25050_, _24966_, _24885_);
  and _29650_ (_25051_, _25050_, _24883_);
  or _29651_ (_25052_, _25051_, _25049_);
  and _29652_ (_25053_, _25052_, _24895_);
  and _29653_ (_25054_, _25053_, _25048_);
  and _29654_ (_25055_, _24899_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _29655_ (_25056_, _25055_, _24904_);
  and _29656_ (_25057_, _24901_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _29657_ (_25058_, _25057_, _25035_);
  nand _29658_ (_25059_, _25058_, _25056_);
  or _29659_ (_25060_, _25039_, _24905_);
  and _29660_ (_25061_, _25060_, _25059_);
  or _29661_ (_25062_, _25061_, _24912_);
  or _29662_ (_25063_, _25049_, _24987_);
  and _29663_ (_25064_, _25063_, _24986_);
  and _29664_ (_25065_, _25064_, _25062_);
  and _29665_ (_25066_, _25039_, _24910_);
  or _29666_ (_25067_, _25066_, _24907_);
  or _29667_ (_25068_, _25067_, _25065_);
  and _29668_ (_25069_, _24918_, _24908_);
  and _29669_ (_25070_, _25049_, _24918_);
  or _29670_ (_25071_, _25070_, _25069_);
  and _29671_ (_25072_, _25071_, _25068_);
  or _29672_ (_25073_, _25072_, _25054_);
  and _29673_ (_25074_, _25073_, _24954_);
  or _29674_ (_25075_, _25074_, _25036_);
  and _29675_ (_09413_, _25075_, _22762_);
  and _29676_ (_25076_, _24852_, _23824_);
  and _29677_ (_25077_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  or _29678_ (_09433_, _25077_, _25076_);
  and _29679_ (_25078_, _23901_, _23655_);
  and _29680_ (_25079_, _25078_, _24370_);
  and _29681_ (_25080_, _25079_, _23778_);
  not _29682_ (_25081_, _25079_);
  and _29683_ (_25082_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  or _29684_ (_09490_, _25082_, _25080_);
  and _29685_ (_25083_, _25079_, _23824_);
  and _29686_ (_25084_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  or _29687_ (_09519_, _25084_, _25083_);
  and _29688_ (_25085_, _25079_, _23649_);
  and _29689_ (_25086_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  or _29690_ (_27185_, _25086_, _25085_);
  and _29691_ (_25087_, _25079_, _24050_);
  and _29692_ (_25088_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  or _29693_ (_09609_, _25088_, _25087_);
  and _29694_ (_25089_, _25079_, _23707_);
  and _29695_ (_25090_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  or _29696_ (_09650_, _25090_, _25089_);
  and _29697_ (_25091_, _24370_, _23656_);
  and _29698_ (_25092_, _25091_, _23824_);
  not _29699_ (_25093_, _25091_);
  and _29700_ (_25094_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  or _29701_ (_09680_, _25094_, _25092_);
  and _29702_ (_25095_, _24862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _29703_ (_25096_, _25095_, _24951_);
  and _29704_ (_09728_, _25096_, _22762_);
  nand _29705_ (_25097_, _24915_, _24896_);
  or _29706_ (_25098_, _25097_, _24902_);
  nor _29707_ (_25099_, _25098_, _24895_);
  and _29708_ (_25100_, _24862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  not _29709_ (_25101_, _24870_);
  nand _29710_ (_25102_, _24893_, _25101_);
  nor _29711_ (_25103_, _25102_, _24880_);
  and _29712_ (_25104_, _25103_, _24954_);
  or _29713_ (_25105_, _25104_, _25100_);
  or _29714_ (_25106_, _25105_, _25099_);
  and _29715_ (_09750_, _25106_, _22762_);
  nor _29716_ (_25108_, _24910_, _24907_);
  or _29717_ (_25109_, _24912_, _24904_);
  and _29718_ (_25110_, _24902_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _29719_ (_25111_, _25110_, _25109_);
  and _29720_ (_25112_, _25111_, _25108_);
  and _29721_ (_25113_, _25112_, _24918_);
  nor _29722_ (_25114_, _24885_, _24882_);
  or _29723_ (_25115_, _24891_, _24887_);
  and _29724_ (_25116_, _24880_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _29725_ (_25117_, _25116_, _25115_);
  and _29726_ (_25118_, _25117_, _25114_);
  and _29727_ (_25119_, _25118_, _24895_);
  or _29728_ (_25120_, _25119_, _25113_);
  or _29729_ (_25121_, _25120_, _24862_);
  or _29730_ (_25122_, _24954_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _29731_ (_25123_, _25122_, _22762_);
  and _29732_ (_09772_, _25123_, _25121_);
  nor _29733_ (_25125_, _24901_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _29734_ (_25126_, _25125_, _24899_);
  or _29735_ (_25127_, _25126_, _24904_);
  and _29736_ (_25128_, _25127_, _24987_);
  or _29737_ (_25129_, _25128_, _24910_);
  and _29738_ (_25130_, _25129_, _25069_);
  or _29739_ (_25131_, _24878_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _29740_ (_25132_, _25131_, _24874_);
  or _29741_ (_25133_, _25132_, _24891_);
  and _29742_ (_25134_, _25133_, _24966_);
  or _29743_ (_25135_, _25134_, _24885_);
  and _29744_ (_25136_, _24895_, _24883_);
  and _29745_ (_25137_, _25136_, _25135_);
  or _29746_ (_25138_, _25137_, _24862_);
  or _29747_ (_25139_, _25138_, _25130_);
  or _29748_ (_25140_, _24954_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _29749_ (_25141_, _25140_, _22762_);
  and _29750_ (_09791_, _25141_, _25139_);
  and _29751_ (_25142_, _24370_, _24275_);
  and _29752_ (_25143_, _25142_, _23778_);
  not _29753_ (_25144_, _25142_);
  and _29754_ (_25145_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  or _29755_ (_27199_, _25145_, _25143_);
  and _29756_ (_25146_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _22762_);
  and _29757_ (_09843_, _25146_, _24862_);
  and _29758_ (_25148_, _25091_, _23747_);
  and _29759_ (_25150_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  or _29760_ (_27187_, _25150_, _25148_);
  and _29761_ (_25151_, _25091_, _23946_);
  and _29762_ (_25153_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  or _29763_ (_09958_, _25153_, _25151_);
  and _29764_ (_25154_, _25091_, _23707_);
  and _29765_ (_25155_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  or _29766_ (_09981_, _25155_, _25154_);
  and _29767_ (_25156_, _24370_, _23752_);
  and _29768_ (_25157_, _25156_, _23898_);
  not _29769_ (_25158_, _25156_);
  and _29770_ (_25159_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or _29771_ (_10015_, _25159_, _25157_);
  and _29772_ (_25160_, _25156_, _23824_);
  and _29773_ (_25161_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or _29774_ (_10138_, _25161_, _25160_);
  nor _29775_ (_25162_, _23003_, _22970_);
  and _29776_ (_25163_, _25162_, _22943_);
  and _29777_ (_25164_, _25163_, _24643_);
  and _29778_ (_25165_, _25164_, _24118_);
  nand _29779_ (_25166_, _25165_, _23594_);
  or _29780_ (_25167_, _25165_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _29781_ (_25168_, _25167_, _24645_);
  and _29782_ (_25169_, _25168_, _25166_);
  and _29783_ (_25170_, _23065_, _23002_);
  and _29784_ (_25171_, _25170_, _24295_);
  and _29785_ (_25172_, _25171_, _24656_);
  and _29786_ (_25173_, _25172_, _23753_);
  not _29787_ (_25174_, _25173_);
  or _29788_ (_25175_, _25174_, _23738_);
  or _29789_ (_25176_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _29790_ (_25178_, _25176_, _24069_);
  and _29791_ (_25179_, _25178_, _25175_);
  not _29792_ (_25181_, _24068_);
  and _29793_ (_25182_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _29794_ (_25183_, _25182_, rst);
  or _29795_ (_25184_, _25183_, _25179_);
  or _29796_ (_10161_, _25184_, _25169_);
  and _29797_ (_25185_, _25164_, _24291_);
  nand _29798_ (_25186_, _25185_, _23594_);
  or _29799_ (_25187_, _25185_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _29800_ (_25188_, _25187_, _24645_);
  and _29801_ (_25189_, _25188_, _25186_);
  or _29802_ (_25190_, _25174_, _23816_);
  or _29803_ (_25191_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _29804_ (_25192_, _25191_, _24069_);
  and _29805_ (_25193_, _25192_, _25190_);
  and _29806_ (_25194_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _29807_ (_25195_, _25194_, rst);
  or _29808_ (_25196_, _25195_, _25193_);
  or _29809_ (_10186_, _25196_, _25189_);
  and _29810_ (_25197_, _25164_, _24067_);
  nand _29811_ (_25198_, _25197_, _23594_);
  or _29812_ (_25199_, _25197_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _29813_ (_25200_, _25199_, _24645_);
  and _29814_ (_25201_, _25200_, _25198_);
  or _29815_ (_25202_, _25174_, _23892_);
  or _29816_ (_25203_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _29817_ (_25204_, _25203_, _24069_);
  and _29818_ (_25205_, _25204_, _25202_);
  and _29819_ (_25206_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _29820_ (_25207_, _25206_, rst);
  or _29821_ (_25208_, _25207_, _25205_);
  or _29822_ (_10212_, _25208_, _25201_);
  and _29823_ (_25209_, _25164_, _24678_);
  nand _29824_ (_25210_, _25209_, _23594_);
  or _29825_ (_25211_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _29826_ (_25212_, _25211_, _24645_);
  and _29827_ (_25213_, _25212_, _25210_);
  nand _29828_ (_25214_, _25173_, _23772_);
  and _29829_ (_25215_, _25214_, _24069_);
  and _29830_ (_25216_, _25215_, _25211_);
  not _29831_ (_25217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor _29832_ (_25218_, _24068_, _25217_);
  or _29833_ (_25219_, _25218_, rst);
  or _29834_ (_25220_, _25219_, _25216_);
  or _29835_ (_10236_, _25220_, _25213_);
  and _29836_ (_25221_, _25156_, _23649_);
  and _29837_ (_25222_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or _29838_ (_10291_, _25222_, _25221_);
  and _29839_ (_25223_, _25156_, _24050_);
  and _29840_ (_25224_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or _29841_ (_27188_, _25224_, _25223_);
  and _29842_ (_25225_, _25164_, _24705_);
  nand _29843_ (_25226_, _25225_, _23594_);
  or _29844_ (_25227_, _25225_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _29845_ (_25228_, _25227_, _24645_);
  and _29846_ (_25229_, _25228_, _25226_);
  or _29847_ (_25230_, _25174_, _24043_);
  or _29848_ (_25231_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _29849_ (_25232_, _25231_, _24069_);
  and _29850_ (_25233_, _25232_, _25230_);
  not _29851_ (_25234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor _29852_ (_25235_, _24068_, _25234_);
  or _29853_ (_25236_, _25235_, rst);
  or _29854_ (_25237_, _25236_, _25233_);
  or _29855_ (_10409_, _25237_, _25229_);
  and _29856_ (_25238_, _25164_, _24125_);
  nand _29857_ (_25239_, _25238_, _23594_);
  or _29858_ (_25240_, _25238_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _29859_ (_25241_, _25240_, _24645_);
  and _29860_ (_25242_, _25241_, _25239_);
  or _29861_ (_25243_, _25174_, _23939_);
  or _29862_ (_25244_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _29863_ (_25245_, _25244_, _24069_);
  and _29864_ (_25246_, _25245_, _25243_);
  and _29865_ (_25247_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _29866_ (_25248_, _25247_, rst);
  or _29867_ (_25249_, _25248_, _25246_);
  or _29868_ (_10540_, _25249_, _25242_);
  and _29869_ (_25250_, _24358_, _23649_);
  and _29870_ (_25251_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  or _29871_ (_10604_, _25251_, _25250_);
  and _29872_ (_25252_, _24766_, _23991_);
  not _29873_ (_25253_, _25252_);
  and _29874_ (_25254_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  and _29875_ (_25255_, _25252_, _24050_);
  or _29876_ (_10628_, _25255_, _25254_);
  and _29877_ (_25256_, _24358_, _23747_);
  and _29878_ (_25257_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  or _29879_ (_10652_, _25257_, _25256_);
  and _29880_ (_25258_, _23002_, _22970_);
  and _29881_ (_25259_, _25258_, _22943_);
  and _29882_ (_25260_, _25259_, _24643_);
  and _29883_ (_25261_, _25260_, _24067_);
  nand _29884_ (_25262_, _25261_, _23594_);
  or _29885_ (_25263_, _25261_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _29886_ (_25264_, _25263_, _24645_);
  and _29887_ (_25265_, _25264_, _25262_);
  and _29888_ (_25266_, _25171_, _24734_);
  not _29889_ (_25267_, _25266_);
  or _29890_ (_25268_, _25267_, _23892_);
  or _29891_ (_25269_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _29892_ (_25270_, _25269_, _24069_);
  and _29893_ (_25271_, _25270_, _25268_);
  and _29894_ (_25272_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _29895_ (_25273_, _25272_, rst);
  or _29896_ (_25274_, _25273_, _25271_);
  or _29897_ (_10718_, _25274_, _25265_);
  and _29898_ (_25275_, _25260_, _24125_);
  nand _29899_ (_25276_, _25275_, _23594_);
  or _29900_ (_25277_, _25275_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _29901_ (_25278_, _25277_, _24645_);
  and _29902_ (_25279_, _25278_, _25276_);
  or _29903_ (_25280_, _25267_, _23939_);
  or _29904_ (_25281_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _29905_ (_25282_, _25281_, _24069_);
  and _29906_ (_25283_, _25282_, _25280_);
  and _29907_ (_25284_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _29908_ (_25286_, _25284_, rst);
  or _29909_ (_25287_, _25286_, _25283_);
  or _29910_ (_10757_, _25287_, _25279_);
  and _29911_ (_25289_, _25260_, _24296_);
  nand _29912_ (_25290_, _25289_, _23594_);
  or _29913_ (_25291_, _25289_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _29914_ (_25292_, _25291_, _24645_);
  and _29915_ (_25293_, _25292_, _25290_);
  or _29916_ (_25294_, _25267_, _23642_);
  or _29917_ (_25296_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _29918_ (_25297_, _25296_, _24069_);
  and _29919_ (_25299_, _25297_, _25294_);
  not _29920_ (_25300_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor _29921_ (_25301_, _24068_, _25300_);
  or _29922_ (_25302_, _25301_, rst);
  or _29923_ (_25303_, _25302_, _25299_);
  or _29924_ (_10779_, _25303_, _25293_);
  and _29925_ (_25304_, _25260_, _24118_);
  nand _29926_ (_25305_, _25304_, _23594_);
  or _29927_ (_25306_, _25304_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _29928_ (_25307_, _25306_, _24645_);
  and _29929_ (_25308_, _25307_, _25305_);
  or _29930_ (_25309_, _25267_, _23738_);
  or _29931_ (_25310_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _29932_ (_25311_, _25310_, _24069_);
  and _29933_ (_25312_, _25311_, _25309_);
  and _29934_ (_25313_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _29935_ (_25314_, _25313_, rst);
  or _29936_ (_25315_, _25314_, _25312_);
  or _29937_ (_10829_, _25315_, _25308_);
  and _29938_ (_25316_, _25260_, _24291_);
  nand _29939_ (_25317_, _25316_, _23594_);
  or _29940_ (_25318_, _25316_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _29941_ (_25319_, _25318_, _24645_);
  and _29942_ (_25320_, _25319_, _25317_);
  or _29943_ (_25321_, _25267_, _23816_);
  or _29944_ (_25322_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _29945_ (_25323_, _25322_, _24069_);
  and _29946_ (_25324_, _25323_, _25321_);
  and _29947_ (_25325_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _29948_ (_25326_, _25325_, rst);
  or _29949_ (_25327_, _25326_, _25324_);
  or _29950_ (_10855_, _25327_, _25320_);
  and _29951_ (_25328_, _25260_, _24678_);
  nand _29952_ (_25329_, _25328_, _23594_);
  or _29953_ (_25330_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _29954_ (_25331_, _25330_, _24645_);
  and _29955_ (_25332_, _25331_, _25329_);
  nand _29956_ (_25333_, _25266_, _23772_);
  and _29957_ (_25334_, _25333_, _24069_);
  and _29958_ (_25335_, _25334_, _25330_);
  not _29959_ (_25336_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor _29960_ (_25337_, _24068_, _25336_);
  or _29961_ (_25338_, _25337_, rst);
  or _29962_ (_25339_, _25338_, _25335_);
  or _29963_ (_10891_, _25339_, _25332_);
  and _29964_ (_25340_, _24356_, _23911_);
  and _29965_ (_25341_, _25340_, _23649_);
  not _29966_ (_25342_, _25340_);
  and _29967_ (_25343_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  or _29968_ (_27081_, _25343_, _25341_);
  and _29969_ (_25345_, _25340_, _23747_);
  and _29970_ (_25346_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  or _29971_ (_11051_, _25346_, _25345_);
  and _29972_ (_25348_, _25340_, _23824_);
  and _29973_ (_25349_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  or _29974_ (_11091_, _25349_, _25348_);
  and _29975_ (_25350_, _25163_, _24812_);
  and _29976_ (_25352_, _25350_, _24118_);
  nand _29977_ (_25353_, _25352_, _23594_);
  or _29978_ (_25354_, _25352_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _29979_ (_25355_, _25354_, _24645_);
  and _29980_ (_25356_, _25355_, _25353_);
  and _29981_ (_25358_, _25350_, _24678_);
  not _29982_ (_25359_, _25358_);
  or _29983_ (_25360_, _25359_, _23738_);
  or _29984_ (_25361_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _29985_ (_25362_, _25361_, _24069_);
  and _29986_ (_25363_, _25362_, _25360_);
  and _29987_ (_25364_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _29988_ (_25365_, _25364_, rst);
  or _29989_ (_25367_, _25365_, _25363_);
  or _29990_ (_11413_, _25367_, _25356_);
  and _29991_ (_25368_, _25350_, _24291_);
  nand _29992_ (_25369_, _25368_, _23594_);
  or _29993_ (_25370_, _25368_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _29994_ (_25371_, _25370_, _24645_);
  and _29995_ (_25372_, _25371_, _25369_);
  or _29996_ (_25373_, _25359_, _23816_);
  or _29997_ (_25374_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _29998_ (_25375_, _25374_, _24069_);
  and _29999_ (_25376_, _25375_, _25373_);
  and _30000_ (_25377_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _30001_ (_25378_, _25377_, rst);
  or _30002_ (_25379_, _25378_, _25376_);
  or _30003_ (_11482_, _25379_, _25372_);
  and _30004_ (_25380_, _25350_, _24067_);
  nand _30005_ (_25381_, _25380_, _23594_);
  or _30006_ (_25382_, _25380_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _30007_ (_25383_, _25382_, _24645_);
  and _30008_ (_25384_, _25383_, _25381_);
  or _30009_ (_25385_, _25359_, _23892_);
  or _30010_ (_25386_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _30011_ (_25387_, _25386_, _24069_);
  and _30012_ (_25388_, _25387_, _25385_);
  and _30013_ (_25389_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _30014_ (_25390_, _25389_, rst);
  or _30015_ (_25391_, _25390_, _25388_);
  or _30016_ (_11558_, _25391_, _25384_);
  nand _30017_ (_25393_, _25358_, _23594_);
  or _30018_ (_25394_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _30019_ (_25395_, _25394_, _24645_);
  and _30020_ (_25396_, _25395_, _25393_);
  nand _30021_ (_25397_, _25358_, _23772_);
  and _30022_ (_25398_, _25397_, _24069_);
  and _30023_ (_25399_, _25398_, _25394_);
  not _30024_ (_25400_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor _30025_ (_25401_, _24068_, _25400_);
  or _30026_ (_25402_, _25401_, rst);
  or _30027_ (_25403_, _25402_, _25399_);
  or _30028_ (_11583_, _25403_, _25396_);
  and _30029_ (_25404_, _25340_, _23707_);
  and _30030_ (_25405_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  or _30031_ (_11681_, _25405_, _25404_);
  and _30032_ (_25406_, _25340_, _24050_);
  and _30033_ (_25407_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  or _30034_ (_11792_, _25407_, _25406_);
  and _30035_ (_25408_, _25350_, _24705_);
  nand _30036_ (_25409_, _25408_, _23594_);
  or _30037_ (_25410_, _25408_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _30038_ (_25411_, _25410_, _24645_);
  and _30039_ (_25412_, _25411_, _25409_);
  or _30040_ (_25414_, _25359_, _24043_);
  or _30041_ (_25415_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _30042_ (_25416_, _25415_, _24069_);
  and _30043_ (_25417_, _25416_, _25414_);
  not _30044_ (_25418_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor _30045_ (_25419_, _24068_, _25418_);
  or _30046_ (_25420_, _25419_, rst);
  or _30047_ (_25421_, _25420_, _25417_);
  or _30048_ (_11878_, _25421_, _25412_);
  and _30049_ (_25422_, _25350_, _24125_);
  nand _30050_ (_25423_, _25422_, _23594_);
  or _30051_ (_25425_, _25422_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _30052_ (_25426_, _25425_, _24645_);
  and _30053_ (_25427_, _25426_, _25423_);
  or _30054_ (_25429_, _25359_, _23939_);
  or _30055_ (_25430_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _30056_ (_25431_, _25430_, _24069_);
  and _30057_ (_25432_, _25431_, _25429_);
  and _30058_ (_25433_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _30059_ (_25434_, _25433_, rst);
  or _30060_ (_25435_, _25434_, _25432_);
  or _30061_ (_11954_, _25435_, _25427_);
  and _30062_ (_25437_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  and _30063_ (_25438_, _25252_, _23898_);
  or _30064_ (_11987_, _25438_, _25437_);
  and _30065_ (_25439_, _25259_, _24812_);
  and _30066_ (_25441_, _25439_, _24291_);
  nand _30067_ (_25442_, _25441_, _23594_);
  or _30068_ (_25443_, _25441_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _30069_ (_25444_, _25443_, _24645_);
  and _30070_ (_25445_, _25444_, _25442_);
  and _30071_ (_25446_, _25171_, _24064_);
  not _30072_ (_25447_, _25446_);
  or _30073_ (_25448_, _25447_, _23816_);
  or _30074_ (_25449_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _30075_ (_25450_, _25449_, _24069_);
  and _30076_ (_25451_, _25450_, _25448_);
  and _30077_ (_25453_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _30078_ (_25455_, _25453_, rst);
  or _30079_ (_25456_, _25455_, _25451_);
  or _30080_ (_12139_, _25456_, _25445_);
  and _30081_ (_25459_, _25439_, _24067_);
  nand _30082_ (_25460_, _25459_, _23594_);
  or _30083_ (_25461_, _25459_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _30084_ (_25462_, _25461_, _24645_);
  and _30085_ (_25464_, _25462_, _25460_);
  or _30086_ (_25466_, _25447_, _23892_);
  or _30087_ (_25467_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _30088_ (_25468_, _25467_, _24069_);
  and _30089_ (_25469_, _25468_, _25466_);
  and _30090_ (_25470_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _30091_ (_25472_, _25470_, rst);
  or _30092_ (_25473_, _25472_, _25469_);
  or _30093_ (_12170_, _25473_, _25464_);
  and _30094_ (_25474_, _25439_, _24678_);
  nand _30095_ (_25475_, _25474_, _23594_);
  or _30096_ (_25476_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _30097_ (_25477_, _25476_, _24645_);
  and _30098_ (_25479_, _25477_, _25475_);
  nand _30099_ (_25480_, _25446_, _23772_);
  and _30100_ (_25481_, _25476_, _24069_);
  and _30101_ (_25482_, _25481_, _25480_);
  not _30102_ (_25483_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor _30103_ (_25484_, _24068_, _25483_);
  or _30104_ (_25485_, _25484_, rst);
  or _30105_ (_25486_, _25485_, _25482_);
  or _30106_ (_12192_, _25486_, _25479_);
  and _30107_ (_25488_, _24356_, _24010_);
  and _30108_ (_25489_, _25488_, _24050_);
  not _30109_ (_25490_, _25488_);
  and _30110_ (_25491_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or _30111_ (_12223_, _25491_, _25489_);
  and _30112_ (_25493_, _25488_, _23946_);
  and _30113_ (_25494_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or _30114_ (_12344_, _25494_, _25493_);
  and _30115_ (_25495_, _25439_, _24125_);
  nand _30116_ (_25496_, _25495_, _23594_);
  or _30117_ (_25497_, _25495_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _30118_ (_25498_, _25497_, _24645_);
  and _30119_ (_25499_, _25498_, _25496_);
  or _30120_ (_25500_, _25447_, _23939_);
  or _30121_ (_25501_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _30122_ (_25502_, _25501_, _24069_);
  and _30123_ (_25503_, _25502_, _25500_);
  and _30124_ (_25504_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _30125_ (_25505_, _25504_, rst);
  or _30126_ (_25506_, _25505_, _25503_);
  or _30127_ (_12395_, _25506_, _25499_);
  and _30128_ (_25507_, _25439_, _24705_);
  nand _30129_ (_25508_, _25507_, _23594_);
  or _30130_ (_25509_, _25507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _30131_ (_25510_, _25509_, _24645_);
  and _30132_ (_25511_, _25510_, _25508_);
  or _30133_ (_25512_, _25447_, _24043_);
  or _30134_ (_25514_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _30135_ (_25515_, _25514_, _24069_);
  and _30136_ (_25516_, _25515_, _25512_);
  not _30137_ (_25517_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor _30138_ (_25518_, _24068_, _25517_);
  or _30139_ (_25519_, _25518_, rst);
  or _30140_ (_25520_, _25519_, _25516_);
  or _30141_ (_12507_, _25520_, _25511_);
  and _30142_ (_25521_, _25439_, _24296_);
  nand _30143_ (_25523_, _25521_, _23594_);
  or _30144_ (_25524_, _25521_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _30145_ (_25525_, _25524_, _24645_);
  and _30146_ (_25526_, _25525_, _25523_);
  or _30147_ (_25527_, _25447_, _23642_);
  or _30148_ (_25528_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _30149_ (_25529_, _25528_, _24069_);
  and _30150_ (_25530_, _25529_, _25527_);
  not _30151_ (_25531_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor _30152_ (_25532_, _24068_, _25531_);
  or _30153_ (_25533_, _25532_, rst);
  or _30154_ (_25534_, _25533_, _25530_);
  or _30155_ (_12529_, _25534_, _25526_);
  and _30156_ (_25536_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  and _30157_ (_25537_, _25252_, _23747_);
  or _30158_ (_27043_, _25537_, _25536_);
  and _30159_ (_25538_, _25340_, _23778_);
  and _30160_ (_25539_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  or _30161_ (_27080_, _25539_, _25538_);
  and _30162_ (_25540_, _25488_, _23707_);
  and _30163_ (_25541_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or _30164_ (_12805_, _25541_, _25540_);
  and _30165_ (_25542_, _24766_, _23903_);
  not _30166_ (_25543_, _25542_);
  and _30167_ (_25544_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  and _30168_ (_25545_, _25542_, _23946_);
  or _30169_ (_12920_, _25545_, _25544_);
  and _30170_ (_25546_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  and _30171_ (_25547_, _25542_, _24050_);
  or _30172_ (_12950_, _25547_, _25546_);
  and _30173_ (_25548_, _25488_, _23898_);
  and _30174_ (_25549_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or _30175_ (_14450_, _25549_, _25548_);
  nor _30176_ (_25550_, _22768_, _23373_);
  and _30177_ (_25551_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _30178_ (_25552_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _30179_ (_25553_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or _30180_ (_25554_, _25553_, _25552_);
  and _30181_ (_25555_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _30182_ (_25556_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or _30183_ (_25557_, _25556_, _25555_);
  or _30184_ (_25558_, _25557_, _25554_);
  and _30185_ (_25559_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _30186_ (_25560_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _30187_ (_25561_, _25560_, _25559_);
  or _30188_ (_25562_, _25561_, _25558_);
  and _30189_ (_25563_, _25562_, _23839_);
  or _30190_ (_25564_, _25563_, _25551_);
  and _30191_ (_25565_, _25564_, _22768_);
  nor _30192_ (_25566_, _25565_, _25550_);
  nor _30193_ (_26897_[0], _25566_, rst);
  and _30194_ (_25568_, _25488_, _23778_);
  and _30195_ (_25570_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or _30196_ (_14601_, _25570_, _25568_);
  and _30197_ (_25571_, _24356_, _24085_);
  and _30198_ (_25572_, _25571_, _23707_);
  not _30199_ (_25573_, _25571_);
  and _30200_ (_25574_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or _30201_ (_14938_, _25574_, _25572_);
  or _30202_ (_25576_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _30203_ (_25577_, _25576_, _22762_);
  or _30204_ (_25579_, _24079_, _23939_);
  and _30205_ (_15132_, _25579_, _25577_);
  and _30206_ (_25581_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _30207_ (_25582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand _30208_ (_25583_, _25582_, _24152_);
  nor _30209_ (_25584_, _25583_, _24149_);
  and _30210_ (_25586_, _24234_, _25584_);
  and _30211_ (_25587_, _25586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _30212_ (_25588_, _25587_, _24145_);
  nand _30213_ (_25590_, _25588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _30214_ (_25591_, _25588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _30215_ (_25592_, _25591_, _24132_);
  and _30216_ (_25593_, _25592_, _25590_);
  and _30217_ (_25594_, _25019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _30218_ (_25595_, _24256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _30219_ (_25596_, _25595_, _25014_);
  or _30220_ (_25597_, _25596_, _25594_);
  nor _30221_ (_25598_, _25597_, _25593_);
  nor _30222_ (_25599_, _25598_, _24127_);
  and _30223_ (_25601_, _24127_, _23738_);
  or _30224_ (_25602_, _25601_, _25599_);
  and _30225_ (_25603_, _25602_, _24166_);
  or _30226_ (_15153_, _25603_, _25581_);
  and _30227_ (_25604_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  and _30228_ (_25605_, _25542_, _23707_);
  or _30229_ (_15784_, _25605_, _25604_);
  and _30230_ (_25607_, _25488_, _23747_);
  and _30231_ (_25608_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or _30232_ (_17267_, _25608_, _25607_);
  or _30233_ (_25609_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _30234_ (_25610_, _25609_, _22762_);
  or _30235_ (_25611_, _24079_, _24043_);
  and _30236_ (_17294_, _25611_, _25610_);
  and _30237_ (_25612_, _25488_, _23824_);
  and _30238_ (_25613_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or _30239_ (_17417_, _25613_, _25612_);
  and _30240_ (_25615_, _23755_, _23747_);
  and _30241_ (_25616_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  or _30242_ (_17600_, _25616_, _25615_);
  and _30243_ (_25618_, \oc8051_top_1.oc8051_sfr1.wait_data , _22762_);
  and _30244_ (_25619_, _25618_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _30245_ (_25620_, _24567_, _24552_);
  and _30246_ (_25621_, _24584_, _24471_);
  and _30247_ (_25622_, _25621_, _24448_);
  or _30248_ (_25623_, _25622_, _25620_);
  or _30249_ (_25624_, _25623_, _24568_);
  and _30250_ (_25625_, _24593_, _24471_);
  and _30251_ (_25626_, _25625_, _24567_);
  and _30252_ (_25627_, _24592_, _24538_);
  and _30253_ (_25629_, _25627_, _24567_);
  nor _30254_ (_25630_, _25629_, _25626_);
  and _30255_ (_25631_, _25621_, _24613_);
  and _30256_ (_25633_, _24618_, _24447_);
  nor _30257_ (_25634_, _25633_, _25631_);
  nand _30258_ (_25635_, _25634_, _25630_);
  and _30259_ (_25636_, _24552_, _24448_);
  and _30260_ (_25638_, _24598_, _24471_);
  and _30261_ (_25639_, _25638_, _24556_);
  or _30262_ (_25640_, _25639_, _25636_);
  or _30263_ (_25641_, _25640_, _25635_);
  or _30264_ (_25642_, _25641_, _25624_);
  and _30265_ (_25644_, _22768_, _22762_);
  and _30266_ (_25645_, _25644_, _25642_);
  or _30267_ (_26865_, _25645_, _25619_);
  and _30268_ (_25646_, _25571_, _23778_);
  and _30269_ (_25647_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or _30270_ (_17981_, _25647_, _25646_);
  and _30271_ (_25649_, _24010_, _23076_);
  and _30272_ (_25650_, _25649_, _23649_);
  not _30273_ (_25651_, _25649_);
  and _30274_ (_25652_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or _30275_ (_18188_, _25652_, _25650_);
  and _30276_ (_25653_, _25571_, _23898_);
  and _30277_ (_25654_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or _30278_ (_18303_, _25654_, _25653_);
  and _30279_ (_25656_, _24370_, _23069_);
  and _30280_ (_25657_, _25656_, _23946_);
  not _30281_ (_25659_, _25656_);
  and _30282_ (_25660_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or _30283_ (_18519_, _25660_, _25657_);
  not _30284_ (_25661_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _30285_ (_25662_, _24626_, _25661_);
  not _30286_ (_25663_, _24560_);
  and _30287_ (_25664_, _25663_, _25662_);
  nand _30288_ (_25665_, _24415_, _24412_);
  and _30289_ (_25666_, _25665_, _24408_);
  and _30290_ (_25667_, _25666_, _24554_);
  and _30291_ (_25668_, _25667_, _24552_);
  and _30292_ (_25669_, _25668_, _22767_);
  or _30293_ (_25671_, _25669_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _30294_ (_25672_, _25671_, _25664_);
  or _30295_ (_25674_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _22766_);
  and _30296_ (_25675_, _25674_, _22762_);
  and _30297_ (_26868_[2], _25675_, _25672_);
  and _30298_ (_25676_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _30299_ (_25677_, _24128_, _23939_);
  not _30300_ (_25678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _30301_ (_25679_, _24252_, _24256_);
  and _30302_ (_25680_, _24145_, _24131_);
  and _30303_ (_25681_, _24239_, _25680_);
  nand _30304_ (_25682_, _25681_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _30305_ (_25683_, _25682_, _24256_);
  nor _30306_ (_25684_, _25683_, _25679_);
  nor _30307_ (_25685_, _25684_, _25678_);
  and _30308_ (_25686_, _25683_, _25681_);
  and _30309_ (_25687_, _25014_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _30310_ (_25688_, _25687_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _30311_ (_25689_, _25688_, _25679_);
  or _30312_ (_25690_, _25689_, _25686_);
  or _30313_ (_25691_, _25690_, _25685_);
  or _30314_ (_25692_, _25691_, _24127_);
  and _30315_ (_25693_, _25692_, _24166_);
  and _30316_ (_25694_, _25693_, _25677_);
  or _30317_ (_18600_, _25694_, _25676_);
  and _30318_ (_25695_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  and _30319_ (_25696_, _25542_, _23778_);
  or _30320_ (_27042_, _25696_, _25695_);
  nor _30321_ (_25697_, _22768_, _23100_);
  and _30322_ (_25698_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _30323_ (_25699_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _30324_ (_25700_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _30325_ (_25701_, _25700_, _25699_);
  and _30326_ (_25702_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _30327_ (_25703_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _30328_ (_25704_, _25703_, _25702_);
  and _30329_ (_25705_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _30330_ (_25706_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _30331_ (_25707_, _25706_, _25705_);
  and _30332_ (_25708_, _25707_, _25704_);
  and _30333_ (_25709_, _25708_, _25701_);
  nor _30334_ (_25710_, _25709_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _30335_ (_25711_, _25710_, _25698_);
  nor _30336_ (_25712_, _25711_, _23950_);
  nor _30337_ (_25713_, _25712_, _25697_);
  nor _30338_ (_26897_[7], _25713_, rst);
  and _30339_ (_25714_, _25571_, _23747_);
  and _30340_ (_25715_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or _30341_ (_19421_, _25715_, _25714_);
  nor _30342_ (_25716_, _22768_, _23227_);
  and _30343_ (_25717_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _30344_ (_25718_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _30345_ (_25719_, _25718_, _25717_);
  and _30346_ (_25720_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _30347_ (_25721_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _30348_ (_25722_, _25721_, _25720_);
  and _30349_ (_25723_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _30350_ (_25724_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _30351_ (_25725_, _25724_, _25723_);
  and _30352_ (_25726_, _25725_, _25722_);
  and _30353_ (_25727_, _25726_, _25719_);
  and _30354_ (_25728_, _22768_, _23839_);
  not _30355_ (_25729_, _25728_);
  nor _30356_ (_25730_, _25729_, _25727_);
  nor _30357_ (_25731_, _25730_, _25716_);
  nor _30358_ (_26887_[4], _25731_, rst);
  and _30359_ (_25733_, _23986_, _23076_);
  and _30360_ (_25734_, _25733_, _23649_);
  not _30361_ (_25735_, _25733_);
  and _30362_ (_25736_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or _30363_ (_19920_, _25736_, _25734_);
  and _30364_ (_25737_, _23946_, _23755_);
  and _30365_ (_25738_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  or _30366_ (_19941_, _25738_, _25737_);
  and _30367_ (_25739_, _23903_, _23754_);
  and _30368_ (_25740_, _25739_, _23946_);
  not _30369_ (_25741_, _25739_);
  and _30370_ (_25742_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or _30371_ (_19972_, _25742_, _25740_);
  and _30372_ (_25743_, _25571_, _23649_);
  and _30373_ (_25744_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or _30374_ (_20043_, _25744_, _25743_);
  and _30375_ (_25745_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  and _30376_ (_25746_, _25542_, _23824_);
  or _30377_ (_20570_, _25746_, _25745_);
  and _30378_ (_25748_, _23784_, _23664_);
  and _30379_ (_25749_, _25748_, _23898_);
  not _30380_ (_25750_, _25748_);
  and _30381_ (_25751_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or _30382_ (_27069_, _25751_, _25749_);
  and _30383_ (_25752_, _24050_, _23790_);
  and _30384_ (_25753_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  or _30385_ (_27253_, _25753_, _25752_);
  and _30386_ (_25754_, _24356_, _23784_);
  and _30387_ (_25755_, _25754_, _23898_);
  not _30388_ (_25756_, _25754_);
  and _30389_ (_25757_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  or _30390_ (_21247_, _25757_, _25755_);
  and _30391_ (_25759_, _25754_, _23747_);
  and _30392_ (_25760_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  or _30393_ (_21348_, _25760_, _25759_);
  and _30394_ (_25761_, _25754_, _23824_);
  and _30395_ (_25762_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  or _30396_ (_21419_, _25762_, _25761_);
  and _30397_ (_26860_[4], _24464_, _22762_);
  and _30398_ (_25763_, _24766_, _24005_);
  not _30399_ (_25764_, _25763_);
  and _30400_ (_25765_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and _30401_ (_25766_, _25763_, _23946_);
  or _30402_ (_21820_, _25766_, _25765_);
  and _30403_ (_26885_[0], _24408_, _22762_);
  and _30404_ (_26885_[1], _24417_, _22762_);
  and _30405_ (_26885_[2], _24440_, _22762_);
  and _30406_ (_25769_, _23052_, _22971_);
  and _30407_ (_25770_, _25171_, _24069_);
  and _30408_ (_25772_, _25770_, _25769_);
  and _30409_ (_25773_, _25772_, _23662_);
  not _30410_ (_25774_, _25773_);
  and _30411_ (_25775_, _25774_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _30412_ (_25776_, _25769_, _23662_);
  and _30413_ (_25777_, _25776_, _25770_);
  and _30414_ (_25779_, _25777_, _23738_);
  nor _30415_ (_25780_, _25779_, _25775_);
  nor _30416_ (_26885_[3], _25780_, rst);
  or _30417_ (_25782_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  not _30418_ (_25783_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nand _30419_ (_25784_, _23953_, _25783_);
  and _30420_ (_25785_, _25784_, _22762_);
  and _30421_ (_26903_[0], _25785_, _25782_);
  or _30422_ (_25787_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  not _30423_ (_25788_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand _30424_ (_25789_, _23953_, _25788_);
  and _30425_ (_25790_, _25789_, _22762_);
  and _30426_ (_26903_[1], _25790_, _25787_);
  or _30427_ (_25791_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  not _30428_ (_25793_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand _30429_ (_25794_, _23953_, _25793_);
  and _30430_ (_25795_, _25794_, _22762_);
  and _30431_ (_26903_[2], _25795_, _25791_);
  or _30432_ (_25797_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  not _30433_ (_25798_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nand _30434_ (_25799_, _23953_, _25798_);
  and _30435_ (_25801_, _25799_, _22762_);
  and _30436_ (_26903_[3], _25801_, _25797_);
  or _30437_ (_25802_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  not _30438_ (_25803_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nand _30439_ (_25804_, _23953_, _25803_);
  and _30440_ (_25805_, _25804_, _22762_);
  and _30441_ (_26903_[4], _25805_, _25802_);
  or _30442_ (_25806_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  not _30443_ (_25807_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nand _30444_ (_25808_, _23953_, _25807_);
  and _30445_ (_25809_, _25808_, _22762_);
  and _30446_ (_26903_[5], _25809_, _25806_);
  or _30447_ (_25810_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  not _30448_ (_25811_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand _30449_ (_25812_, _23953_, _25811_);
  and _30450_ (_25813_, _25812_, _22762_);
  and _30451_ (_26903_[6], _25813_, _25810_);
  or _30452_ (_25816_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  not _30453_ (_25817_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nand _30454_ (_25818_, _23953_, _25817_);
  and _30455_ (_25820_, _25818_, _22762_);
  and _30456_ (_26903_[7], _25820_, _25816_);
  or _30457_ (_25821_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  not _30458_ (_25822_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand _30459_ (_25823_, _23953_, _25822_);
  and _30460_ (_25824_, _25823_, _22762_);
  and _30461_ (_26903_[8], _25824_, _25821_);
  or _30462_ (_25825_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  not _30463_ (_25826_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand _30464_ (_25827_, _23953_, _25826_);
  and _30465_ (_25828_, _25827_, _22762_);
  and _30466_ (_26903_[9], _25828_, _25825_);
  or _30467_ (_25829_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  not _30468_ (_25830_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand _30469_ (_25831_, _23953_, _25830_);
  and _30470_ (_25832_, _25831_, _22762_);
  and _30471_ (_26903_[10], _25832_, _25829_);
  or _30472_ (_25833_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  not _30473_ (_25834_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand _30474_ (_25835_, _23953_, _25834_);
  and _30475_ (_25836_, _25835_, _22762_);
  and _30476_ (_26903_[11], _25836_, _25833_);
  or _30477_ (_25837_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  not _30478_ (_25838_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nand _30479_ (_25839_, _23953_, _25838_);
  and _30480_ (_25840_, _25839_, _22762_);
  and _30481_ (_26903_[12], _25840_, _25837_);
  or _30482_ (_25841_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  not _30483_ (_25842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand _30484_ (_25843_, _23953_, _25842_);
  and _30485_ (_25844_, _25843_, _22762_);
  and _30486_ (_26903_[13], _25844_, _25841_);
  or _30487_ (_25845_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  not _30488_ (_25846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand _30489_ (_25847_, _23953_, _25846_);
  and _30490_ (_25848_, _25847_, _22762_);
  and _30491_ (_26903_[14], _25848_, _25845_);
  or _30492_ (_25849_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  not _30493_ (_25850_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand _30494_ (_25851_, _23953_, _25850_);
  and _30495_ (_25852_, _25851_, _22762_);
  and _30496_ (_26903_[15], _25852_, _25849_);
  or _30497_ (_25853_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  not _30498_ (_25854_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand _30499_ (_25855_, _23953_, _25854_);
  and _30500_ (_25856_, _25855_, _22762_);
  and _30501_ (_26903_[16], _25856_, _25853_);
  or _30502_ (_25857_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  not _30503_ (_25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand _30504_ (_25859_, _23953_, _25858_);
  and _30505_ (_25860_, _25859_, _22762_);
  and _30506_ (_26903_[17], _25860_, _25857_);
  or _30507_ (_25861_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  not _30508_ (_25862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand _30509_ (_25863_, _23953_, _25862_);
  and _30510_ (_25864_, _25863_, _22762_);
  and _30511_ (_26903_[18], _25864_, _25861_);
  or _30512_ (_25865_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  not _30513_ (_25866_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand _30514_ (_25867_, _23953_, _25866_);
  and _30515_ (_25868_, _25867_, _22762_);
  and _30516_ (_26903_[19], _25868_, _25865_);
  or _30517_ (_25869_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  not _30518_ (_25870_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand _30519_ (_25871_, _23953_, _25870_);
  and _30520_ (_25873_, _25871_, _22762_);
  and _30521_ (_26903_[20], _25873_, _25869_);
  or _30522_ (_25875_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  not _30523_ (_25876_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand _30524_ (_25877_, _23953_, _25876_);
  and _30525_ (_25878_, _25877_, _22762_);
  and _30526_ (_26903_[21], _25878_, _25875_);
  or _30527_ (_25879_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  not _30528_ (_25880_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand _30529_ (_25881_, _23953_, _25880_);
  and _30530_ (_25882_, _25881_, _22762_);
  and _30531_ (_26903_[22], _25882_, _25879_);
  or _30532_ (_25883_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  not _30533_ (_25884_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand _30534_ (_25885_, _23953_, _25884_);
  and _30535_ (_25886_, _25885_, _22762_);
  and _30536_ (_26903_[23], _25886_, _25883_);
  and _30537_ (_25887_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  not _30538_ (_25888_, _23953_);
  and _30539_ (_25889_, _25888_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or _30540_ (_25890_, _25889_, _25887_);
  and _30541_ (_26903_[24], _25890_, _22762_);
  or _30542_ (_25891_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  not _30543_ (_25892_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand _30544_ (_25893_, _23953_, _25892_);
  and _30545_ (_25894_, _25893_, _22762_);
  and _30546_ (_26903_[25], _25894_, _25891_);
  or _30547_ (_25895_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  not _30548_ (_25896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand _30549_ (_25897_, _23953_, _25896_);
  and _30550_ (_25898_, _25897_, _22762_);
  and _30551_ (_26903_[26], _25898_, _25895_);
  or _30552_ (_25899_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  not _30553_ (_25900_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand _30554_ (_25901_, _23953_, _25900_);
  and _30555_ (_25902_, _25901_, _22762_);
  and _30556_ (_26903_[27], _25902_, _25899_);
  or _30557_ (_25903_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  not _30558_ (_25904_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand _30559_ (_25905_, _23953_, _25904_);
  and _30560_ (_25906_, _25905_, _22762_);
  and _30561_ (_26903_[28], _25906_, _25903_);
  or _30562_ (_25907_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  not _30563_ (_25908_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand _30564_ (_25909_, _23953_, _25908_);
  and _30565_ (_25910_, _25909_, _22762_);
  and _30566_ (_26903_[29], _25910_, _25907_);
  or _30567_ (_25911_, _23953_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  not _30568_ (_25912_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand _30569_ (_25913_, _23953_, _25912_);
  and _30570_ (_25914_, _25913_, _22762_);
  and _30571_ (_26903_[30], _25914_, _25911_);
  and _30572_ (_25915_, _25754_, _24050_);
  and _30573_ (_25916_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  or _30574_ (_22542_, _25916_, _25915_);
  and _30575_ (_25917_, _25774_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _30576_ (_25918_, _25777_, _23642_);
  nor _30577_ (_25919_, _25918_, _25917_);
  nor _30578_ (_25920_, _25919_, _22971_);
  and _30579_ (_25921_, _25919_, _22971_);
  nor _30580_ (_25922_, _25921_, _25920_);
  nor _30581_ (_25923_, _24408_, _23018_);
  and _30582_ (_25924_, _24408_, _23018_);
  nor _30583_ (_25925_, _25924_, _25923_);
  and _30584_ (_25926_, _22905_, _22948_);
  and _30585_ (_25927_, _25926_, _23052_);
  and _30586_ (_25928_, _25927_, _24066_);
  and _30587_ (_25929_, _25928_, _23073_);
  and _30588_ (_25930_, _25929_, _25925_);
  and _30589_ (_25931_, _25780_, _23003_);
  nor _30590_ (_25932_, _25780_, _23003_);
  nor _30591_ (_25933_, _25932_, _25931_);
  and _30592_ (_25934_, _25933_, _25930_);
  and _30593_ (_25935_, _25934_, _25922_);
  and _30594_ (_25936_, _25780_, _24408_);
  and _30595_ (_25937_, _25936_, _25919_);
  and _30596_ (_25938_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _30597_ (_25939_, _25780_, _24612_);
  and _30598_ (_25940_, _25939_, _25919_);
  and _30599_ (_25941_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor _30600_ (_25942_, _25941_, _25938_);
  nor _30601_ (_25943_, _25780_, _24612_);
  and _30602_ (_25945_, _25943_, _25919_);
  and _30603_ (_25946_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor _30604_ (_25947_, _25780_, _24408_);
  and _30605_ (_25948_, _25947_, _25919_);
  and _30606_ (_25949_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _30607_ (_25950_, _25949_, _25946_);
  and _30608_ (_25952_, _25950_, _25942_);
  not _30609_ (_25953_, _25919_);
  and _30610_ (_25954_, _25947_, _25953_);
  and _30611_ (_25955_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _30612_ (_25956_, _25943_, _25953_);
  and _30613_ (_25957_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor _30614_ (_25958_, _25957_, _25955_);
  and _30615_ (_25959_, _25939_, _25953_);
  and _30616_ (_25960_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _30617_ (_25961_, _25936_, _25953_);
  and _30618_ (_25962_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor _30619_ (_25963_, _25962_, _25960_);
  and _30620_ (_25964_, _25963_, _25958_);
  and _30621_ (_25965_, _25964_, _25952_);
  nor _30622_ (_25966_, _25965_, _25935_);
  and _30623_ (_25967_, _25935_, _24685_);
  nor _30624_ (_25968_, _25967_, _25966_);
  nor _30625_ (_26886_[0], _25968_, rst);
  and _30626_ (_25969_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _30627_ (_25970_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor _30628_ (_25971_, _25970_, _25969_);
  and _30629_ (_25973_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _30630_ (_25974_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor _30631_ (_25975_, _25974_, _25973_);
  and _30632_ (_25976_, _25975_, _25971_);
  and _30633_ (_25977_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _30634_ (_25978_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _30635_ (_25979_, _25978_, _25977_);
  and _30636_ (_25980_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _30637_ (_25981_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor _30638_ (_25982_, _25981_, _25980_);
  and _30639_ (_25983_, _25982_, _25979_);
  and _30640_ (_25984_, _25983_, _25976_);
  nor _30641_ (_25985_, _25984_, _25935_);
  and _30642_ (_25986_, _25935_, _23892_);
  nor _30643_ (_25987_, _25986_, _25985_);
  nor _30644_ (_26886_[1], _25987_, rst);
  and _30645_ (_25988_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _30646_ (_25989_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor _30647_ (_25990_, _25989_, _25988_);
  and _30648_ (_25991_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _30649_ (_25992_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _30650_ (_25993_, _25992_, _25991_);
  and _30651_ (_25994_, _25993_, _25990_);
  and _30652_ (_25995_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _30653_ (_25996_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor _30654_ (_25997_, _25996_, _25995_);
  and _30655_ (_25998_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and _30656_ (_26000_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor _30657_ (_26001_, _26000_, _25998_);
  and _30658_ (_26002_, _26001_, _25997_);
  and _30659_ (_26003_, _26002_, _25994_);
  nor _30660_ (_26004_, _26003_, _25935_);
  and _30661_ (_26005_, _25935_, _23816_);
  nor _30662_ (_26006_, _26005_, _26004_);
  nor _30663_ (_26886_[2], _26006_, rst);
  and _30664_ (_26007_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _30665_ (_26008_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor _30666_ (_26009_, _26008_, _26007_);
  and _30667_ (_26010_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _30668_ (_26011_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor _30669_ (_26012_, _26011_, _26010_);
  and _30670_ (_26013_, _26012_, _26009_);
  and _30671_ (_26014_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _30672_ (_26015_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor _30673_ (_26016_, _26015_, _26014_);
  and _30674_ (_26017_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and _30675_ (_26018_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _30676_ (_26019_, _26018_, _26017_);
  and _30677_ (_26020_, _26019_, _26016_);
  and _30678_ (_26021_, _26020_, _26013_);
  nor _30679_ (_26022_, _26021_, _25935_);
  and _30680_ (_26023_, _25935_, _23738_);
  nor _30681_ (_26024_, _26023_, _26022_);
  nor _30682_ (_26886_[3], _26024_, rst);
  and _30683_ (_26026_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _30684_ (_26027_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor _30685_ (_26028_, _26027_, _26026_);
  and _30686_ (_26029_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _30687_ (_26030_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor _30688_ (_26031_, _26030_, _26029_);
  and _30689_ (_26032_, _26031_, _26028_);
  and _30690_ (_26033_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _30691_ (_26034_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor _30692_ (_26035_, _26034_, _26033_);
  and _30693_ (_26036_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _30694_ (_26037_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _30695_ (_26038_, _26037_, _26036_);
  and _30696_ (_26039_, _26038_, _26035_);
  and _30697_ (_26040_, _26039_, _26032_);
  nor _30698_ (_26041_, _26040_, _25935_);
  and _30699_ (_26042_, _25935_, _23642_);
  nor _30700_ (_26043_, _26042_, _26041_);
  nor _30701_ (_26886_[4], _26043_, rst);
  and _30702_ (_26044_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _30703_ (_26045_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor _30704_ (_26046_, _26045_, _26044_);
  and _30705_ (_26047_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _30706_ (_26048_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor _30707_ (_26049_, _26048_, _26047_);
  and _30708_ (_26051_, _26049_, _26046_);
  and _30709_ (_26052_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _30710_ (_26053_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor _30711_ (_26055_, _26053_, _26052_);
  and _30712_ (_26056_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _30713_ (_26058_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor _30714_ (_26060_, _26058_, _26056_);
  and _30715_ (_26061_, _26060_, _26055_);
  and _30716_ (_26062_, _26061_, _26051_);
  nor _30717_ (_26063_, _26062_, _25935_);
  and _30718_ (_26064_, _25935_, _23939_);
  nor _30719_ (_26065_, _26064_, _26063_);
  nor _30720_ (_26886_[5], _26065_, rst);
  and _30721_ (_26067_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and _30722_ (_26069_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor _30723_ (_26070_, _26069_, _26067_);
  and _30724_ (_26072_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _30725_ (_26073_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor _30726_ (_26074_, _26073_, _26072_);
  and _30727_ (_26075_, _26074_, _26070_);
  and _30728_ (_26076_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and _30729_ (_26077_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nor _30730_ (_26078_, _26077_, _26076_);
  and _30731_ (_26079_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _30732_ (_26080_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor _30733_ (_26082_, _26080_, _26079_);
  and _30734_ (_26083_, _26082_, _26078_);
  and _30735_ (_26084_, _26083_, _26075_);
  nor _30736_ (_26085_, _26084_, _25935_);
  and _30737_ (_26086_, _25935_, _24043_);
  nor _30738_ (_26088_, _26086_, _26085_);
  nor _30739_ (_26886_[6], _26088_, rst);
  and _30740_ (_26089_, _23824_, _23755_);
  and _30741_ (_26090_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  or _30742_ (_22628_, _26090_, _26089_);
  and _30743_ (_26091_, _25754_, _23946_);
  and _30744_ (_26092_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  or _30745_ (_22629_, _26092_, _26091_);
  and _30746_ (_26094_, _25754_, _23649_);
  and _30747_ (_26095_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  or _30748_ (_27034_, _26095_, _26094_);
  nand _30749_ (_26096_, _24293_, _23702_);
  nor _30750_ (_26097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not _30751_ (_26098_, _26097_);
  not _30752_ (_26099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _30753_ (_26100_, _26099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _30754_ (_26101_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  not _30755_ (_26102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not _30756_ (_26103_, t0_i);
  and _30757_ (_26104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _26103_);
  nor _30758_ (_26105_, _26104_, _26102_);
  not _30759_ (_26106_, _26105_);
  not _30760_ (_26107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _30761_ (_26108_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor _30762_ (_26109_, _26108_, _26107_);
  and _30763_ (_26110_, _26109_, _26106_);
  and _30764_ (_26111_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _30765_ (_26112_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _30766_ (_26113_, _26112_, _26111_);
  and _30767_ (_26114_, _26113_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _30768_ (_26115_, _26114_, _26110_);
  and _30769_ (_26116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _30770_ (_26117_, _26116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _30771_ (_26118_, _26117_, _26115_);
  nor _30772_ (_26119_, _26118_, _26097_);
  nor _30773_ (_26120_, _26119_, _26101_);
  nand _30774_ (_26121_, _26120_, _26098_);
  or _30775_ (_26122_, _26121_, _24299_);
  and _30776_ (_26123_, _26122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _30777_ (_26124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand _30778_ (_26125_, _26124_, _26115_);
  or _30779_ (_26126_, _26125_, _26120_);
  nor _30780_ (_26127_, _26126_, _24299_);
  or _30781_ (_26128_, _26127_, _26123_);
  or _30782_ (_26129_, _26128_, _24293_);
  and _30783_ (_26130_, _26129_, _22762_);
  and _30784_ (_22630_, _26130_, _26096_);
  nor _30785_ (_26131_, _22768_, _23275_);
  and _30786_ (_26133_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _30787_ (_26134_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _30788_ (_26135_, _26134_, _26133_);
  and _30789_ (_26136_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _30790_ (_26137_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _30791_ (_26138_, _26137_, _26136_);
  and _30792_ (_26139_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _30793_ (_26140_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _30794_ (_26141_, _26140_, _26139_);
  and _30795_ (_26142_, _26141_, _26138_);
  and _30796_ (_26143_, _26142_, _26135_);
  nor _30797_ (_26144_, _26143_, _25729_);
  nor _30798_ (_26145_, _26144_, _26131_);
  nor _30799_ (_26887_[3], _26145_, rst);
  nor _30800_ (_26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _30801_ (_26147_, _26146_, _23392_);
  nor _30802_ (_26148_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor _30803_ (_26149_, _26148_, _26147_);
  and _30804_ (_26150_, _23397_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _30805_ (_26151_, _26150_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _30806_ (_26152_, _23179_, _23141_);
  nor _30807_ (_26153_, _26152_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _30808_ (_26154_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _30809_ (_26155_, _23462_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _30810_ (_26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _30811_ (_26157_, _23216_, _26156_);
  nand _30812_ (_26158_, _26157_, _26155_);
  or _30813_ (_26159_, _23250_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _30814_ (_26160_, _23177_, _26156_);
  nand _30815_ (_26161_, _26160_, _26159_);
  and _30816_ (_26162_, _26161_, _26158_);
  or _30817_ (_26163_, _23332_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _30818_ (_26164_, _23250_, _26156_);
  nand _30819_ (_26165_, _26164_, _26163_);
  or _30820_ (_26166_, _23216_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _30821_ (_26167_, _23141_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _30822_ (_26168_, _26167_, _26166_);
  and _30823_ (_26169_, _26168_, _26165_);
  nand _30824_ (_26170_, _26169_, _26162_);
  and _30825_ (_26171_, _26170_, _26154_);
  nor _30826_ (_26172_, _26171_, _26153_);
  or _30827_ (_26173_, _23364_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _30828_ (_26174_, _23462_, _26156_);
  nand _30829_ (_26175_, _26174_, _26173_);
  and _30830_ (_26176_, _26175_, _26154_);
  and _30831_ (_26177_, _26168_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _30832_ (_26178_, _26177_, _26176_);
  not _30833_ (_26179_, _26178_);
  nor _30834_ (_26180_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not _30835_ (_26181_, _26180_);
  nand _30836_ (_26182_, _26146_, _23131_);
  and _30837_ (_26183_, _26182_, _26181_);
  not _30838_ (_26184_, _26183_);
  or _30839_ (_26185_, _23397_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _30840_ (_26186_, _23332_, _26156_);
  and _30841_ (_26187_, _26186_, _26185_);
  or _30842_ (_26188_, _26187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _30843_ (_26189_, _26161_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _30844_ (_26190_, _26189_, _26188_);
  or _30845_ (_26191_, _26190_, _26184_);
  and _30846_ (_26192_, _23364_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _30847_ (_26193_, _26192_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _30848_ (_26194_, _26158_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _30849_ (_26195_, _26194_, _26193_);
  nor _30850_ (_26196_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not _30851_ (_26197_, _26196_);
  nand _30852_ (_26198_, _26146_, _23171_);
  and _30853_ (_26199_, _26198_, _26197_);
  not _30854_ (_26200_, _26199_);
  or _30855_ (_26201_, _26200_, _26195_);
  nand _30856_ (_26202_, _26189_, _26188_);
  or _30857_ (_26203_, _26202_, _26183_);
  and _30858_ (_26204_, _26203_, _26191_);
  not _30859_ (_26205_, _26204_);
  or _30860_ (_26206_, _26205_, _26201_);
  and _30861_ (_26207_, _26206_, _26191_);
  nand _30862_ (_26208_, _26194_, _26193_);
  or _30863_ (_26209_, _26199_, _26208_);
  and _30864_ (_26210_, _26209_, _26201_);
  and _30865_ (_26211_, _26210_, _26204_);
  nor _30866_ (_26212_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not _30867_ (_26213_, _26212_);
  not _30868_ (_26214_, _26146_);
  or _30869_ (_26215_, _26214_, _23208_);
  nand _30870_ (_26216_, _26215_, _26213_);
  or _30871_ (_26217_, _26150_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _30872_ (_26218_, _26165_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _30873_ (_26219_, _26218_, _26217_);
  or _30874_ (_26220_, _26219_, _26216_);
  nor _30875_ (_26221_, _26175_, _26154_);
  nand _30876_ (_26222_, _26146_, _23244_);
  nor _30877_ (_26223_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not _30878_ (_26224_, _26223_);
  and _30879_ (_26225_, _26224_, _26222_);
  not _30880_ (_26226_, _26225_);
  or _30881_ (_26227_, _26226_, _26221_);
  and _30882_ (_26228_, _26215_, _26213_);
  nand _30883_ (_26229_, _26218_, _26217_);
  or _30884_ (_26230_, _26229_, _26228_);
  nand _30885_ (_26231_, _26230_, _26220_);
  or _30886_ (_26232_, _26231_, _26227_);
  nand _30887_ (_26233_, _26232_, _26220_);
  nand _30888_ (_26234_, _26233_, _26211_);
  and _30889_ (_26235_, _26234_, _26207_);
  and _30890_ (_26236_, _26187_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _30891_ (_26237_, _26236_);
  nor _30892_ (_26238_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not _30893_ (_26239_, _26238_);
  nand _30894_ (_26240_, _26146_, _23291_);
  and _30895_ (_26241_, _26240_, _26239_);
  nand _30896_ (_26242_, _26241_, _26237_);
  or _30897_ (_26243_, _26241_, _26237_);
  nand _30898_ (_26244_, _26243_, _26242_);
  nand _30899_ (_26245_, _26192_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _30900_ (_26246_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not _30901_ (_26247_, _26246_);
  or _30902_ (_26248_, _26214_, _23326_);
  and _30903_ (_26249_, _26248_, _26247_);
  nand _30904_ (_26250_, _26249_, _26245_);
  nor _30905_ (_26251_, _26146_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not _30906_ (_26252_, _26251_);
  or _30907_ (_26253_, _26214_, _23359_);
  nand _30908_ (_26254_, _26253_, _26252_);
  and _30909_ (_26255_, _26254_, _26151_);
  or _30910_ (_26256_, _26249_, _26245_);
  nand _30911_ (_26257_, _26256_, _26250_);
  or _30912_ (_26258_, _26257_, _26255_);
  and _30913_ (_26259_, _26258_, _26250_);
  or _30914_ (_26260_, _26259_, _26244_);
  nand _30915_ (_26261_, _26260_, _26242_);
  not _30916_ (_26262_, _26221_);
  or _30917_ (_26263_, _26225_, _26262_);
  and _30918_ (_26264_, _26263_, _26227_);
  and _30919_ (_26265_, _26230_, _26220_);
  and _30920_ (_26266_, _26265_, _26264_);
  and _30921_ (_26267_, _26266_, _26211_);
  nand _30922_ (_26268_, _26267_, _26261_);
  nand _30923_ (_26269_, _26268_, _26235_);
  and _30924_ (_26270_, _26179_, _26172_);
  nand _30925_ (_26271_, _26270_, _26269_);
  and _30926_ (_26272_, _26271_, _26184_);
  not _30927_ (_26273_, _26272_);
  and _30928_ (_26274_, _26270_, _26269_);
  and _30929_ (_26275_, _26219_, _26216_);
  not _30930_ (_26276_, _26227_);
  and _30931_ (_26277_, _26264_, _26261_);
  nor _30932_ (_26278_, _26277_, _26276_);
  or _30933_ (_26279_, _26278_, _26275_);
  and _30934_ (_26280_, _26279_, _26220_);
  not _30935_ (_26281_, _26280_);
  nand _30936_ (_26282_, _26281_, _26210_);
  nand _30937_ (_26283_, _26282_, _26201_);
  nand _30938_ (_26284_, _26283_, _26205_);
  nand _30939_ (_26285_, _26284_, _26274_);
  and _30940_ (_26286_, _26285_, _26273_);
  and _30941_ (_26287_, _26286_, _26179_);
  nor _30942_ (_26288_, _26286_, _26179_);
  or _30943_ (_26289_, _26281_, _26210_);
  nand _30944_ (_26290_, _26289_, _26282_);
  nand _30945_ (_26291_, _26290_, _26274_);
  and _30946_ (_26292_, _26271_, _26200_);
  not _30947_ (_26293_, _26292_);
  and _30948_ (_26294_, _26293_, _26291_);
  nand _30949_ (_26295_, _26294_, _26202_);
  nor _30950_ (_26296_, _26295_, _26288_);
  nor _30951_ (_26297_, _26296_, _26287_);
  or _30952_ (_26298_, _26288_, _26287_);
  or _30953_ (_26299_, _26294_, _26202_);
  and _30954_ (_26300_, _26299_, _26295_);
  not _30955_ (_26301_, _26300_);
  nor _30956_ (_26302_, _26301_, _26298_);
  nand _30957_ (_26303_, _26231_, _26278_);
  or _30958_ (_26304_, _26231_, _26278_);
  nand _30959_ (_26305_, _26304_, _26303_);
  nand _30960_ (_26306_, _26305_, _26274_);
  and _30961_ (_26307_, _26271_, _26216_);
  not _30962_ (_26308_, _26307_);
  and _30963_ (_26309_, _26308_, _26306_);
  and _30964_ (_26310_, _26309_, _26208_);
  nor _30965_ (_26311_, _26264_, _26261_);
  or _30966_ (_26312_, _26311_, _26277_);
  and _30967_ (_26313_, _26312_, _26274_);
  and _30968_ (_26314_, _26271_, _26226_);
  nor _30969_ (_26315_, _26314_, _26313_);
  and _30970_ (_26316_, _26315_, _26229_);
  not _30971_ (_26317_, _26316_);
  nor _30972_ (_26318_, _26309_, _26208_);
  or _30973_ (_26319_, _26318_, _26310_);
  nor _30974_ (_26320_, _26319_, _26317_);
  nor _30975_ (_26321_, _26320_, _26310_);
  and _30976_ (_26322_, _26259_, _26244_);
  not _30977_ (_26323_, _26322_);
  and _30978_ (_26324_, _26323_, _26260_);
  or _30979_ (_26325_, _26324_, _26271_);
  or _30980_ (_26326_, _26274_, _26241_);
  and _30981_ (_26327_, _26326_, _26325_);
  nor _30982_ (_26328_, _26327_, _26262_);
  not _30983_ (_26329_, _26328_);
  not _30984_ (_26330_, _26151_);
  or _30985_ (_26331_, _26271_, _26330_);
  nand _30986_ (_26332_, _26331_, _26254_);
  or _30987_ (_26333_, _26331_, _26254_);
  and _30988_ (_26334_, _26333_, _26332_);
  nand _30989_ (_26335_, _26334_, _26245_);
  or _30990_ (_26336_, _26334_, _26245_);
  and _30991_ (_26337_, _26336_, _26335_);
  nor _30992_ (_26338_, _26330_, _26149_);
  not _30993_ (_26339_, _26338_);
  nand _30994_ (_26340_, _26339_, _26337_);
  and _30995_ (_26341_, _26340_, _26335_);
  and _30996_ (_26342_, _26257_, _26255_);
  not _30997_ (_26343_, _26342_);
  and _30998_ (_26344_, _26343_, _26258_);
  or _30999_ (_26345_, _26344_, _26271_);
  or _31000_ (_26346_, _26274_, _26249_);
  and _31001_ (_26347_, _26346_, _26345_);
  nand _31002_ (_26348_, _26347_, _26237_);
  or _31003_ (_26349_, _26347_, _26237_);
  and _31004_ (_26350_, _26349_, _26348_);
  not _31005_ (_26351_, _26350_);
  or _31006_ (_26352_, _26351_, _26341_);
  and _31007_ (_26353_, _26327_, _26262_);
  not _31008_ (_26354_, _26353_);
  and _31009_ (_26355_, _26354_, _26348_);
  nand _31010_ (_26356_, _26355_, _26352_);
  and _31011_ (_26357_, _26356_, _26329_);
  nor _31012_ (_26358_, _26315_, _26229_);
  nor _31013_ (_26359_, _26358_, _26316_);
  not _31014_ (_26360_, _26359_);
  nor _31015_ (_26361_, _26319_, _26360_);
  nand _31016_ (_26362_, _26361_, _26357_);
  nand _31017_ (_26363_, _26362_, _26321_);
  nand _31018_ (_26364_, _26363_, _26302_);
  nand _31019_ (_26365_, _26364_, _26297_);
  and _31020_ (_26366_, _26365_, _26172_);
  nand _31021_ (_26367_, _26366_, _26151_);
  and _31022_ (_26368_, _26367_, _26149_);
  nor _31023_ (_26369_, _26367_, _26149_);
  or _31024_ (_26370_, _26369_, _26368_);
  nand _31025_ (_26371_, _26370_, _23599_);
  nor _31026_ (_26372_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _31027_ (_26373_, _26372_);
  and _31028_ (_26374_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  not _31029_ (_26375_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _31030_ (_26376_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _26375_);
  not _31031_ (_26377_, _26376_);
  or _31032_ (_26378_, _26377_, _23296_);
  not _31033_ (_26379_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _31034_ (_26380_, _26379_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _31035_ (_26381_, _26380_);
  or _31036_ (_26383_, _26381_, _23214_);
  and _31037_ (_26384_, _26383_, _26378_);
  or _31038_ (_26385_, _26380_, _26376_);
  or _31039_ (_26386_, _26385_, _23400_);
  and _31040_ (_26387_, _26386_, _26373_);
  and _31041_ (_26388_, _26387_, _26384_);
  and _31042_ (_26389_, _26372_, _23141_);
  nor _31043_ (_26390_, _26389_, _26388_);
  and _31044_ (_26391_, _26390_, _23359_);
  or _31045_ (_26392_, _26377_, _23404_);
  or _31046_ (_26393_, _26381_, _23263_);
  and _31047_ (_26394_, _26393_, _26392_);
  or _31048_ (_26395_, _26385_, _23418_);
  and _31049_ (_26396_, _26395_, _26373_);
  nand _31050_ (_26397_, _26396_, _26394_);
  or _31051_ (_26398_, _26373_, _23177_);
  and _31052_ (_26399_, _26398_, _26397_);
  and _31053_ (_26400_, _26399_, _23326_);
  nand _31054_ (_26401_, _26400_, _26391_);
  and _31055_ (_26402_, _26399_, _23616_);
  nand _31056_ (_26403_, _26398_, _26397_);
  or _31057_ (_26404_, _26403_, _23612_);
  and _31058_ (_26405_, _26390_, _23326_);
  and _31059_ (_26406_, _26405_, _26404_);
  nand _31060_ (_26407_, _26406_, _26402_);
  nand _31061_ (_26408_, _26407_, _26401_);
  or _31062_ (_26409_, _26389_, _26388_);
  or _31063_ (_26410_, _26409_, _23291_);
  or _31064_ (_26411_, _26403_, _23244_);
  or _31065_ (_26412_, _26411_, _26410_);
  nand _31066_ (_26413_, _26411_, _26410_);
  and _31067_ (_26414_, _26413_, _26412_);
  and _31068_ (_26415_, _26414_, _26408_);
  and _31069_ (_26416_, _26390_, _23525_);
  and _31070_ (_26417_, _26416_, _26402_);
  or _31071_ (_26418_, _26409_, _23522_);
  or _31072_ (_26419_, _26418_, _26411_);
  and _31073_ (_26420_, _26399_, _23208_);
  or _31074_ (_26421_, _26420_, _26416_);
  and _31075_ (_26422_, _26421_, _26419_);
  nand _31076_ (_26423_, _26422_, _26417_);
  or _31077_ (_26424_, _26422_, _26417_);
  and _31078_ (_26425_, _26424_, _26423_);
  nand _31079_ (_26426_, _26425_, _26415_);
  not _31080_ (_26427_, _26418_);
  or _31081_ (_26428_, _26419_, _23171_);
  and _31082_ (_26429_, _26399_, _24028_);
  not _31083_ (_26430_, _26429_);
  nand _31084_ (_26431_, _26430_, _26419_);
  and _31085_ (_26432_, _26431_, _26428_);
  nand _31086_ (_26433_, _26432_, _26427_);
  or _31087_ (_26434_, _26429_, _26427_);
  nand _31088_ (_26435_, _26434_, _26433_);
  or _31089_ (_26436_, _26435_, _26426_);
  or _31090_ (_26437_, _26409_, _23392_);
  nor _31091_ (_26438_, _26437_, _26404_);
  or _31092_ (_26439_, _26400_, _26391_);
  and _31093_ (_26440_, _26439_, _26401_);
  and _31094_ (_26441_, _26440_, _26438_);
  or _31095_ (_26442_, _26406_, _26402_);
  and _31096_ (_26443_, _26442_, _26407_);
  and _31097_ (_26444_, _26443_, _26441_);
  nand _31098_ (_26445_, _26414_, _26408_);
  or _31099_ (_26446_, _26414_, _26408_);
  and _31100_ (_26447_, _26446_, _26445_);
  and _31101_ (_26448_, _26447_, _26444_);
  or _31102_ (_26449_, _26425_, _26415_);
  and _31103_ (_26450_, _26449_, _26426_);
  nand _31104_ (_26451_, _26450_, _26448_);
  not _31105_ (_26452_, _26451_);
  and _31106_ (_26453_, _26426_, _26423_);
  nand _31107_ (_26454_, _26453_, _26435_);
  or _31108_ (_26455_, _26453_, _26435_);
  and _31109_ (_26456_, _26455_, _26454_);
  nand _31110_ (_26457_, _26456_, _26452_);
  nand _31111_ (_26458_, _26457_, _26436_);
  nor _31112_ (_26459_, _26435_, _26423_);
  not _31113_ (_26460_, _26428_);
  and _31114_ (_26461_, _26432_, _26427_);
  or _31115_ (_26462_, _26403_, _23131_);
  or _31116_ (_26463_, _26409_, _23171_);
  or _31117_ (_26464_, _26463_, _26462_);
  nand _31118_ (_26465_, _26463_, _26462_);
  and _31119_ (_26466_, _26465_, _26464_);
  nand _31120_ (_26467_, _26466_, _26461_);
  or _31121_ (_26468_, _26466_, _26461_);
  and _31122_ (_26469_, _26468_, _26467_);
  nand _31123_ (_26470_, _26469_, _26460_);
  or _31124_ (_26471_, _26469_, _26460_);
  and _31125_ (_26472_, _26471_, _26470_);
  nand _31126_ (_26473_, _26472_, _26459_);
  or _31127_ (_26474_, _26472_, _26459_);
  and _31128_ (_26475_, _26474_, _26473_);
  nand _31129_ (_26476_, _26475_, _26458_);
  or _31130_ (_26477_, _26475_, _26458_);
  and _31131_ (_26478_, _26477_, _26476_);
  nand _31132_ (_26479_, _26478_, _26374_);
  or _31133_ (_26480_, _26478_, _26374_);
  and _31134_ (_26481_, _26480_, _26479_);
  and _31135_ (_26482_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or _31136_ (_26483_, _26456_, _26452_);
  and _31137_ (_26484_, _26483_, _26457_);
  nand _31138_ (_26485_, _26484_, _26482_);
  or _31139_ (_26486_, _26484_, _26482_);
  nand _31140_ (_26487_, _26486_, _26485_);
  and _31141_ (_26488_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  or _31142_ (_26489_, _26450_, _26448_);
  and _31143_ (_26490_, _26489_, _26451_);
  nand _31144_ (_26491_, _26490_, _26488_);
  or _31145_ (_26492_, _26490_, _26488_);
  and _31146_ (_26493_, _26492_, _26491_);
  and _31147_ (_26494_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nand _31148_ (_26495_, _26447_, _26444_);
  or _31149_ (_26496_, _26447_, _26444_);
  and _31150_ (_26497_, _26496_, _26495_);
  nand _31151_ (_26498_, _26497_, _26494_);
  and _31152_ (_26499_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nand _31153_ (_26500_, _26443_, _26441_);
  or _31154_ (_26501_, _26443_, _26441_);
  and _31155_ (_26502_, _26501_, _26500_);
  nand _31156_ (_26503_, _26502_, _26499_);
  and _31157_ (_26504_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand _31158_ (_26505_, _26440_, _26438_);
  or _31159_ (_26506_, _26440_, _26438_);
  and _31160_ (_26507_, _26506_, _26505_);
  and _31161_ (_26508_, _26507_, _26504_);
  not _31162_ (_26509_, _26508_);
  or _31163_ (_26510_, _26502_, _26499_);
  nand _31164_ (_26511_, _26510_, _26503_);
  or _31165_ (_26512_, _26511_, _26509_);
  nand _31166_ (_26513_, _26512_, _26503_);
  or _31167_ (_26514_, _26497_, _26494_);
  and _31168_ (_26515_, _26514_, _26498_);
  nand _31169_ (_26516_, _26515_, _26513_);
  nand _31170_ (_26517_, _26516_, _26498_);
  nand _31171_ (_26518_, _26517_, _26493_);
  and _31172_ (_26519_, _26518_, _26491_);
  or _31173_ (_26520_, _26519_, _26487_);
  nand _31174_ (_26521_, _26520_, _26485_);
  nand _31175_ (_26522_, _26521_, _26481_);
  nand _31176_ (_26523_, _26522_, _26479_);
  and _31177_ (_26524_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  nand _31178_ (_26525_, _26476_, _26473_);
  and _31179_ (_26526_, _26390_, _23536_);
  and _31180_ (_26527_, _26526_, _26430_);
  and _31181_ (_26528_, _26470_, _26467_);
  not _31182_ (_26529_, _26528_);
  nand _31183_ (_26530_, _26529_, _26527_);
  or _31184_ (_26531_, _26529_, _26527_);
  and _31185_ (_26532_, _26531_, _26530_);
  nand _31186_ (_26533_, _26532_, _26525_);
  or _31187_ (_26534_, _26532_, _26525_);
  and _31188_ (_26535_, _26534_, _26533_);
  nand _31189_ (_26536_, _26535_, _26524_);
  or _31190_ (_26537_, _26535_, _26524_);
  and _31191_ (_26538_, _26537_, _26536_);
  and _31192_ (_26539_, _26538_, _26523_);
  nor _31193_ (_26540_, _26538_, _26523_);
  nor _31194_ (_26541_, _26540_, _26539_);
  and _31195_ (_26542_, _26541_, _23596_);
  and _31196_ (_26543_, _23521_, _23422_);
  nor _31197_ (_26544_, _26543_, _23492_);
  and _31198_ (_26545_, _26544_, _23087_);
  not _31199_ (_26546_, _26545_);
  and _31200_ (_26547_, _23480_, _26544_);
  and _31201_ (_26548_, _23571_, _23456_);
  not _31202_ (_26549_, _26548_);
  nand _31203_ (_26550_, _23602_, _23359_);
  and _31204_ (_26551_, _23582_, _23536_);
  and _31205_ (_26552_, _23579_, _23567_);
  nor _31206_ (_26553_, _26552_, _26551_);
  or _31207_ (_26554_, _23539_, _23392_);
  and _31208_ (_26555_, _26554_, _23767_);
  and _31209_ (_26556_, _26555_, _23764_);
  and _31210_ (_26557_, _26556_, _26553_);
  and _31211_ (_26558_, _26557_, _26550_);
  nand _31212_ (_26559_, _26558_, _26549_);
  nor _31213_ (_26560_, _26559_, _26547_);
  and _31214_ (_26561_, _26560_, _23760_);
  and _31215_ (_26562_, _26561_, _26546_);
  not _31216_ (_26563_, _26562_);
  nor _31217_ (_26564_, _26563_, _26542_);
  nand _31218_ (_26565_, _26564_, _26371_);
  and _31219_ (_26566_, _24566_, _24542_);
  and _31220_ (_26567_, _24616_, _24613_);
  and _31221_ (_26568_, _25666_, _24446_);
  nor _31222_ (_26569_, _26568_, _26567_);
  nor _31223_ (_26570_, _26569_, _24382_);
  nor _31224_ (_26571_, _26566_, _26570_);
  not _31225_ (_26572_, _24382_);
  and _31226_ (_26573_, _26567_, _26572_);
  not _31227_ (_26574_, _26573_);
  and _31228_ (_26575_, _24593_, _24567_);
  and _31229_ (_26576_, _26575_, _26572_);
  nor _31230_ (_26577_, _26576_, _24628_);
  and _31231_ (_26578_, _26577_, _26574_);
  not _31232_ (_26579_, _24566_);
  nor _31233_ (_26580_, _25630_, _26579_);
  and _31234_ (_26581_, _25667_, _24618_);
  and _31235_ (_26582_, _24554_, _25665_);
  and _31236_ (_26583_, _24606_, _26582_);
  or _31237_ (_26584_, _26583_, _26581_);
  and _31238_ (_26585_, _24440_, _24417_);
  and _31239_ (_26586_, _24538_, _24553_);
  and _31240_ (_26587_, _26586_, _26585_);
  and _31241_ (_26588_, _26587_, _24535_);
  and _31242_ (_26589_, _24538_, _24445_);
  and _31243_ (_26590_, _26589_, _24535_);
  or _31244_ (_26591_, _26590_, _26588_);
  or _31245_ (_26592_, _26591_, _26584_);
  and _31246_ (_26593_, _26592_, _24566_);
  nor _31247_ (_26594_, _26593_, _26580_);
  nand _31248_ (_26595_, _26594_, _26578_);
  and _31249_ (_26596_, _26575_, _24471_);
  nor _31250_ (_26597_, _26596_, _25629_);
  and _31251_ (_26598_, _24606_, _24445_);
  or _31252_ (_26599_, _26598_, _24607_);
  and _31253_ (_26600_, _26589_, _24584_);
  nor _31254_ (_26601_, _26600_, _26599_);
  nand _31255_ (_26602_, _26601_, _26597_);
  nor _31256_ (_26603_, _25620_, _24542_);
  not _31257_ (_26604_, _26603_);
  or _31258_ (_26605_, _26604_, _26584_);
  or _31259_ (_26606_, _26605_, _26602_);
  and _31260_ (_26607_, _26606_, _24566_);
  or _31261_ (_26608_, _26576_, _24569_);
  or _31262_ (_26609_, _26608_, _26607_);
  nor _31263_ (_26610_, _26609_, _26595_);
  and _31264_ (_26611_, _26610_, _26571_);
  or _31265_ (_26612_, _26611_, _26566_);
  and _31266_ (_26613_, _26612_, _26565_);
  and _31267_ (_26614_, _24616_, _24471_);
  and _31268_ (_26615_, _26614_, _25667_);
  and _31269_ (_26616_, _24596_, _24535_);
  or _31270_ (_26618_, _26616_, _26615_);
  and _31271_ (_26619_, _25667_, _24606_);
  and _31272_ (_26620_, _24604_, _24447_);
  and _31273_ (_26621_, _24584_, _24567_);
  or _31274_ (_26622_, _26621_, _26620_);
  or _31275_ (_26623_, _26622_, _26619_);
  or _31276_ (_26624_, _26623_, _26618_);
  and _31277_ (_26625_, _24471_, _24445_);
  and _31278_ (_26626_, _26625_, _24535_);
  or _31279_ (_26627_, _26626_, _24614_);
  or _31280_ (_26628_, _24593_, _24589_);
  and _31281_ (_26629_, _25667_, _26628_);
  or _31282_ (_26630_, _25638_, _24546_);
  and _31283_ (_26631_, _26630_, _25667_);
  or _31284_ (_26632_, _26631_, _26629_);
  or _31285_ (_26633_, _26632_, _26627_);
  not _31286_ (_26634_, _26597_);
  and _31287_ (_26635_, _24613_, _24536_);
  and _31288_ (_26636_, _25633_, _24612_);
  or _31289_ (_26637_, _26636_, _26635_);
  or _31290_ (_26638_, _26637_, _26634_);
  or _31291_ (_26639_, _26638_, _26633_);
  or _31292_ (_26640_, _26639_, _26624_);
  and _31293_ (_26641_, _24606_, _24567_);
  or _31294_ (_26643_, _26581_, _26641_);
  and _31295_ (_26644_, _24613_, _24541_);
  and _31296_ (_26645_, _24616_, _24538_);
  and _31297_ (_26646_, _26645_, _25667_);
  or _31298_ (_26647_, _26646_, _26644_);
  or _31299_ (_26648_, _26647_, _26643_);
  and _31300_ (_26650_, _24588_, _24471_);
  and _31301_ (_26651_, _25667_, _26650_);
  and _31302_ (_26652_, _24567_, _24536_);
  or _31303_ (_26653_, _26652_, _26651_);
  and _31304_ (_26654_, _26650_, _24447_);
  or _31305_ (_26655_, _25621_, _24606_);
  and _31306_ (_26656_, _26655_, _24613_);
  or _31307_ (_26657_, _26656_, _26654_);
  or _31308_ (_26658_, _26657_, _26653_);
  or _31309_ (_26659_, _26658_, _26648_);
  and _31310_ (_26660_, _24613_, _24552_);
  and _31311_ (_26661_, _24589_, _24447_);
  or _31312_ (_26662_, _26661_, _26660_);
  and _31313_ (_26663_, _25667_, _24604_);
  and _31314_ (_26665_, _25621_, _25667_);
  or _31315_ (_26666_, _26665_, _26663_);
  and _31316_ (_26668_, _24613_, _24546_);
  or _31317_ (_26669_, _25668_, _26668_);
  or _31318_ (_26670_, _26669_, _26666_);
  or _31319_ (_26671_, _26670_, _26662_);
  or _31320_ (_26672_, _26671_, _26659_);
  or _31321_ (_26673_, _26672_, _26640_);
  nand _31322_ (_26674_, _26673_, _26572_);
  nor _31323_ (_26675_, _24628_, _24569_);
  nand _31324_ (_26676_, _26675_, _26674_);
  nand _31325_ (_26677_, _26676_, _22766_);
  and _31326_ (_26678_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _31327_ (_26679_, _26678_);
  and _31328_ (_26680_, _26679_, _26677_);
  nor _31329_ (_26681_, _26680_, _24634_);
  and _31330_ (_26682_, _26681_, _24576_);
  and _31331_ (_26683_, _24067_, _23002_);
  and _31332_ (_26684_, _26683_, _24077_);
  not _31333_ (_26685_, _26684_);
  nor _31334_ (_26686_, _26685_, _23702_);
  and _31335_ (_26687_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _31336_ (_26688_, _26684_, _23738_);
  nor _31337_ (_26689_, _26688_, _26687_);
  and _31338_ (_26691_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _31339_ (_26692_, _26684_, _23816_);
  or _31340_ (_26693_, _26692_, _26691_);
  nand _31341_ (_26694_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nand _31342_ (_26695_, _26684_, _23892_);
  and _31343_ (_26696_, _26695_, _26694_);
  or _31344_ (_26697_, _26684_, _23012_);
  nand _31345_ (_26698_, _26684_, _24685_);
  and _31346_ (_26699_, _26698_, _26697_);
  and _31347_ (_26700_, _26699_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _31348_ (_26701_, _26700_, _26696_);
  not _31349_ (_26702_, _26701_);
  nor _31350_ (_26703_, _26702_, _26693_);
  and _31351_ (_26704_, _26703_, _26689_);
  and _31352_ (_26705_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _31353_ (_26707_, _26684_, _23642_);
  nor _31354_ (_26708_, _26707_, _26705_);
  and _31355_ (_26709_, _26708_, _26704_);
  and _31356_ (_26710_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _31357_ (_26711_, _26684_, _23939_);
  nor _31358_ (_26712_, _26711_, _26710_);
  and _31359_ (_26713_, _26712_, _26709_);
  and _31360_ (_26714_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and _31361_ (_26715_, _26684_, _24043_);
  nor _31362_ (_26716_, _26715_, _26714_);
  and _31363_ (_26717_, _26716_, _26713_);
  and _31364_ (_26718_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and _31365_ (_26719_, _26718_, _26717_);
  nor _31366_ (_26721_, _26718_, _26717_);
  or _31367_ (_26722_, _26721_, _22920_);
  or _31368_ (_26723_, _26722_, _26719_);
  and _31369_ (_26724_, _26723_, _22924_);
  nor _31370_ (_26725_, _26724_, _26684_);
  or _31371_ (_26727_, _26725_, _26686_);
  nand _31372_ (_26728_, _26727_, _26682_);
  not _31373_ (_26729_, _24634_);
  and _31374_ (_26730_, _26680_, _26729_);
  and _31375_ (_26732_, _26730_, _24576_);
  nand _31376_ (_26733_, _25956_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nand _31377_ (_26734_, _25948_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _31378_ (_26735_, _26734_, _26733_);
  nand _31379_ (_26736_, _25945_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand _31380_ (_26737_, _25937_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _31381_ (_26738_, _26737_, _26736_);
  and _31382_ (_26739_, _26738_, _26735_);
  nand _31383_ (_26740_, _25954_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nand _31384_ (_26741_, _25940_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _31385_ (_26742_, _26741_, _26740_);
  nand _31386_ (_26743_, _25961_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nand _31387_ (_26744_, _25959_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _31388_ (_26745_, _26744_, _26743_);
  and _31389_ (_26746_, _26745_, _26742_);
  and _31390_ (_26747_, _26746_, _26739_);
  nor _31391_ (_26749_, _26747_, _25935_);
  not _31392_ (_26750_, _23702_);
  and _31393_ (_26751_, _25935_, _26750_);
  or _31394_ (_26752_, _26751_, _26749_);
  nand _31395_ (_26753_, _26752_, _26732_);
  nor _31396_ (_26754_, _26680_, _26729_);
  nor _31397_ (_26755_, _22768_, _23104_);
  and _31398_ (_26756_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _31399_ (_26757_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _31400_ (_26758_, _26757_, _26756_);
  and _31401_ (_26759_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _31402_ (_26760_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _31403_ (_26761_, _26760_, _26759_);
  and _31404_ (_26762_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _31405_ (_26763_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _31406_ (_26765_, _26763_, _26762_);
  and _31407_ (_26766_, _26765_, _26761_);
  and _31408_ (_26767_, _26766_, _26758_);
  nor _31409_ (_26768_, _26767_, _25729_);
  nor _31410_ (_26770_, _26768_, _26755_);
  not _31411_ (_26772_, _26770_);
  nand _31412_ (_26773_, _26772_, _26754_);
  and _31413_ (_26775_, _26773_, _24576_);
  and _31414_ (_26776_, _26775_, _26753_);
  nand _31415_ (_26777_, _26776_, _26728_);
  and _31416_ (_26778_, _26777_, _22943_);
  nor _31417_ (_26779_, _26777_, _22943_);
  nor _31418_ (_26781_, _26779_, _26778_);
  not _31419_ (_26782_, _26682_);
  nor _31420_ (_26783_, _26716_, _26713_);
  nor _31421_ (_26784_, _26783_, _26717_);
  nor _31422_ (_26785_, _26784_, _22920_);
  nor _31423_ (_26786_, _26785_, _23025_);
  nor _31424_ (_26787_, _26786_, _26684_);
  nor _31425_ (_26788_, _26787_, _26715_);
  nor _31426_ (_26789_, _26788_, _26782_);
  not _31427_ (_26790_, _26789_);
  not _31428_ (_26791_, _26732_);
  nor _31429_ (_26792_, _26088_, _26791_);
  not _31430_ (_26793_, _26792_);
  and _31431_ (_26794_, _24634_, _24577_);
  and _31432_ (_26795_, _26681_, _24577_);
  nor _31433_ (_26796_, _26795_, _26794_);
  nor _31434_ (_26797_, _22768_, _23154_);
  and _31435_ (_26798_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _31436_ (_26799_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _31437_ (_26800_, _26799_, _26798_);
  and _31438_ (_26801_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _31439_ (_26802_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _31440_ (_26803_, _26802_, _26801_);
  and _31441_ (_26804_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _31442_ (_26806_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _31443_ (_26807_, _26806_, _26804_);
  and _31444_ (_26808_, _26807_, _26803_);
  and _31445_ (_26809_, _26808_, _26800_);
  nor _31446_ (_26810_, _26809_, _25729_);
  nor _31447_ (_26811_, _26810_, _26797_);
  not _31448_ (_26812_, _26811_);
  and _31449_ (_26813_, _26812_, _26754_);
  not _31450_ (_26814_, _26813_);
  and _31451_ (_26815_, _26814_, _26796_);
  and _31452_ (_26816_, _26815_, _26793_);
  and _31453_ (_26817_, _26816_, _26790_);
  nor _31454_ (_26818_, _26817_, _23034_);
  and _31455_ (_26819_, _26817_, _23034_);
  nor _31456_ (_26820_, _26819_, _26818_);
  nor _31457_ (_26821_, _26712_, _26709_);
  nor _31458_ (_26822_, _26821_, _26713_);
  nor _31459_ (_26823_, _26822_, _22920_);
  nor _31460_ (_26824_, _26823_, _23044_);
  nor _31461_ (_26825_, _26824_, _26684_);
  nor _31462_ (_26826_, _26825_, _26711_);
  nor _31463_ (_26827_, _26826_, _26782_);
  not _31464_ (_26829_, _26827_);
  nor _31465_ (_26830_, _26065_, _26791_);
  not _31466_ (_26831_, _26830_);
  and _31467_ (_26832_, _26754_, _24576_);
  nor _31468_ (_26833_, _22768_, _23191_);
  and _31469_ (_26835_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _31470_ (_26836_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _31471_ (_26837_, _26836_, _26835_);
  and _31472_ (_26838_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _31473_ (_26839_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _31474_ (_26840_, _26839_, _26838_);
  and _31475_ (_26841_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _31476_ (_00001_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _31477_ (_00002_, _00001_, _26841_);
  and _31478_ (_00003_, _00002_, _26840_);
  and _31479_ (_00004_, _00003_, _26837_);
  nor _31480_ (_00005_, _00004_, _25729_);
  nor _31481_ (_00006_, _00005_, _26833_);
  not _31482_ (_00007_, _00006_);
  and _31483_ (_00008_, _00007_, _26832_);
  not _31484_ (_00009_, _00008_);
  and _31485_ (_00010_, _26794_, _26680_);
  nor _31486_ (_00011_, _26795_, _00010_);
  and _31487_ (_00012_, _00011_, _00009_);
  and _31488_ (_00013_, _00012_, _26831_);
  and _31489_ (_00014_, _00013_, _26829_);
  nor _31490_ (_00015_, _00014_, _23052_);
  and _31491_ (_00016_, _00014_, _23052_);
  nor _31492_ (_00017_, _00016_, _00015_);
  nor _31493_ (_00018_, _26024_, _26791_);
  not _31494_ (_00019_, _26145_);
  and _31495_ (_00020_, _26832_, _00019_);
  nor _31496_ (_00021_, _00020_, _00018_);
  not _31497_ (_00022_, _26689_);
  or _31498_ (_00023_, _26702_, _26693_);
  and _31499_ (_00024_, _00023_, _00022_);
  nor _31500_ (_00025_, _00024_, _26704_);
  nor _31501_ (_00026_, _00025_, _22920_);
  nor _31502_ (_00027_, _00026_, _22990_);
  nor _31503_ (_00028_, _00027_, _26684_);
  nor _31504_ (_00029_, _00028_, _26688_);
  not _31505_ (_00030_, _00029_);
  and _31506_ (_00031_, _00030_, _26682_);
  and _31507_ (_00032_, _24634_, _24576_);
  and _31508_ (_00033_, _00032_, _26680_);
  not _31509_ (_00034_, _00033_);
  nor _31510_ (_00035_, _00034_, _25780_);
  nor _31511_ (_00036_, _00035_, _00031_);
  and _31512_ (_00037_, _00036_, _00021_);
  nor _31513_ (_00038_, _00037_, _23002_);
  and _31514_ (_00039_, _00037_, _23002_);
  nor _31515_ (_00040_, _00039_, _00038_);
  nor _31516_ (_00041_, _26708_, _26704_);
  nor _31517_ (_00042_, _00041_, _26709_);
  nor _31518_ (_00043_, _00042_, _22920_);
  nor _31519_ (_00044_, _00043_, _22954_);
  nor _31520_ (_00045_, _00044_, _26684_);
  nor _31521_ (_00046_, _00045_, _26707_);
  not _31522_ (_00047_, _00046_);
  and _31523_ (_00048_, _00047_, _26682_);
  not _31524_ (_00049_, _00048_);
  nor _31525_ (_00050_, _26043_, _26791_);
  not _31526_ (_00051_, _25731_);
  and _31527_ (_00052_, _26754_, _00051_);
  not _31528_ (_00053_, _00052_);
  and _31529_ (_00054_, _00033_, _25953_);
  nor _31530_ (_00055_, _00054_, _26794_);
  nand _31531_ (_00056_, _00055_, _00053_);
  nor _31532_ (_00057_, _00056_, _00050_);
  and _31533_ (_00058_, _00057_, _00049_);
  nor _31534_ (_00059_, _00058_, _22970_);
  and _31535_ (_00060_, _00058_, _22970_);
  nor _31536_ (_00061_, _00060_, _00059_);
  or _31537_ (_00062_, _00061_, _00040_);
  or _31538_ (_00063_, _00062_, _00017_);
  or _31539_ (_00064_, _00063_, _26820_);
  nor _31540_ (_00065_, _00064_, _26781_);
  nor _31541_ (_00066_, _25987_, _26791_);
  nor _31542_ (_00067_, _24634_, _24576_);
  and _31543_ (_00068_, _00032_, _24417_);
  or _31544_ (_00069_, _00068_, _00067_);
  and _31545_ (_00070_, _00069_, _26680_);
  nor _31546_ (_00071_, _26700_, _26696_);
  nor _31547_ (_00072_, _00071_, _26701_);
  nor _31548_ (_00073_, _00072_, _22920_);
  nor _31549_ (_00074_, _00073_, _22975_);
  nor _31550_ (_00075_, _00074_, _26684_);
  not _31551_ (_00076_, _00075_);
  and _31552_ (_00077_, _00076_, _26695_);
  not _31553_ (_00078_, _00077_);
  and _31554_ (_00079_, _00078_, _26682_);
  nor _31555_ (_00080_, _22768_, _23343_);
  and _31556_ (_00081_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _31557_ (_00082_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _31558_ (_00083_, _00082_, _00081_);
  and _31559_ (_00084_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _31560_ (_00085_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _31561_ (_00086_, _00085_, _00084_);
  and _31562_ (_00087_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _31563_ (_00088_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _31564_ (_00089_, _00088_, _00087_);
  and _31565_ (_00091_, _00089_, _00086_);
  and _31566_ (_00092_, _00091_, _00083_);
  nor _31567_ (_00093_, _00092_, _25729_);
  nor _31568_ (_00094_, _00093_, _00080_);
  not _31569_ (_00095_, _00094_);
  and _31570_ (_00096_, _00095_, _26832_);
  or _31571_ (_00097_, _00096_, _00079_);
  or _31572_ (_00098_, _00097_, _00070_);
  nor _31573_ (_00099_, _00098_, _00066_);
  and _31574_ (_00100_, _00099_, _24289_);
  nor _31575_ (_00101_, _00099_, _24289_);
  or _31576_ (_00102_, _00101_, _00100_);
  not _31577_ (_00103_, _00102_);
  nor _31578_ (_00104_, _25968_, _26791_);
  not _31579_ (_00105_, _00104_);
  nor _31580_ (_00106_, _26699_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor _31581_ (_00107_, _00106_, _26700_);
  nor _31582_ (_00108_, _00107_, _22920_);
  nor _31583_ (_00109_, _00108_, _23014_);
  nor _31584_ (_00110_, _00109_, _26684_);
  not _31585_ (_00111_, _00110_);
  and _31586_ (_00112_, _00111_, _26698_);
  not _31587_ (_00113_, _00112_);
  and _31588_ (_00114_, _00113_, _26682_);
  nand _31589_ (_00115_, _00033_, _24408_);
  nor _31590_ (_00116_, _22768_, _23375_);
  and _31591_ (_00117_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _31592_ (_00118_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _31593_ (_00119_, _00118_, _00117_);
  and _31594_ (_00120_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _31595_ (_00121_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _31596_ (_00122_, _00121_, _00120_);
  and _31597_ (_00123_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _31598_ (_00124_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _31599_ (_00125_, _00124_, _00123_);
  and _31600_ (_00126_, _00125_, _00122_);
  and _31601_ (_00127_, _00126_, _00119_);
  nor _31602_ (_00128_, _00127_, _25729_);
  nor _31603_ (_00129_, _00128_, _00116_);
  not _31604_ (_00130_, _00129_);
  nand _31605_ (_00131_, _00130_, _26832_);
  nand _31606_ (_00132_, _00131_, _00115_);
  nor _31607_ (_00133_, _00132_, _00114_);
  and _31608_ (_00134_, _00133_, _00105_);
  nor _31609_ (_00135_, _00134_, _23018_);
  and _31610_ (_00136_, _00134_, _23018_);
  nor _31611_ (_00137_, _00136_, _00135_);
  not _31612_ (_00138_, _00137_);
  nor _31613_ (_00139_, _26006_, _26791_);
  not _31614_ (_00140_, _00139_);
  and _31615_ (_00141_, _00033_, _24440_);
  and _31616_ (_00142_, _26702_, _26693_);
  nor _31617_ (_00143_, _00142_, _26703_);
  nor _31618_ (_00144_, _00143_, _22920_);
  nor _31619_ (_00145_, _00144_, _23057_);
  nor _31620_ (_00146_, _00145_, _26684_);
  nor _31621_ (_00147_, _00146_, _26692_);
  not _31622_ (_00148_, _00147_);
  and _31623_ (_00149_, _00148_, _26682_);
  nor _31624_ (_00150_, _22768_, _23322_);
  and _31625_ (_00151_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _31626_ (_00152_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _31627_ (_00153_, _00152_, _00151_);
  and _31628_ (_00154_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _31629_ (_00155_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _31630_ (_00156_, _00155_, _00154_);
  and _31631_ (_00157_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _31632_ (_00158_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _31633_ (_00159_, _00158_, _00157_);
  and _31634_ (_00160_, _00159_, _00156_);
  and _31635_ (_00161_, _00160_, _00153_);
  nor _31636_ (_00162_, _00161_, _25729_);
  nor _31637_ (_00163_, _00162_, _00150_);
  not _31638_ (_00164_, _00163_);
  and _31639_ (_00165_, _00164_, _26832_);
  or _31640_ (_00166_, _00165_, _00149_);
  nor _31641_ (_00167_, _00166_, _00141_);
  and _31642_ (_00168_, _00167_, _00140_);
  nor _31643_ (_00169_, _00168_, _23065_);
  and _31644_ (_00170_, _00168_, _23065_);
  nor _31645_ (_00171_, _00170_, _00169_);
  nor _31646_ (_00172_, _00171_, _25181_);
  and _31647_ (_00173_, _00172_, _00138_);
  and _31648_ (_00174_, _00173_, _00103_);
  and _31649_ (_00175_, _00174_, _00065_);
  and _31650_ (_00176_, _22943_, _22948_);
  and _31651_ (_00177_, _00176_, _00175_);
  not _31652_ (_00178_, _00177_);
  nor _31653_ (_00179_, _26597_, _26579_);
  nor _31654_ (_00180_, _26597_, _24382_);
  nor _31655_ (_00181_, _00180_, _00179_);
  not _31656_ (_00182_, _00181_);
  nor _31657_ (_00183_, _24654_, _24070_);
  and _31658_ (_00184_, _00183_, _00065_);
  and _31659_ (_00185_, _00184_, _00182_);
  and _31660_ (_00186_, _23471_, _23483_);
  nor _31661_ (_00187_, _23471_, _23483_);
  nor _31662_ (_00188_, _00187_, _00186_);
  not _31663_ (_00189_, _00188_);
  nor _31664_ (_00190_, _23469_, _23259_);
  nor _31665_ (_00191_, _00190_, _23470_);
  nor _31666_ (_00192_, _23468_, _23262_);
  nor _31667_ (_00193_, _00192_, _23469_);
  nor _31668_ (_00194_, _23467_, _23266_);
  and _31669_ (_00195_, _23467_, _23266_);
  nor _31670_ (_00196_, _00195_, _00194_);
  not _31671_ (_00197_, _00196_);
  and _31672_ (_00198_, _23460_, _23411_);
  nor _31673_ (_00199_, _00198_, _23461_);
  nor _31674_ (_00201_, _26544_, _23416_);
  nor _31675_ (_00202_, _23458_, _23414_);
  nor _31676_ (_00204_, _00202_, _23459_);
  and _31677_ (_00205_, _00204_, _00201_);
  and _31678_ (_00207_, _00205_, _00199_);
  not _31679_ (_00208_, _24569_);
  and _31680_ (_00209_, _00181_, _00208_);
  and _31681_ (_00210_, _00209_, _00207_);
  and _31682_ (_00211_, _00210_, _00197_);
  and _31683_ (_00212_, _00211_, _00193_);
  and _31684_ (_00213_, _00212_, _00191_);
  and _31685_ (_00214_, _00213_, _00189_);
  nor _31686_ (_00215_, _00181_, _23561_);
  not _31687_ (_00216_, _00215_);
  and _31688_ (_00217_, _00181_, _24534_);
  nor _31689_ (_00218_, _00217_, _00208_);
  and _31690_ (_00219_, _00218_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _31691_ (_00220_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _31692_ (_00221_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _31693_ (_00222_, _00221_, _00220_);
  nor _31694_ (_00223_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _31695_ (_00224_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _31696_ (_00225_, _00224_, _00223_);
  and _31697_ (_00226_, _00225_, _00222_);
  and _31698_ (_00227_, _00226_, _24630_);
  nor _31699_ (_00228_, _00227_, _00219_);
  and _31700_ (_00229_, _00228_, _00216_);
  not _31701_ (_00230_, _00229_);
  nor _31702_ (_00231_, _00230_, _00214_);
  nor _31703_ (_00232_, _26600_, _26584_);
  not _31704_ (_00233_, _24567_);
  and _31705_ (_00234_, _24593_, _24538_);
  or _31706_ (_00235_, _24589_, _24541_);
  nor _31707_ (_00236_, _00235_, _00234_);
  nor _31708_ (_00237_, _00236_, _00233_);
  nor _31709_ (_00238_, _00237_, _26591_);
  and _31710_ (_00239_, _00238_, _00232_);
  not _31711_ (_00240_, _00239_);
  and _31712_ (_00241_, _00240_, _00231_);
  and _31713_ (_00242_, _26603_, _24615_);
  not _31714_ (_00243_, _00242_);
  nor _31715_ (_00244_, _00243_, _00241_);
  nand _31716_ (_00245_, _25629_, _24544_);
  and _31717_ (_00246_, _24568_, _24471_);
  nor _31718_ (_00247_, _00246_, _26596_);
  and _31719_ (_00248_, _00247_, _00245_);
  or _31720_ (_00249_, _00248_, _00231_);
  and _31721_ (_00250_, _00249_, _00244_);
  nor _31722_ (_00251_, _24628_, _24566_);
  nor _31723_ (_00252_, _00251_, _00250_);
  nor _31724_ (_00253_, _00252_, _26570_);
  not _31725_ (_00254_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _31726_ (_00255_, _22766_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _31727_ (_00256_, _00255_, _00254_);
  not _31728_ (_00257_, _00256_);
  not _31729_ (_00258_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _31730_ (_00259_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _22766_);
  and _31731_ (_00260_, _00259_, _00258_);
  and _31732_ (_00261_, _24733_, _23662_);
  and _31733_ (_00262_, _00261_, _25770_);
  nor _31734_ (_00263_, _00262_, _00260_);
  and _31735_ (_00264_, _00263_, _00257_);
  nor _31736_ (_00265_, _23052_, _23034_);
  and _31737_ (_00266_, _00265_, _24645_);
  and _31738_ (_00267_, _00266_, _25259_);
  not _31739_ (_00268_, _00267_);
  and _31740_ (_00270_, _00268_, _00264_);
  not _31741_ (_00271_, _00270_);
  and _31742_ (_00272_, _00271_, _24630_);
  nor _31743_ (_00273_, _23053_, _23034_);
  and _31744_ (_00274_, _00273_, _24645_);
  and _31745_ (_00276_, _00274_, _25163_);
  nor _31746_ (_00277_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not _31747_ (_00278_, _00277_);
  nor _31748_ (_00280_, _00278_, _00276_);
  and _31749_ (_00281_, _00280_, _25774_);
  not _31750_ (_00282_, _00281_);
  and _31751_ (_00283_, _00282_, _00218_);
  nor _31752_ (_00284_, _00283_, _00272_);
  not _31753_ (_00285_, _00284_);
  nor _31754_ (_00286_, _00285_, _00253_);
  not _31755_ (_00287_, _00286_);
  nor _31756_ (_00288_, _00287_, _00185_);
  and _31757_ (_00289_, _00288_, _00178_);
  and _31758_ (_00290_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  not _31759_ (_00291_, _25566_);
  and _31760_ (_00292_, _26573_, _00291_);
  and _31761_ (_00293_, _24567_, _26572_);
  and _31762_ (_00294_, _00293_, _24593_);
  nor _31763_ (_00295_, _26591_, _24568_);
  and _31764_ (_00297_, _00295_, _26603_);
  and _31765_ (_00298_, _00297_, _25630_);
  and _31766_ (_00300_, _00298_, _00232_);
  nor _31767_ (_00301_, _00300_, _26579_);
  nor _31768_ (_00302_, _00301_, _00294_);
  not _31769_ (_00303_, _26571_);
  and _31770_ (_00304_, _26594_, _26578_);
  and _31771_ (_00305_, _00304_, _00303_);
  and _31772_ (_00306_, _00305_, _00302_);
  and _31773_ (_00307_, _00306_, _00130_);
  or _31774_ (_00308_, _00307_, _00292_);
  or _31775_ (_00310_, _00308_, _00290_);
  and _31776_ (_00311_, _26595_, _00291_);
  and _31777_ (_00312_, _00304_, _00130_);
  or _31778_ (_00313_, _00312_, _00311_);
  nor _31779_ (_00314_, _00313_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _31780_ (_00315_, _00313_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _31781_ (_00316_, _00315_, _00314_);
  nor _31782_ (_00317_, _00305_, _00302_);
  and _31783_ (_00318_, _00317_, _00316_);
  nor _31784_ (_00319_, _00318_, _00310_);
  nand _31785_ (_00320_, _00319_, _00289_);
  or _31786_ (_00321_, _00320_, _26613_);
  or _31787_ (_00322_, _00289_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _31788_ (_00323_, _00322_, _22762_);
  and _31789_ (_26890_[0], _00323_, _00321_);
  not _31790_ (_00324_, _26536_);
  nor _31791_ (_00325_, _26539_, _00324_);
  and _31792_ (_00326_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  and _31793_ (_00327_, _26530_, _26464_);
  nand _31794_ (_00328_, _00327_, _26533_);
  nand _31795_ (_00329_, _00328_, _00326_);
  or _31796_ (_00330_, _00328_, _00326_);
  nand _31797_ (_00331_, _00330_, _00329_);
  or _31798_ (_00332_, _00331_, _00325_);
  nand _31799_ (_00333_, _00331_, _00325_);
  and _31800_ (_00334_, _00333_, _00332_);
  nand _31801_ (_00335_, _00334_, _23596_);
  nand _31802_ (_00336_, _26365_, _26172_);
  or _31803_ (_00337_, _26339_, _26337_);
  and _31804_ (_00338_, _00337_, _26340_);
  or _31805_ (_00339_, _00338_, _00336_);
  or _31806_ (_00340_, _26366_, _26334_);
  and _31807_ (_00341_, _00340_, _00339_);
  nand _31808_ (_00342_, _00341_, _23599_);
  nor _31809_ (_00343_, _23419_, _23367_);
  or _31810_ (_00344_, _00343_, _23485_);
  and _31811_ (_00345_, _00344_, _23492_);
  nor _31812_ (_00346_, _00344_, _23492_);
  or _31813_ (_00347_, _00346_, _00345_);
  and _31814_ (_00348_, _00347_, _23480_);
  nor _31815_ (_00349_, _23457_, _23417_);
  nor _31816_ (_00350_, _00349_, _23458_);
  nor _31817_ (_00351_, _00350_, _23088_);
  nor _31818_ (_00352_, _00351_, _00348_);
  nor _31819_ (_00353_, _23530_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _31820_ (_00354_, _00353_, _23359_);
  nor _31821_ (_00355_, _00353_, _23359_);
  nor _31822_ (_00356_, _00355_, _00354_);
  nor _31823_ (_00357_, _00356_, _23539_);
  not _31824_ (_00358_, _00357_);
  not _31825_ (_00359_, _23604_);
  nor _31826_ (_00360_, _00359_, _23392_);
  not _31827_ (_00361_, _00360_);
  nand _31828_ (_00362_, _23602_, _23326_);
  and _31829_ (_00363_, _23579_, _23359_);
  not _31830_ (_00364_, _00363_);
  and _31831_ (_00365_, _00364_, _00362_);
  and _31832_ (_00366_, _00365_, _00361_);
  and _31833_ (_00367_, _00366_, _23889_);
  and _31834_ (_00368_, _00367_, _00358_);
  and _31835_ (_00369_, _00368_, _23878_);
  and _31836_ (_00370_, _00369_, _00352_);
  and _31837_ (_00371_, _00370_, _00342_);
  and _31838_ (_00372_, _00371_, _00335_);
  not _31839_ (_00373_, _00372_);
  and _31840_ (_00374_, _00373_, _26612_);
  nor _31841_ (_00375_, _22768_, _23341_);
  and _31842_ (_00376_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and _31843_ (_00377_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _31844_ (_00378_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _31845_ (_00379_, _00378_, _00377_);
  and _31846_ (_00380_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _31847_ (_00381_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or _31848_ (_00382_, _00381_, _00380_);
  or _31849_ (_00383_, _00382_, _00379_);
  and _31850_ (_00384_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _31851_ (_00386_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _31852_ (_00387_, _00386_, _00384_);
  or _31853_ (_00388_, _00387_, _00383_);
  and _31854_ (_00389_, _00388_, _23839_);
  or _31855_ (_00390_, _00389_, _00376_);
  and _31856_ (_00391_, _00390_, _22768_);
  nor _31857_ (_00392_, _00391_, _00375_);
  or _31858_ (_00393_, _00392_, _00304_);
  or _31859_ (_00394_, _26595_, _00094_);
  and _31860_ (_00395_, _00394_, _00393_);
  or _31861_ (_00396_, _00395_, _23336_);
  nand _31862_ (_00397_, _00395_, _23336_);
  and _31863_ (_00398_, _00397_, _00396_);
  and _31864_ (_00399_, _00398_, _00315_);
  not _31865_ (_00400_, _00305_);
  and _31866_ (_00401_, _00400_, _26609_);
  or _31867_ (_00402_, _00398_, _00315_);
  nand _31868_ (_00403_, _00402_, _00401_);
  or _31869_ (_00404_, _00403_, _00399_);
  and _31870_ (_00405_, _26610_, _00303_);
  and _31871_ (_00406_, _00405_, _00095_);
  nor _31872_ (_00407_, _00392_, _26574_);
  and _31873_ (_00408_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _31874_ (_00409_, _00408_, _00407_);
  nor _31875_ (_00410_, _00409_, _00406_);
  and _31876_ (_00411_, _00410_, _00404_);
  nand _31877_ (_00412_, _00411_, _00289_);
  or _31878_ (_00413_, _00412_, _00374_);
  or _31879_ (_00414_, _00289_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _31880_ (_00415_, _00414_, _22762_);
  and _31881_ (_26890_[1], _00415_, _00413_);
  not _31882_ (_00416_, _00289_);
  not _31883_ (_00417_, _26352_);
  and _31884_ (_00418_, _26351_, _26341_);
  nor _31885_ (_00419_, _00418_, _00417_);
  or _31886_ (_00420_, _00419_, _00336_);
  or _31887_ (_00421_, _26366_, _26347_);
  and _31888_ (_00422_, _00421_, _00420_);
  nand _31889_ (_00423_, _00422_, _23599_);
  and _31890_ (_00424_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  nand _31891_ (_00425_, _00332_, _00329_);
  nand _31892_ (_00426_, _00425_, _00424_);
  or _31893_ (_00427_, _00425_, _00424_);
  and _31894_ (_00428_, _00427_, _00426_);
  nand _31895_ (_00429_, _00428_, _23596_);
  nor _31896_ (_00430_, _00204_, _23088_);
  or _31897_ (_00431_, _23603_, _23291_);
  and _31898_ (_00432_, _23579_, _23326_);
  not _31899_ (_00433_, _00432_);
  nand _31900_ (_00434_, _23604_, _23359_);
  and _31901_ (_00435_, _00434_, _00433_);
  and _31902_ (_00436_, _00435_, _00431_);
  and _31903_ (_00437_, _00436_, _23811_);
  not _31904_ (_00438_, _00437_);
  nor _31905_ (_00439_, _00438_, _00430_);
  nor _31906_ (_00440_, _23495_, _23493_);
  nor _31907_ (_00441_, _00440_, _23481_);
  and _31908_ (_00442_, _00441_, _23497_);
  and _31909_ (_00443_, _23529_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _31910_ (_00444_, _00355_, _23610_);
  nor _31911_ (_00445_, _00444_, _00443_);
  nor _31912_ (_00446_, _00445_, _23539_);
  nor _31913_ (_00447_, _00446_, _00442_);
  and _31914_ (_00448_, _00447_, _00439_);
  and _31915_ (_00449_, _00448_, _23803_);
  and _31916_ (_00450_, _00449_, _00429_);
  nand _31917_ (_00451_, _00450_, _00423_);
  and _31918_ (_00452_, _00451_, _26612_);
  and _31919_ (_00453_, _00405_, _00164_);
  nor _31920_ (_00454_, _22768_, _23302_);
  and _31921_ (_00455_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and _31922_ (_00456_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _31923_ (_00457_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or _31924_ (_00458_, _00457_, _00456_);
  and _31925_ (_00459_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _31926_ (_00460_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or _31927_ (_00461_, _00460_, _00459_);
  or _31928_ (_00462_, _00461_, _00458_);
  and _31929_ (_00463_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _31930_ (_00464_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _31931_ (_00465_, _00464_, _00463_);
  or _31932_ (_00466_, _00465_, _00462_);
  and _31933_ (_00467_, _00466_, _23839_);
  or _31934_ (_00468_, _00467_, _00455_);
  and _31935_ (_00469_, _00468_, _22768_);
  nor _31936_ (_00470_, _00469_, _00454_);
  not _31937_ (_00471_, _00470_);
  and _31938_ (_00472_, _00471_, _26573_);
  and _31939_ (_00473_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _31940_ (_00474_, _00473_, _00472_);
  or _31941_ (_00475_, _00474_, _00453_);
  not _31942_ (_00476_, _00396_);
  or _31943_ (_00477_, _00399_, _00476_);
  and _31944_ (_00478_, _00471_, _26595_);
  and _31945_ (_00479_, _00304_, _00164_);
  nor _31946_ (_00480_, _00479_, _00478_);
  nor _31947_ (_00481_, _00480_, _23307_);
  and _31948_ (_00482_, _00480_, _23307_);
  nor _31949_ (_00483_, _00482_, _00481_);
  or _31950_ (_00484_, _00483_, _00477_);
  and _31951_ (_00485_, _00483_, _00477_);
  not _31952_ (_00486_, _00485_);
  and _31953_ (_00487_, _00486_, _00317_);
  and _31954_ (_00488_, _00487_, _00484_);
  or _31955_ (_00489_, _00488_, _00475_);
  or _31956_ (_00490_, _00489_, _00452_);
  or _31957_ (_00491_, _00490_, _00416_);
  not _31958_ (_00492_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _31959_ (_00493_, _23953_, _00492_);
  and _31960_ (_00494_, _23953_, _00492_);
  nor _31961_ (_00495_, _00494_, _00493_);
  or _31962_ (_00496_, _00495_, _00289_);
  and _31963_ (_00497_, _00496_, _22762_);
  and _31964_ (_26890_[2], _00497_, _00491_);
  or _31965_ (_00498_, _00331_, _26536_);
  nand _31966_ (_00499_, _00498_, _00329_);
  and _31967_ (_00500_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _31968_ (_00501_, _00500_, _00424_);
  and _31969_ (_00502_, _00501_, _00499_);
  and _31970_ (_00503_, _00330_, _00329_);
  and _31971_ (_00504_, _00503_, _26538_);
  and _31972_ (_00505_, _00501_, _00504_);
  and _31973_ (_00506_, _00505_, _26523_);
  or _31974_ (_00507_, _00506_, _00502_);
  not _31975_ (_00508_, _00507_);
  not _31976_ (_00509_, _00500_);
  nand _31977_ (_00510_, _00509_, _00426_);
  and _31978_ (_00511_, _00510_, _00508_);
  nand _31979_ (_00512_, _00511_, _23596_);
  or _31980_ (_00513_, _26353_, _26328_);
  and _31981_ (_00514_, _26352_, _26348_);
  or _31982_ (_00515_, _00514_, _00513_);
  nand _31983_ (_00516_, _00514_, _00513_);
  nand _31984_ (_00517_, _00516_, _00515_);
  nand _31985_ (_00518_, _00517_, _26366_);
  or _31986_ (_00519_, _26366_, _26327_);
  and _31987_ (_00520_, _00519_, _00518_);
  nand _31988_ (_00521_, _00520_, _23599_);
  nor _31989_ (_00522_, _00199_, _23088_);
  not _31990_ (_00523_, _00522_);
  and _31991_ (_00524_, _23497_, _23491_);
  or _31992_ (_00525_, _00524_, _23481_);
  nor _31993_ (_00526_, _00525_, _23498_);
  not _31994_ (_00527_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _31995_ (_00528_, _23529_, _00527_);
  nor _31996_ (_00529_, _00528_, _23616_);
  and _31997_ (_00530_, _23579_, _23616_);
  nor _31998_ (_00531_, _23530_, _23539_);
  nor _31999_ (_00532_, _00531_, _00530_);
  nor _32000_ (_00533_, _00532_, _00529_);
  not _32001_ (_00534_, _00533_);
  or _32002_ (_00535_, _23603_, _23244_);
  nand _32003_ (_00536_, _23604_, _23326_);
  and _32004_ (_00537_, _00536_, _00535_);
  and _32005_ (_00538_, _00537_, _23736_);
  and _32006_ (_00539_, _00538_, _00534_);
  and _32007_ (_00540_, _00539_, _23725_);
  not _32008_ (_00541_, _00540_);
  nor _32009_ (_00542_, _00541_, _00526_);
  and _32010_ (_00543_, _00542_, _00523_);
  and _32011_ (_00544_, _00543_, _00521_);
  nand _32012_ (_00545_, _00544_, _00512_);
  and _32013_ (_00546_, _00545_, _26612_);
  and _32014_ (_00547_, _00405_, _00019_);
  and _32015_ (_00548_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _32016_ (_00549_, _22768_, _23273_);
  and _32017_ (_00550_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and _32018_ (_00551_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _32019_ (_00552_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _32020_ (_00553_, _00552_, _00551_);
  and _32021_ (_00554_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _32022_ (_00555_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _32023_ (_00556_, _00555_, _00554_);
  and _32024_ (_00557_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _32025_ (_00558_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _32026_ (_00559_, _00558_, _00557_);
  and _32027_ (_00560_, _00559_, _00556_);
  and _32028_ (_00561_, _00560_, _00553_);
  nor _32029_ (_00563_, _00561_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _32030_ (_00564_, _00563_, _00550_);
  nor _32031_ (_00565_, _00564_, _23950_);
  nor _32032_ (_00566_, _00565_, _00549_);
  not _32033_ (_00567_, _00566_);
  and _32034_ (_00568_, _00567_, _26573_);
  or _32035_ (_00569_, _00568_, _00548_);
  or _32036_ (_00570_, _00569_, _00547_);
  or _32037_ (_00571_, _00485_, _00481_);
  and _32038_ (_00572_, _00567_, _26595_);
  and _32039_ (_00573_, _00304_, _00019_);
  nor _32040_ (_00574_, _00573_, _00572_);
  nor _32041_ (_00575_, _00574_, _23268_);
  and _32042_ (_00576_, _00574_, _23268_);
  nor _32043_ (_00577_, _00576_, _00575_);
  nand _32044_ (_00578_, _00577_, _00571_);
  or _32045_ (_00579_, _00577_, _00571_);
  and _32046_ (_00580_, _00579_, _00578_);
  and _32047_ (_00581_, _00580_, _00317_);
  or _32048_ (_00582_, _00581_, _00570_);
  or _32049_ (_00583_, _00582_, _00546_);
  and _32050_ (_00584_, _00583_, _00289_);
  and _32051_ (_00585_, _00493_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _32052_ (_00586_, _00493_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _32053_ (_00587_, _00586_, _00585_);
  and _32054_ (_00588_, _00587_, _00416_);
  or _32055_ (_00589_, _00588_, _00584_);
  and _32056_ (_26890_[3], _00589_, _22762_);
  nand _32057_ (_00590_, _26359_, _26357_);
  or _32058_ (_00591_, _26359_, _26357_);
  and _32059_ (_00592_, _00591_, _00590_);
  or _32060_ (_00593_, _00592_, _00336_);
  or _32061_ (_00594_, _26366_, _26315_);
  and _32062_ (_00595_, _00594_, _00593_);
  and _32063_ (_00596_, _00595_, _23599_);
  and _32064_ (_00597_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _32065_ (_00598_, _00597_, _00507_);
  nor _32066_ (_00599_, _00597_, _00507_);
  nor _32067_ (_00600_, _00599_, _00598_);
  and _32068_ (_00601_, _00600_, _23596_);
  and _32069_ (_00602_, _00196_, _23087_);
  or _32070_ (_00603_, _23501_, _23266_);
  nor _32071_ (_00604_, _23502_, _23481_);
  and _32072_ (_00605_, _00604_, _00603_);
  or _32073_ (_00606_, _23531_, _23525_);
  nor _32074_ (_00607_, _23532_, _23539_);
  and _32075_ (_00608_, _00607_, _00606_);
  and _32076_ (_00609_, _23602_, _23208_);
  and _32077_ (_00610_, _23579_, _23525_);
  nor _32078_ (_00611_, _00359_, _23291_);
  or _32079_ (_00612_, _00611_, _00610_);
  or _32080_ (_00613_, _00612_, _00609_);
  or _32081_ (_00614_, _00613_, _00608_);
  or _32082_ (_00615_, _00614_, _23641_);
  or _32083_ (_00616_, _00615_, _00605_);
  or _32084_ (_00618_, _00616_, _00602_);
  or _32085_ (_00619_, _00618_, _00601_);
  or _32086_ (_00620_, _00619_, _00596_);
  and _32087_ (_00621_, _00620_, _26612_);
  and _32088_ (_00622_, _00405_, _00051_);
  nor _32089_ (_00623_, _22768_, _23225_);
  and _32090_ (_00624_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and _32091_ (_00625_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _32092_ (_00627_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _32093_ (_00628_, _00627_, _00625_);
  and _32094_ (_00629_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _32095_ (_00630_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _32096_ (_00631_, _00630_, _00629_);
  and _32097_ (_00632_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _32098_ (_00633_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _32099_ (_00634_, _00633_, _00632_);
  and _32100_ (_00635_, _00634_, _00631_);
  and _32101_ (_00636_, _00635_, _00628_);
  nor _32102_ (_00637_, _00636_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _32103_ (_00638_, _00637_, _00624_);
  nor _32104_ (_00639_, _00638_, _23950_);
  nor _32105_ (_00640_, _00639_, _00623_);
  not _32106_ (_00641_, _00640_);
  and _32107_ (_00642_, _00641_, _26573_);
  and _32108_ (_00643_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _32109_ (_00644_, _00643_, _00642_);
  or _32110_ (_00645_, _00644_, _00622_);
  and _32111_ (_00646_, _00641_, _26595_);
  and _32112_ (_00647_, _00304_, _00051_);
  nor _32113_ (_00648_, _00647_, _00646_);
  or _32114_ (_00649_, _00648_, _23220_);
  nand _32115_ (_00650_, _00648_, _23220_);
  and _32116_ (_00651_, _00650_, _00649_);
  nor _32117_ (_00652_, _00575_, _00571_);
  nor _32118_ (_00653_, _00652_, _00576_);
  or _32119_ (_00654_, _00653_, _00651_);
  nand _32120_ (_00655_, _00653_, _00651_);
  and _32121_ (_00656_, _00655_, _00317_);
  and _32122_ (_00657_, _00656_, _00654_);
  nor _32123_ (_00658_, _00657_, _00645_);
  nand _32124_ (_00659_, _00658_, _00289_);
  or _32125_ (_00660_, _00659_, _00621_);
  and _32126_ (_00661_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _32127_ (_00662_, _00661_, _00493_);
  nor _32128_ (_00663_, _00585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _32129_ (_00664_, _00663_, _00662_);
  or _32130_ (_00665_, _00664_, _00289_);
  and _32131_ (_00666_, _00665_, _22762_);
  and _32132_ (_26890_[4], _00666_, _00660_);
  and _32133_ (_00667_, _00590_, _26317_);
  nand _32134_ (_00668_, _26319_, _00667_);
  or _32135_ (_00669_, _26319_, _00667_);
  and _32136_ (_00670_, _00669_, _00668_);
  or _32137_ (_00671_, _00670_, _00336_);
  or _32138_ (_00672_, _26366_, _26309_);
  and _32139_ (_00673_, _00672_, _00671_);
  and _32140_ (_00674_, _00673_, _23599_);
  and _32141_ (_00675_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _32142_ (_00676_, _00675_, _00597_);
  nand _32143_ (_00677_, _00676_, _00507_);
  or _32144_ (_00678_, _00675_, _00598_);
  and _32145_ (_00679_, _00678_, _00677_);
  and _32146_ (_00680_, _00679_, _23596_);
  nor _32147_ (_00681_, _23264_, _23219_);
  nor _32148_ (_00682_, _00681_, _23506_);
  or _32149_ (_00683_, _00682_, _23502_);
  nor _32150_ (_00684_, _23503_, _23481_);
  and _32151_ (_00685_, _00684_, _00683_);
  nor _32152_ (_00686_, _00193_, _23088_);
  and _32153_ (_00687_, _23532_, _23208_);
  nor _32154_ (_00688_, _23532_, _23208_);
  nor _32155_ (_00689_, _23523_, _23131_);
  nor _32156_ (_00690_, _00689_, _23531_);
  and _32157_ (_00691_, _00690_, _23521_);
  or _32158_ (_00692_, _00691_, _00688_);
  or _32159_ (_00693_, _00692_, _00687_);
  and _32160_ (_00694_, _00691_, _23522_);
  nor _32161_ (_00695_, _00694_, _23539_);
  and _32162_ (_00696_, _00695_, _00693_);
  and _32163_ (_00697_, _23579_, _23208_);
  nor _32164_ (_00698_, _00359_, _23244_);
  nor _32165_ (_00699_, _23603_, _23171_);
  or _32166_ (_00700_, _00699_, _00698_);
  nor _32167_ (_00701_, _00700_, _00697_);
  nand _32168_ (_00702_, _00701_, _23935_);
  nor _32169_ (_00703_, _00702_, _00696_);
  nand _32170_ (_00704_, _00703_, _23926_);
  or _32171_ (_00705_, _00704_, _00686_);
  or _32172_ (_00706_, _00705_, _00685_);
  or _32173_ (_00707_, _00706_, _00680_);
  or _32174_ (_00708_, _00707_, _00674_);
  and _32175_ (_00709_, _00708_, _26612_);
  nand _32176_ (_00710_, _00655_, _00649_);
  nor _32177_ (_00711_, _22768_, _23188_);
  and _32178_ (_00712_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and _32179_ (_00713_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _32180_ (_00714_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _32181_ (_00715_, _00714_, _00713_);
  and _32182_ (_00716_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _32183_ (_00717_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _32184_ (_00718_, _00717_, _00716_);
  and _32185_ (_00719_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and _32186_ (_00720_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor _32187_ (_00721_, _00720_, _00719_);
  and _32188_ (_00722_, _00721_, _00718_);
  and _32189_ (_00723_, _00722_, _00715_);
  nor _32190_ (_00724_, _00723_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _32191_ (_00725_, _00724_, _00712_);
  nor _32192_ (_00726_, _00725_, _23950_);
  nor _32193_ (_00727_, _00726_, _00711_);
  nor _32194_ (_00728_, _00727_, _00304_);
  and _32195_ (_00729_, _00304_, _00007_);
  nor _32196_ (_00730_, _00729_, _00728_);
  nor _32197_ (_00731_, _00730_, _23183_);
  and _32198_ (_00732_, _00730_, _23183_);
  nor _32199_ (_00733_, _00732_, _00731_);
  or _32200_ (_00734_, _00733_, _00710_);
  and _32201_ (_00735_, _00733_, _00710_);
  not _32202_ (_00736_, _00735_);
  and _32203_ (_00737_, _00736_, _00401_);
  nand _32204_ (_00738_, _00737_, _00734_);
  nand _32205_ (_00739_, _00405_, _00007_);
  and _32206_ (_00741_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _32207_ (_00742_, _00728_, _26570_);
  nor _32208_ (_00743_, _00742_, _00741_);
  and _32209_ (_00744_, _00743_, _00739_);
  and _32210_ (_00745_, _00744_, _00738_);
  nand _32211_ (_00746_, _00745_, _00289_);
  or _32212_ (_00747_, _00746_, _00709_);
  nor _32213_ (_00748_, _00662_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _32214_ (_00749_, _00662_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _32215_ (_00750_, _00749_, _00748_);
  or _32216_ (_00751_, _00750_, _00289_);
  and _32217_ (_00752_, _00751_, _22762_);
  and _32218_ (_26890_[5], _00752_, _00747_);
  not _32219_ (_00753_, _23599_);
  and _32220_ (_00754_, _26363_, _26300_);
  nor _32221_ (_00755_, _26363_, _26300_);
  or _32222_ (_00756_, _00755_, _00754_);
  and _32223_ (_00757_, _00756_, _26366_);
  nor _32224_ (_00758_, _26366_, _26294_);
  or _32225_ (_00759_, _00758_, _00757_);
  or _32226_ (_00760_, _00759_, _00753_);
  and _32227_ (_00761_, _26373_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  not _32228_ (_00762_, _00761_);
  nor _32229_ (_00763_, _00762_, _00677_);
  and _32230_ (_00765_, _00762_, _00677_);
  or _32231_ (_00766_, _00765_, _00763_);
  or _32232_ (_00767_, _00766_, _23597_);
  nor _32233_ (_00768_, _00191_, _23088_);
  not _32234_ (_00769_, _00768_);
  nor _32235_ (_00770_, _23511_, _23503_);
  nor _32236_ (_00771_, _00770_, _23481_);
  and _32237_ (_00772_, _00771_, _23514_);
  and _32238_ (_00773_, _24041_, _24026_);
  not _32239_ (_00774_, _00688_);
  nor _32240_ (_00775_, _00694_, _00774_);
  nor _32241_ (_00776_, _00775_, _24028_);
  not _32242_ (_00777_, _00776_);
  and _32243_ (_00778_, _00775_, _24028_);
  nor _32244_ (_00779_, _00778_, _23539_);
  and _32245_ (_00780_, _00779_, _00777_);
  nand _32246_ (_00781_, _23604_, _23208_);
  or _32247_ (_00782_, _23603_, _23131_);
  and _32248_ (_00783_, _23579_, _24028_);
  not _32249_ (_00784_, _00783_);
  and _32250_ (_00785_, _00784_, _00782_);
  nand _32251_ (_00786_, _00785_, _00781_);
  nor _32252_ (_00787_, _00786_, _00780_);
  and _32253_ (_00788_, _00787_, _00773_);
  not _32254_ (_00789_, _00788_);
  nor _32255_ (_00790_, _00789_, _00772_);
  and _32256_ (_00791_, _00790_, _00769_);
  and _32257_ (_00792_, _00791_, _00767_);
  and _32258_ (_00793_, _00792_, _00760_);
  not _32259_ (_00794_, _00793_);
  and _32260_ (_00795_, _00794_, _26612_);
  and _32261_ (_00796_, _00405_, _26812_);
  and _32262_ (_00797_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _32263_ (_00798_, _22768_, _23152_);
  and _32264_ (_00799_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and _32265_ (_00800_, _23849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _32266_ (_00801_, _23857_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or _32267_ (_00802_, _00801_, _00800_);
  and _32268_ (_00803_, _23846_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _32269_ (_00804_, _23853_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or _32270_ (_00805_, _00804_, _00803_);
  or _32271_ (_00806_, _00805_, _00802_);
  and _32272_ (_00807_, _23842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _32273_ (_00808_, _23844_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _32274_ (_00809_, _00808_, _00807_);
  or _32275_ (_00810_, _00809_, _00806_);
  and _32276_ (_00811_, _00810_, _23839_);
  or _32277_ (_00812_, _00811_, _00799_);
  and _32278_ (_00813_, _00812_, _22768_);
  nor _32279_ (_00814_, _00813_, _00798_);
  not _32280_ (_00815_, _00814_);
  and _32281_ (_00816_, _00815_, _26573_);
  or _32282_ (_00817_, _00816_, _00797_);
  or _32283_ (_00818_, _00817_, _00796_);
  or _32284_ (_00819_, _00735_, _00731_);
  and _32285_ (_00820_, _00815_, _26595_);
  and _32286_ (_00821_, _00304_, _26812_);
  nor _32287_ (_00822_, _00821_, _00820_);
  or _32288_ (_00823_, _00822_, _23147_);
  nand _32289_ (_00824_, _00822_, _23147_);
  and _32290_ (_00825_, _00824_, _00823_);
  or _32291_ (_00826_, _00825_, _00819_);
  nand _32292_ (_00827_, _00825_, _00819_);
  and _32293_ (_00829_, _00827_, _00317_);
  and _32294_ (_00830_, _00829_, _00826_);
  or _32295_ (_00831_, _00830_, _00818_);
  or _32296_ (_00833_, _00831_, _00795_);
  and _32297_ (_00834_, _00833_, _00289_);
  and _32298_ (_00835_, _00749_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _32299_ (_00836_, _00749_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _32300_ (_00837_, _00836_, _00835_);
  and _32301_ (_00838_, _00837_, _00416_);
  or _32302_ (_00839_, _00838_, _00834_);
  and _32303_ (_26890_[6], _00839_, _22762_);
  or _32304_ (_00840_, _26366_, _26286_);
  not _32305_ (_00841_, _00754_);
  nand _32306_ (_00842_, _00841_, _26295_);
  and _32307_ (_00843_, _00842_, _26298_);
  or _32308_ (_00844_, _00843_, _00336_);
  and _32309_ (_00845_, _00844_, _00840_);
  and _32310_ (_00846_, _00845_, _23599_);
  not _32311_ (_00847_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  or _32312_ (_00848_, _26372_, _00847_);
  nor _32313_ (_00849_, _00848_, _00763_);
  and _32314_ (_00850_, _00763_, _00847_);
  or _32315_ (_00851_, _00850_, _00849_);
  and _32316_ (_00852_, _00851_, _23596_);
  and _32317_ (_00853_, _00188_, _23087_);
  nand _32318_ (_00854_, _23516_, _23483_);
  and _32319_ (_00855_, _23518_, _23480_);
  and _32320_ (_00856_, _00855_, _00854_);
  nor _32321_ (_00857_, _00691_, _23533_);
  and _32322_ (_00858_, _00857_, _23131_);
  nor _32323_ (_00859_, _00857_, _23131_);
  or _32324_ (_00860_, _00859_, _00858_);
  and _32325_ (_00861_, _00860_, _23528_);
  and _32326_ (_00862_, _23568_, _23456_);
  and _32327_ (_00863_, _23563_, _23567_);
  and _32328_ (_00864_, _23579_, _23536_);
  nor _32329_ (_00865_, _00359_, _23171_);
  or _32330_ (_00866_, _00865_, _00864_);
  or _32331_ (_00867_, _00866_, _00863_);
  or _32332_ (_00868_, _00867_, _00862_);
  nor _32333_ (_00869_, _00868_, _00861_);
  nand _32334_ (_00870_, _00869_, _23701_);
  or _32335_ (_00871_, _00870_, _00856_);
  or _32336_ (_00872_, _00871_, _00853_);
  or _32337_ (_00873_, _00872_, _00852_);
  or _32338_ (_00875_, _00873_, _00846_);
  and _32339_ (_00876_, _00875_, _26612_);
  and _32340_ (_00877_, _00405_, _26772_);
  nor _32341_ (_00878_, _26574_, _25713_);
  and _32342_ (_00879_, _24628_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _32343_ (_00880_, _00879_, _00878_);
  or _32344_ (_00881_, _00880_, _00877_);
  or _32345_ (_00882_, _00881_, _00876_);
  nand _32346_ (_00883_, _00827_, _00823_);
  nor _32347_ (_00884_, _00304_, _25713_);
  and _32348_ (_00885_, _00304_, _26772_);
  nor _32349_ (_00886_, _00885_, _00884_);
  nor _32350_ (_00887_, _00886_, _23089_);
  and _32351_ (_00888_, _00886_, _23089_);
  nor _32352_ (_00889_, _00888_, _00887_);
  or _32353_ (_00890_, _00889_, _00883_);
  nand _32354_ (_00891_, _00889_, _00883_);
  and _32355_ (_00892_, _00891_, _00890_);
  nand _32356_ (_00893_, _00892_, _00317_);
  nand _32357_ (_00894_, _00893_, _00289_);
  or _32358_ (_00895_, _00894_, _00882_);
  nor _32359_ (_00896_, _00835_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _32360_ (_00897_, _00835_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _32361_ (_00898_, _00897_, _00896_);
  or _32362_ (_00899_, _00898_, _00289_);
  and _32363_ (_00900_, _00899_, _22762_);
  and _32364_ (_26890_[7], _00900_, _00895_);
  and _32365_ (_00901_, _26565_, _24628_);
  nor _32366_ (_00902_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32367_ (_00903_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23370_);
  nor _32368_ (_00904_, _00903_, _00902_);
  not _32369_ (_00905_, _00904_);
  or _32370_ (_00906_, _00905_, _23519_);
  and _32371_ (_00907_, _00905_, _23519_);
  nor _32372_ (_00908_, _00907_, _23481_);
  and _32373_ (_00909_, _00908_, _00906_);
  nand _32374_ (_00910_, _26366_, _23599_);
  nor _32375_ (_00911_, _23540_, _23537_);
  and _32376_ (_00912_, _00911_, _23680_);
  nor _32377_ (_00913_, _00912_, _23397_);
  not _32378_ (_00914_, _23609_);
  and _32379_ (_00915_, _00912_, _23397_);
  or _32380_ (_00916_, _00915_, _00914_);
  nor _32381_ (_00917_, _00916_, _00913_);
  and _32382_ (_00918_, _23579_, _23397_);
  and _32383_ (_00919_, _26399_, _23567_);
  and _32384_ (_00920_, _00919_, _23596_);
  and _32385_ (_00922_, _23571_, _23525_);
  nor _32386_ (_00923_, _23688_, _23392_);
  or _32387_ (_00924_, _00923_, _00922_);
  or _32388_ (_00925_, _00924_, _00920_);
  nor _32389_ (_00926_, _00925_, _00918_);
  not _32390_ (_00927_, _00926_);
  nor _32391_ (_00928_, _00927_, _00917_);
  nand _32392_ (_00929_, _00928_, _00910_);
  or _32393_ (_00930_, _00929_, _00909_);
  and _32394_ (_00931_, _00930_, _26566_);
  and _32395_ (_00932_, _26573_, _00130_);
  not _32396_ (_00933_, _24530_);
  and _32397_ (_00934_, _00405_, _00933_);
  and _32398_ (_00935_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _32399_ (_00936_, _00935_, _00934_);
  or _32400_ (_00937_, _00936_, _00932_);
  or _32401_ (_00938_, _00937_, _00931_);
  or _32402_ (_00939_, _00938_, _00901_);
  not _32403_ (_00940_, _00886_);
  not _32404_ (_00941_, _00888_);
  and _32405_ (_00942_, _00941_, _00883_);
  or _32406_ (_00943_, _00942_, _00887_);
  nand _32407_ (_00944_, _00943_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _32408_ (_00945_, _00943_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _32409_ (_00946_, _00945_, _00944_);
  or _32410_ (_00947_, _00946_, _00940_);
  nand _32411_ (_00948_, _00946_, _00940_);
  and _32412_ (_00949_, _00948_, _00947_);
  and _32413_ (_00950_, _00949_, _00317_);
  or _32414_ (_00951_, _00950_, _00416_);
  or _32415_ (_00952_, _00951_, _00939_);
  nor _32416_ (_00953_, _00897_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _32417_ (_00954_, _00897_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _32418_ (_00955_, _00954_, _00953_);
  or _32419_ (_00956_, _00955_, _00289_);
  and _32420_ (_00957_, _00956_, _22762_);
  and _32421_ (_26890_[8], _00957_, _00952_);
  not _32422_ (_00958_, _26566_);
  nor _32423_ (_00959_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32424_ (_00960_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23338_);
  nor _32425_ (_00961_, _00960_, _00959_);
  not _32426_ (_00962_, _00961_);
  and _32427_ (_00963_, _00962_, _00906_);
  not _32428_ (_00964_, _00963_);
  or _32429_ (_00965_, _00962_, _00906_);
  and _32430_ (_00966_, _00965_, _23480_);
  and _32431_ (_00967_, _00966_, _00964_);
  not _32432_ (_00968_, _00967_);
  and _32433_ (_00969_, _26274_, _23599_);
  not _32434_ (_00970_, _00969_);
  and _32435_ (_00971_, _23579_, _23364_);
  or _32436_ (_00972_, _23418_, _23131_);
  nor _32437_ (_00973_, _00972_, _23678_);
  and _32438_ (_00974_, _00973_, _23521_);
  and _32439_ (_00975_, _23418_, _23131_);
  and _32440_ (_00976_, _00975_, _23674_);
  and _32441_ (_00977_, _00976_, _23456_);
  nor _32442_ (_00978_, _00977_, _00974_);
  nor _32443_ (_00979_, _00978_, _23400_);
  and _32444_ (_00980_, _00978_, _23400_);
  or _32445_ (_00981_, _00980_, _00914_);
  nor _32446_ (_00982_, _00981_, _00979_);
  and _32447_ (_00983_, _26437_, _26404_);
  nor _32448_ (_00984_, _00983_, _26438_);
  and _32449_ (_00985_, _00984_, _23596_);
  and _32450_ (_00986_, _23571_, _23208_);
  and _32451_ (_00987_, _23627_, _23359_);
  or _32452_ (_00988_, _00987_, _00986_);
  or _32453_ (_00989_, _00988_, _00985_);
  or _32454_ (_00990_, _00989_, _00982_);
  nor _32455_ (_00991_, _00990_, _00971_);
  and _32456_ (_00992_, _00991_, _00970_);
  and _32457_ (_00993_, _00992_, _00968_);
  nor _32458_ (_00994_, _00993_, _00958_);
  and _32459_ (_00996_, _26573_, _00095_);
  not _32460_ (_00997_, _24486_);
  and _32461_ (_00998_, _00405_, _00997_);
  or _32462_ (_00999_, _00998_, _00996_);
  and _32463_ (_01000_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _32464_ (_01001_, _01000_, _00999_);
  or _32465_ (_01002_, _01001_, _00994_);
  nor _32466_ (_01003_, _00945_, _00886_);
  nor _32467_ (_01004_, _00944_, _00940_);
  nor _32468_ (_01005_, _01004_, _01003_);
  nand _32469_ (_01006_, _01005_, _23338_);
  or _32470_ (_01007_, _01005_, _23338_);
  and _32471_ (_01008_, _01007_, _00317_);
  and _32472_ (_01009_, _01008_, _01006_);
  or _32473_ (_01010_, _01009_, _01002_);
  not _32474_ (_01011_, _24628_);
  or _32475_ (_01012_, _00372_, _01011_);
  nand _32476_ (_01013_, _01012_, _00289_);
  or _32477_ (_01014_, _01013_, _01010_);
  and _32478_ (_01015_, _00954_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _32479_ (_01016_, _00954_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _32480_ (_01017_, _01016_, _01015_);
  or _32481_ (_01018_, _01017_, _00289_);
  and _32482_ (_01019_, _01018_, _22762_);
  and _32483_ (_26890_[9], _01019_, _01014_);
  and _32484_ (_01021_, _01003_, _23338_);
  and _32485_ (_01022_, _01004_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _32486_ (_01023_, _01022_, _01021_);
  nand _32487_ (_01024_, _01023_, _23309_);
  or _32488_ (_01025_, _01023_, _23309_);
  and _32489_ (_01026_, _01025_, _00401_);
  and _32490_ (_01027_, _01026_, _01024_);
  and _32491_ (_01028_, _00451_, _24628_);
  nor _32492_ (_01029_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32493_ (_01030_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23309_);
  nor _32494_ (_01031_, _01030_, _01029_);
  not _32495_ (_01032_, _01031_);
  and _32496_ (_01033_, _01032_, _00965_);
  not _32497_ (_01034_, _01033_);
  or _32498_ (_01035_, _01032_, _00965_);
  and _32499_ (_01036_, _01035_, _23480_);
  and _32500_ (_01037_, _01036_, _01034_);
  not _32501_ (_01038_, _01037_);
  and _32502_ (_01039_, _00977_, _23400_);
  and _32503_ (_01040_, _00973_, _23364_);
  and _32504_ (_01041_, _01040_, _23521_);
  nor _32505_ (_01042_, _01041_, _01039_);
  and _32506_ (_01043_, _01042_, _23404_);
  nor _32507_ (_01044_, _01042_, _23404_);
  or _32508_ (_01045_, _01044_, _00914_);
  nor _32509_ (_01046_, _01045_, _01043_);
  nor _32510_ (_01047_, _26507_, _26504_);
  nor _32511_ (_01048_, _01047_, _26508_);
  and _32512_ (_01049_, _01048_, _23596_);
  nand _32513_ (_01050_, _00865_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _32514_ (_01051_, _23627_, _23326_);
  and _32515_ (_01052_, _23579_, _23332_);
  and _32516_ (_01053_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or _32517_ (_01054_, _01053_, _01052_);
  nor _32518_ (_01055_, _01054_, _01051_);
  and _32519_ (_01056_, _01055_, _01050_);
  not _32520_ (_01057_, _01056_);
  nor _32521_ (_01058_, _01057_, _01049_);
  not _32522_ (_01059_, _01058_);
  nor _32523_ (_01060_, _01059_, _01046_);
  and _32524_ (_01061_, _01060_, _01038_);
  nor _32525_ (_01062_, _01061_, _00958_);
  and _32526_ (_01063_, _26573_, _00164_);
  not _32527_ (_01064_, _24508_);
  and _32528_ (_01065_, _00405_, _01064_);
  or _32529_ (_01066_, _01065_, _01063_);
  and _32530_ (_01067_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _32531_ (_01068_, _01067_, _01066_);
  nor _32532_ (_01069_, _01068_, _01062_);
  nand _32533_ (_01070_, _01069_, _00289_);
  or _32534_ (_01071_, _01070_, _01028_);
  or _32535_ (_01072_, _01071_, _01027_);
  nor _32536_ (_01073_, _01015_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _32537_ (_01074_, _01015_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _32538_ (_01075_, _01074_, _01073_);
  or _32539_ (_01076_, _01075_, _00289_);
  and _32540_ (_01077_, _01076_, _22762_);
  and _32541_ (_26890_[10], _01077_, _01072_);
  and _32542_ (_01078_, _01074_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _32543_ (_01079_, _01074_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _32544_ (_01080_, _01079_, _01078_);
  or _32545_ (_01081_, _00898_, _00837_);
  and _32546_ (_01082_, _00495_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _32547_ (_01083_, _00955_, _00587_);
  or _32548_ (_01084_, _01083_, _01082_);
  or _32549_ (_01085_, _01017_, _00664_);
  or _32550_ (_01086_, _01085_, _01084_);
  or _32551_ (_01087_, _01075_, _00750_);
  or _32552_ (_01088_, _01087_, _01086_);
  or _32553_ (_01089_, _01088_, _01081_);
  and _32554_ (_01090_, _01089_, _01080_);
  nor _32555_ (_01091_, _01089_, _01080_);
  or _32556_ (_01092_, _01091_, _01090_);
  nand _32557_ (_01093_, _01092_, _00306_);
  and _32558_ (_01094_, _00545_, _24628_);
  nor _32559_ (_01095_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32560_ (_01096_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23270_);
  nor _32561_ (_01097_, _01096_, _01095_);
  not _32562_ (_01098_, _01097_);
  and _32563_ (_01099_, _01098_, _01035_);
  nor _32564_ (_01100_, _01098_, _01035_);
  nor _32565_ (_01101_, _01100_, _01099_);
  and _32566_ (_01102_, _01101_, _23480_);
  not _32567_ (_01103_, _01102_);
  and _32568_ (_01105_, _26511_, _26509_);
  not _32569_ (_01106_, _01105_);
  and _32570_ (_01107_, _01106_, _26512_);
  and _32571_ (_01108_, _01107_, _23596_);
  not _32572_ (_01109_, _01108_);
  and _32573_ (_01110_, _01040_, _23332_);
  nor _32574_ (_01111_, _01110_, _23456_);
  and _32575_ (_01112_, _23400_, _23404_);
  and _32576_ (_01113_, _01112_, _00976_);
  nor _32577_ (_01114_, _01113_, _23521_);
  or _32578_ (_01115_, _01114_, _01111_);
  and _32579_ (_01116_, _01115_, _23296_);
  nor _32580_ (_01117_, _01115_, _23296_);
  nor _32581_ (_01118_, _01117_, _01116_);
  and _32582_ (_01119_, _01118_, _23609_);
  and _32583_ (_01120_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor _32584_ (_01121_, _23688_, _23291_);
  and _32585_ (_01122_, _23579_, _23462_);
  or _32586_ (_01123_, _01122_, _01121_);
  or _32587_ (_01124_, _01123_, _23572_);
  nor _32588_ (_01125_, _01124_, _01120_);
  not _32589_ (_01126_, _01125_);
  nor _32590_ (_01127_, _01126_, _01119_);
  and _32591_ (_01128_, _01127_, _01109_);
  and _32592_ (_01129_, _01128_, _01103_);
  nor _32593_ (_01131_, _01129_, _00958_);
  and _32594_ (_01132_, _26573_, _00019_);
  and _32595_ (_01133_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _32596_ (_01134_, _01133_, _01132_);
  or _32597_ (_01135_, _01134_, _01131_);
  nor _32598_ (_01136_, _01135_, _01094_);
  and _32599_ (_01137_, _01136_, _01093_);
  nand _32600_ (_01138_, _01137_, _00289_);
  nor _32601_ (_01139_, \oc8051_top_1.oc8051_memory_interface1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _32602_ (_01140_, _01139_, _01003_);
  nand _32603_ (_01141_, \oc8051_top_1.oc8051_memory_interface1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _32604_ (_01142_, _01141_, _00944_);
  nor _32605_ (_01143_, _01142_, _00940_);
  nor _32606_ (_01144_, _01143_, _01140_);
  nand _32607_ (_01145_, _01144_, _23270_);
  or _32608_ (_01146_, _01144_, _23270_);
  and _32609_ (_01147_, _01146_, _01145_);
  and _32610_ (_01148_, _01147_, _00317_);
  or _32611_ (_01149_, _01148_, _01138_);
  or _32612_ (_01150_, _01080_, _00289_);
  and _32613_ (_01151_, _01150_, _22762_);
  and _32614_ (_26890_[11], _01151_, _01149_);
  not _32615_ (_01152_, _01091_);
  and _32616_ (_01153_, _01078_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _32617_ (_01154_, _01078_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _32618_ (_01155_, _01154_, _01153_);
  and _32619_ (_01156_, _01155_, _01152_);
  nor _32620_ (_01157_, _01155_, _01152_);
  or _32621_ (_01158_, _01157_, _01156_);
  and _32622_ (_01159_, _01158_, _00306_);
  and _32623_ (_01160_, _00620_, _24628_);
  nor _32624_ (_01161_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32625_ (_01162_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23222_);
  nor _32626_ (_01163_, _01162_, _01161_);
  or _32627_ (_01164_, _01163_, _01100_);
  and _32628_ (_01165_, _01163_, _01100_);
  nor _32629_ (_01166_, _01165_, _23481_);
  and _32630_ (_01167_, _01166_, _01164_);
  or _32631_ (_01168_, _26515_, _26513_);
  and _32632_ (_01169_, _01168_, _26516_);
  and _32633_ (_01170_, _01169_, _23596_);
  and _32634_ (_01171_, _01113_, _23296_);
  and _32635_ (_01172_, _01171_, _23456_);
  and _32636_ (_01173_, _01110_, _23462_);
  and _32637_ (_01174_, _01173_, _23521_);
  nor _32638_ (_01175_, _01174_, _01172_);
  nand _32639_ (_01176_, _01175_, _23263_);
  or _32640_ (_01177_, _01175_, _23263_);
  and _32641_ (_01178_, _01177_, _23609_);
  and _32642_ (_01179_, _01178_, _01176_);
  and _32643_ (_01180_, _23456_, _23525_);
  and _32644_ (_01181_, _23521_, _23250_);
  or _32645_ (_01182_, _01181_, _01180_);
  and _32646_ (_01183_, _01182_, _23627_);
  and _32647_ (_01184_, _23571_, _23567_);
  and _32648_ (_01185_, _23579_, _23250_);
  and _32649_ (_01186_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or _32650_ (_01187_, _01186_, _01185_);
  or _32651_ (_01188_, _01187_, _01184_);
  or _32652_ (_01189_, _01188_, _01183_);
  or _32653_ (_01190_, _01189_, _01179_);
  or _32654_ (_01191_, _01190_, _01170_);
  or _32655_ (_01192_, _01191_, _01167_);
  and _32656_ (_01193_, _01192_, _26566_);
  and _32657_ (_01194_, _26573_, _00051_);
  and _32658_ (_01195_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _32659_ (_01196_, _01195_, _01194_);
  or _32660_ (_01197_, _01196_, _01193_);
  or _32661_ (_01198_, _01197_, _01160_);
  nor _32662_ (_01199_, _01198_, _01159_);
  nand _32663_ (_01200_, _01199_, _00289_);
  and _32664_ (_01201_, _01139_, _23270_);
  and _32665_ (_01202_, _01201_, _01003_);
  or _32666_ (_01203_, _01142_, _23270_);
  nor _32667_ (_01204_, _01203_, _00940_);
  nor _32668_ (_01205_, _01204_, _01202_);
  nand _32669_ (_01206_, _01205_, _23222_);
  or _32670_ (_01207_, _01205_, _23222_);
  and _32671_ (_01208_, _01207_, _01206_);
  and _32672_ (_01209_, _01208_, _00317_);
  or _32673_ (_01210_, _01209_, _01200_);
  or _32674_ (_01211_, _01155_, _00289_);
  and _32675_ (_01212_, _01211_, _22762_);
  and _32676_ (_26890_[12], _01212_, _01210_);
  or _32677_ (_01213_, _01203_, _23222_);
  nor _32678_ (_01214_, _01213_, _00940_);
  and _32679_ (_01215_, _01201_, _23222_);
  and _32680_ (_01216_, _01215_, _01003_);
  nor _32681_ (_01217_, _01216_, _01214_);
  nand _32682_ (_01218_, _01217_, _23185_);
  or _32683_ (_01219_, _01217_, _23185_);
  and _32684_ (_01220_, _01219_, _00401_);
  and _32685_ (_01221_, _01220_, _01218_);
  and _32686_ (_01222_, _00708_, _24628_);
  nor _32687_ (_01223_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32688_ (_01224_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23185_);
  nor _32689_ (_01225_, _01224_, _01223_);
  or _32690_ (_01226_, _01225_, _01165_);
  nand _32691_ (_01227_, _01225_, _01165_);
  and _32692_ (_01228_, _01227_, _23480_);
  and _32693_ (_01229_, _01228_, _01226_);
  or _32694_ (_01230_, _26517_, _26493_);
  and _32695_ (_01231_, _01230_, _26518_);
  and _32696_ (_01232_, _01231_, _23596_);
  and _32697_ (_01233_, _23296_, _23263_);
  and _32698_ (_01234_, _01233_, _01113_);
  nor _32699_ (_01235_, _01234_, _23521_);
  and _32700_ (_01236_, _01173_, _23250_);
  nor _32701_ (_01237_, _01236_, _23456_);
  nor _32702_ (_01238_, _01237_, _01235_);
  nand _32703_ (_01239_, _01238_, _23216_);
  or _32704_ (_01240_, _01238_, _23216_);
  and _32705_ (_01241_, _01240_, _23609_);
  and _32706_ (_01242_, _01241_, _01239_);
  and _32707_ (_01243_, _23521_, _23216_);
  and _32708_ (_01244_, _23456_, _23208_);
  or _32709_ (_01245_, _01244_, _01243_);
  and _32710_ (_01246_, _01245_, _23627_);
  and _32711_ (_01247_, _23571_, _23359_);
  and _32712_ (_01248_, _23579_, _23216_);
  and _32713_ (_01249_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or _32714_ (_01250_, _01249_, _01248_);
  or _32715_ (_01251_, _01250_, _01247_);
  or _32716_ (_01252_, _01251_, _01246_);
  or _32717_ (_01253_, _01252_, _01242_);
  or _32718_ (_01254_, _01253_, _01232_);
  or _32719_ (_01255_, _01254_, _01229_);
  and _32720_ (_01256_, _01255_, _26566_);
  and _32721_ (_01257_, _26573_, _00007_);
  not _32722_ (_01258_, _01157_);
  or _32723_ (_01259_, _01153_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand _32724_ (_01260_, _01153_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _32725_ (_01261_, _01260_, _01259_);
  and _32726_ (_01262_, _01261_, _01258_);
  nor _32727_ (_01263_, _01261_, _01258_);
  or _32728_ (_01264_, _01263_, _01262_);
  and _32729_ (_01265_, _01264_, _00405_);
  or _32730_ (_01266_, _01265_, _01257_);
  and _32731_ (_01267_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _32732_ (_01268_, _01267_, _01266_);
  nor _32733_ (_01269_, _01268_, _01256_);
  nand _32734_ (_01270_, _01269_, _00289_);
  or _32735_ (_01271_, _01270_, _01222_);
  or _32736_ (_01272_, _01271_, _01221_);
  or _32737_ (_01273_, _01261_, _00289_);
  and _32738_ (_01274_, _01273_, _22762_);
  and _32739_ (_26890_[13], _01274_, _01272_);
  nor _32740_ (_01275_, _00793_, _01011_);
  nor _32741_ (_01276_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _32742_ (_01278_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23149_);
  nor _32743_ (_01279_, _01278_, _01276_);
  not _32744_ (_01280_, _01279_);
  and _32745_ (_01281_, _01280_, _01227_);
  not _32746_ (_01282_, _01281_);
  or _32747_ (_01283_, _01280_, _01227_);
  and _32748_ (_01284_, _01283_, _23480_);
  and _32749_ (_01286_, _01284_, _01282_);
  not _32750_ (_01287_, _01286_);
  and _32751_ (_01288_, _26519_, _26487_);
  not _32752_ (_01289_, _01288_);
  and _32753_ (_01290_, _01289_, _26520_);
  and _32754_ (_01291_, _01290_, _23596_);
  and _32755_ (_01292_, _01236_, _23216_);
  and _32756_ (_01293_, _01292_, _23521_);
  and _32757_ (_01294_, _01234_, _23214_);
  and _32758_ (_01295_, _01294_, _23456_);
  or _32759_ (_01297_, _01295_, _01293_);
  and _32760_ (_01298_, _01297_, _23177_);
  nor _32761_ (_01299_, _01297_, _23177_);
  nor _32762_ (_01300_, _01299_, _01298_);
  and _32763_ (_01301_, _01300_, _23609_);
  and _32764_ (_01302_, _23521_, _23179_);
  not _32765_ (_01303_, _01302_);
  and _32766_ (_01304_, _23456_, _23171_);
  nor _32767_ (_01305_, _01304_, _23688_);
  and _32768_ (_01306_, _01305_, _01303_);
  and _32769_ (_01307_, _23579_, _23177_);
  and _32770_ (_01308_, _23571_, _23326_);
  and _32771_ (_01309_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  or _32772_ (_01310_, _01309_, _01308_);
  nor _32773_ (_01311_, _01310_, _01307_);
  not _32774_ (_01312_, _01311_);
  nor _32775_ (_01313_, _01312_, _01306_);
  not _32776_ (_01314_, _01313_);
  nor _32777_ (_01315_, _01314_, _01301_);
  not _32778_ (_01316_, _01315_);
  nor _32779_ (_01317_, _01316_, _01291_);
  and _32780_ (_01318_, _01317_, _01287_);
  nor _32781_ (_01319_, _01318_, _00958_);
  and _32782_ (_01320_, _26573_, _26812_);
  and _32783_ (_01321_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _32784_ (_01322_, _01321_, _01320_);
  or _32785_ (_01323_, _01322_, _01319_);
  or _32786_ (_01324_, _01323_, _01275_);
  or _32787_ (_01325_, _00945_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _32788_ (_01326_, _01325_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _32789_ (_01327_, _01326_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _32790_ (_01328_, _01327_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _32791_ (_01329_, _01328_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _32792_ (_01330_, _01329_, _00886_);
  or _32793_ (_01331_, _01213_, _23185_);
  or _32794_ (_01332_, _01331_, _00940_);
  and _32795_ (_01333_, _01332_, _01330_);
  nand _32796_ (_01334_, _01333_, _23149_);
  or _32797_ (_01335_, _01333_, _23149_);
  and _32798_ (_01336_, _01335_, _00317_);
  and _32799_ (_01337_, _01336_, _01334_);
  or _32800_ (_01338_, _01337_, _01324_);
  not _32801_ (_01339_, _01263_);
  and _32802_ (_01340_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _32803_ (_01341_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _32804_ (_01342_, _01341_, _01074_);
  and _32805_ (_01343_, _01342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _32806_ (_01345_, _01342_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _32807_ (_01346_, _01345_, _01343_);
  and _32808_ (_01347_, _01346_, _01339_);
  nor _32809_ (_01349_, _01346_, _01339_);
  or _32810_ (_01350_, _01349_, _01347_);
  nand _32811_ (_01351_, _01350_, _00306_);
  nand _32812_ (_01352_, _01351_, _00289_);
  or _32813_ (_01353_, _01352_, _01338_);
  or _32814_ (_01354_, _01346_, _00289_);
  and _32815_ (_01355_, _01354_, _22762_);
  and _32816_ (_26890_[14], _01355_, _01353_);
  not _32817_ (_01356_, _24402_);
  not _32818_ (_01357_, _24352_);
  nor _32819_ (_01358_, _01357_, _23866_);
  and _32820_ (_01359_, _01358_, _24436_);
  and _32821_ (_01360_, _01359_, _01356_);
  nor _32822_ (_01361_, _24530_, _24486_);
  and _32823_ (_01362_, _01361_, _01064_);
  and _32824_ (_01363_, _01362_, _01360_);
  nor _32825_ (_01364_, _01064_, _24486_);
  and _32826_ (_01365_, _01364_, _00933_);
  not _32827_ (_01366_, _01365_);
  nor _32828_ (_01367_, _24436_, _01357_);
  and _32829_ (_01368_, _01367_, _23866_);
  nor _32830_ (_01369_, _01368_, _01359_);
  nor _32831_ (_01370_, _01369_, _01366_);
  nor _32832_ (_01371_, _01370_, _01363_);
  nor _32833_ (_01373_, _01371_, _24464_);
  not _32834_ (_01374_, _01373_);
  nor _32835_ (_01375_, _00933_, _24464_);
  and _32836_ (_01376_, _01375_, _01364_);
  and _32837_ (_01377_, _01368_, _24402_);
  and _32838_ (_01378_, _24508_, _24486_);
  and _32839_ (_01379_, _01378_, _24530_);
  and _32840_ (_01380_, _01379_, _01377_);
  nor _32841_ (_01381_, _01380_, _01376_);
  and _32842_ (_01383_, _01359_, _24402_);
  nor _32843_ (_01385_, _01383_, _01377_);
  nor _32844_ (_01387_, _01385_, _01381_);
  not _32845_ (_01388_, _01387_);
  not _32846_ (_01389_, _01360_);
  nor _32847_ (_01390_, _24508_, _24486_);
  and _32848_ (_01391_, _01390_, _01375_);
  not _32849_ (_01392_, _01391_);
  and _32850_ (_01394_, _01064_, _24486_);
  and _32851_ (_01395_, _01394_, _24530_);
  and _32852_ (_01397_, _01395_, _24464_);
  nor _32853_ (_01398_, _01397_, _01378_);
  and _32854_ (_01399_, _01398_, _01392_);
  nor _32855_ (_01400_, _01399_, _01389_);
  and _32856_ (_01401_, _01368_, _01356_);
  and _32857_ (_01402_, _01401_, _01376_);
  and _32858_ (_01403_, _24436_, _23866_);
  and _32859_ (_01404_, _24464_, _24352_);
  and _32860_ (_01405_, _01404_, _01403_);
  and _32861_ (_01406_, _01394_, _00933_);
  nor _32862_ (_01408_, _01406_, _01365_);
  not _32863_ (_01409_, _01408_);
  and _32864_ (_01410_, _01409_, _01405_);
  nor _32865_ (_01411_, _01410_, _01402_);
  not _32866_ (_01413_, _01411_);
  nor _32867_ (_01414_, _01413_, _01400_);
  and _32868_ (_01415_, _01414_, _01388_);
  and _32869_ (_01416_, _01415_, _01374_);
  and _32870_ (_01417_, _24530_, _24464_);
  and _32871_ (_01418_, _01417_, _01364_);
  and _32872_ (_01420_, _01418_, _01401_);
  not _32873_ (_01421_, _01420_);
  and _32874_ (_01422_, _01390_, _01417_);
  and _32875_ (_01423_, _01422_, _01360_);
  not _32876_ (_01424_, _23866_);
  and _32877_ (_01425_, _01367_, _01424_);
  and _32878_ (_01426_, _01425_, _24402_);
  and _32879_ (_01427_, _00933_, _24464_);
  not _32880_ (_01428_, _01427_);
  not _32881_ (_01429_, _01378_);
  nor _32882_ (_01430_, _01429_, _01375_);
  and _32883_ (_01431_, _01430_, _01428_);
  and _32884_ (_01432_, _01431_, _01426_);
  and _32885_ (_01433_, _01406_, _24464_);
  and _32886_ (_01434_, _01433_, _01359_);
  or _32887_ (_01435_, _01434_, _01432_);
  nor _32888_ (_01436_, _01435_, _01423_);
  and _32889_ (_01437_, _01436_, _01421_);
  not _32890_ (_01439_, _01418_);
  nor _32891_ (_01440_, _01377_, _01359_);
  nor _32892_ (_01441_, _01440_, _01439_);
  not _32893_ (_01442_, _01426_);
  and _32894_ (_01443_, _24530_, _00997_);
  and _32895_ (_01444_, _01443_, _01064_);
  nor _32896_ (_01445_, _01444_, _01376_);
  nor _32897_ (_01446_, _01433_, _01395_);
  and _32898_ (_01447_, _01446_, _01445_);
  not _32899_ (_01448_, _24464_);
  and _32900_ (_01449_, _01406_, _01448_);
  and _32901_ (_01450_, _01427_, _01378_);
  nor _32902_ (_01451_, _01450_, _01418_);
  not _32903_ (_01453_, _01451_);
  nor _32904_ (_01454_, _01453_, _01449_);
  and _32905_ (_01456_, _01454_, _01447_);
  nor _32906_ (_01458_, _01456_, _01442_);
  nor _32907_ (_01459_, _01458_, _01441_);
  not _32908_ (_01460_, _01406_);
  and _32909_ (_01461_, _01365_, _24464_);
  nor _32910_ (_01462_, _01461_, _01422_);
  and _32911_ (_01463_, _01462_, _01460_);
  nor _32912_ (_01464_, _01463_, _24352_);
  not _32913_ (_01465_, _01377_);
  nor _32914_ (_01467_, _01433_, _01391_);
  and _32915_ (_01468_, _01467_, _01462_);
  nor _32916_ (_01469_, _01468_, _01465_);
  nor _32917_ (_01470_, _01469_, _01464_);
  and _32918_ (_01471_, _01470_, _01459_);
  and _32919_ (_01472_, _01394_, _01375_);
  and _32920_ (_01473_, _01472_, _01377_);
  and _32921_ (_01474_, _01426_, _01365_);
  nor _32922_ (_01475_, _01474_, _01473_);
  or _32923_ (_01476_, _01449_, _01397_);
  and _32924_ (_01477_, _01476_, _01377_);
  and _32925_ (_01478_, _01378_, _00933_);
  not _32926_ (_01479_, _01478_);
  nor _32927_ (_01480_, _01461_, _01397_);
  and _32928_ (_01481_, _01480_, _01479_);
  not _32929_ (_01482_, _01481_);
  and _32930_ (_01483_, _01482_, _01383_);
  nor _32931_ (_01484_, _01483_, _01477_);
  and _32932_ (_01485_, _01484_, _01475_);
  and _32933_ (_01486_, _01403_, _24352_);
  and _32934_ (_01487_, _01394_, _01448_);
  and _32935_ (_01488_, _01487_, _01486_);
  not _32936_ (_01489_, _01488_);
  and _32937_ (_01490_, _01472_, _01357_);
  and _32938_ (_01491_, _01425_, _01356_);
  nor _32939_ (_01492_, _01491_, _01490_);
  and _32940_ (_01493_, _01492_, _01489_);
  nor _32941_ (_01494_, _01472_, _01461_);
  nor _32942_ (_01496_, _01494_, _01389_);
  and _32943_ (_01497_, _01362_, _24464_);
  nor _32944_ (_01498_, _01497_, _01376_);
  nor _32945_ (_01499_, _01498_, _01389_);
  nor _32946_ (_01500_, _01499_, _01496_);
  and _32947_ (_01501_, _01500_, _01493_);
  and _32948_ (_01502_, _01501_, _01485_);
  and _32949_ (_01503_, _01502_, _01471_);
  and _32950_ (_01504_, _01503_, _01437_);
  and _32951_ (_01505_, _01504_, _01416_);
  and _32952_ (_01506_, _01365_, _01448_);
  and _32953_ (_01507_, _01506_, _01401_);
  or _32954_ (_01508_, _01403_, _01357_);
  and _32955_ (_01509_, _01508_, _01433_);
  or _32956_ (_01510_, _01509_, _01507_);
  nor _32957_ (_01511_, _01510_, _01496_);
  or _32958_ (_01512_, _01450_, _01397_);
  and _32959_ (_01513_, _01512_, _01426_);
  or _32960_ (_01514_, _01402_, _01380_);
  nor _32961_ (_01515_, _01514_, _01513_);
  and _32962_ (_01516_, _01515_, _01511_);
  nand _32963_ (_01517_, _01516_, _01437_);
  nor _32964_ (_01518_, _01517_, _01505_);
  and _32965_ (_01519_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _32966_ (_01520_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _32967_ (_01522_, _01520_, _01519_);
  not _32968_ (_01523_, _01522_);
  nand _32969_ (_01525_, _01523_, _01518_);
  nor _32970_ (_01526_, _01523_, _01518_);
  nor _32971_ (_01527_, _01526_, _25729_);
  and _32972_ (_01528_, _01527_, _01525_);
  nor _32973_ (_01529_, _25728_, _23368_);
  or _32974_ (_01530_, _01529_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _32975_ (_01531_, _01530_, _01528_);
  not _32976_ (_01532_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _32977_ (_01533_, _01532_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _32978_ (_01534_, _01533_, _22762_);
  and _32979_ (_26891_[0], _01534_, _01531_);
  and _32980_ (_01535_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _32981_ (_01536_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _32982_ (_01537_, _01536_, _01535_);
  and _32983_ (_01539_, _01537_, _01519_);
  nor _32984_ (_01540_, _01537_, _01519_);
  nor _32985_ (_01541_, _01540_, _01539_);
  not _32986_ (_01543_, _01541_);
  nor _32987_ (_01544_, _01543_, _01505_);
  and _32988_ (_01545_, _01543_, _01505_);
  nor _32989_ (_01546_, _01545_, _01544_);
  nand _32990_ (_01547_, _01546_, _01526_);
  or _32991_ (_01548_, _01546_, _01526_);
  and _32992_ (_01549_, _01548_, _01547_);
  or _32993_ (_01550_, _01549_, _25729_);
  or _32994_ (_01551_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _32995_ (_01552_, _01551_, _01532_);
  and _32996_ (_01553_, _01552_, _01550_);
  and _32997_ (_01554_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _32998_ (_01555_, _01554_, _01553_);
  and _32999_ (_26891_[1], _01555_, _22762_);
  not _33000_ (_01556_, _01544_);
  and _33001_ (_01557_, _01547_, _01556_);
  not _33002_ (_01558_, _01557_);
  nor _33003_ (_01559_, _01539_, _01535_);
  and _33004_ (_01560_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _33005_ (_01561_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _33006_ (_01562_, _01561_, _01560_);
  not _33007_ (_01563_, _01562_);
  nor _33008_ (_01564_, _01563_, _01559_);
  and _33009_ (_01565_, _01563_, _01559_);
  nor _33010_ (_01567_, _01565_, _01564_);
  and _33011_ (_01568_, _01567_, _01558_);
  nor _33012_ (_01569_, _01567_, _01558_);
  nor _33013_ (_01570_, _01569_, _01568_);
  or _33014_ (_01571_, _01570_, _25729_);
  or _33015_ (_01572_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _33016_ (_01573_, _01572_, _01532_);
  and _33017_ (_01574_, _01573_, _01571_);
  and _33018_ (_01575_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33019_ (_01576_, _01575_, _01574_);
  and _33020_ (_26891_[2], _01576_, _22762_);
  nor _33021_ (_01577_, _01564_, _01560_);
  nor _33022_ (_01578_, _01577_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _33023_ (_01579_, _01577_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _33024_ (_01580_, _01579_, _01578_);
  and _33025_ (_01581_, _01580_, _01568_);
  nor _33026_ (_01582_, _01580_, _01568_);
  nor _33027_ (_01583_, _01582_, _01581_);
  or _33028_ (_01584_, _01583_, _25729_);
  or _33029_ (_01585_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _33030_ (_01586_, _01585_, _01532_);
  and _33031_ (_01587_, _01586_, _01584_);
  and _33032_ (_01588_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33033_ (_01589_, _01588_, _01587_);
  and _33034_ (_26891_[3], _01589_, _22762_);
  nor _33035_ (_01590_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _33036_ (_01591_, _01590_, _00661_);
  nand _33037_ (_01592_, _01591_, _01578_);
  or _33038_ (_01593_, _01591_, _01578_);
  and _33039_ (_01594_, _01593_, _01592_);
  and _33040_ (_01595_, _01594_, _01581_);
  nor _33041_ (_01596_, _01594_, _01581_);
  nor _33042_ (_01597_, _01596_, _01595_);
  or _33043_ (_01598_, _01597_, _25729_);
  or _33044_ (_01599_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _33045_ (_01600_, _01599_, _01532_);
  and _33046_ (_01601_, _01600_, _01598_);
  and _33047_ (_01602_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33048_ (_01603_, _01602_, _01601_);
  and _33049_ (_26891_[4], _01603_, _22762_);
  or _33050_ (_01604_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _01532_);
  and _33051_ (_01605_, _01604_, _22762_);
  nand _33052_ (_01606_, _01590_, _01577_);
  and _33053_ (_01607_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not _33054_ (_01608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _33055_ (_01609_, _01590_, _01608_);
  and _33056_ (_01610_, _01609_, _01577_);
  or _33057_ (_01611_, _01610_, _01607_);
  or _33058_ (_01612_, _01611_, _01595_);
  and _33059_ (_01613_, _01611_, _01594_);
  and _33060_ (_01614_, _01613_, _01581_);
  nor _33061_ (_01615_, _01614_, _25729_);
  and _33062_ (_01616_, _01615_, _01612_);
  nor _33063_ (_01617_, _25728_, _23183_);
  or _33064_ (_01618_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33065_ (_01619_, _01618_, _01616_);
  and _33066_ (_26891_[5], _01619_, _01605_);
  not _33067_ (_01620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _33068_ (_01621_, _01610_, _01620_);
  and _33069_ (_01622_, _01609_, _01620_);
  and _33070_ (_01623_, _01622_, _01577_);
  nor _33071_ (_01624_, _01623_, _01621_);
  not _33072_ (_01625_, _01624_);
  and _33073_ (_01626_, _01625_, _01614_);
  or _33074_ (_01627_, _01625_, _01614_);
  nand _33075_ (_01628_, _01627_, _25728_);
  nor _33076_ (_01629_, _01628_, _01626_);
  nor _33077_ (_01630_, _25728_, _23147_);
  or _33078_ (_01631_, _01630_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33079_ (_01632_, _01631_, _01629_);
  or _33080_ (_01633_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _01532_);
  and _33081_ (_01634_, _01633_, _22762_);
  and _33082_ (_26891_[6], _01634_, _01632_);
  not _33083_ (_01635_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _33084_ (_01636_, _01623_, _01635_);
  and _33085_ (_01637_, _01622_, _01635_);
  and _33086_ (_01638_, _01637_, _01577_);
  nor _33087_ (_01639_, _01638_, _01636_);
  not _33088_ (_01640_, _01639_);
  and _33089_ (_01641_, _01640_, _01626_);
  nor _33090_ (_01642_, _01640_, _01626_);
  nor _33091_ (_01643_, _01642_, _01641_);
  or _33092_ (_01644_, _01643_, _25729_);
  or _33093_ (_01645_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _33094_ (_01646_, _01645_, _01532_);
  and _33095_ (_01647_, _01646_, _01644_);
  and _33096_ (_01648_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _33097_ (_01649_, _01648_, _01647_);
  and _33098_ (_26891_[7], _01649_, _22762_);
  not _33099_ (_01650_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _33100_ (_01651_, _01638_, _01650_);
  and _33101_ (_01652_, _01637_, _01650_);
  and _33102_ (_01653_, _01652_, _01577_);
  or _33103_ (_01654_, _01653_, _01651_);
  and _33104_ (_01655_, _01654_, _01641_);
  nor _33105_ (_01656_, _01654_, _01641_);
  nor _33106_ (_01657_, _01656_, _01655_);
  or _33107_ (_01658_, _01657_, _25729_);
  or _33108_ (_01659_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _33109_ (_01660_, _01659_, _01532_);
  and _33110_ (_01661_, _01660_, _01658_);
  and _33111_ (_01662_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33112_ (_01663_, _01662_, _01661_);
  and _33113_ (_26891_[8], _01663_, _22762_);
  or _33114_ (_01664_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _01532_);
  and _33115_ (_01665_, _01664_, _22762_);
  not _33116_ (_01666_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _33117_ (_01667_, _01652_, _01666_);
  and _33118_ (_01668_, _01667_, _01577_);
  nor _33119_ (_01669_, _01653_, _01666_);
  nor _33120_ (_01670_, _01669_, _01668_);
  not _33121_ (_01671_, _01670_);
  and _33122_ (_01672_, _01671_, _01655_);
  or _33123_ (_01673_, _01671_, _01655_);
  nand _33124_ (_01674_, _01673_, _25728_);
  nor _33125_ (_01675_, _01674_, _01672_);
  nor _33126_ (_01676_, _25728_, _23338_);
  or _33127_ (_01677_, _01676_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33128_ (_01678_, _01677_, _01675_);
  and _33129_ (_26891_[9], _01678_, _01665_);
  not _33130_ (_01679_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _33131_ (_01680_, _01668_, _01679_);
  and _33132_ (_01681_, _01667_, _01679_);
  and _33133_ (_01682_, _01681_, _01577_);
  nor _33134_ (_01683_, _01682_, _01680_);
  not _33135_ (_01684_, _01683_);
  and _33136_ (_01685_, _01684_, _01672_);
  nor _33137_ (_01686_, _01684_, _01672_);
  nor _33138_ (_01687_, _01686_, _01685_);
  or _33139_ (_01688_, _01687_, _25729_);
  or _33140_ (_01689_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _33141_ (_01691_, _01689_, _01532_);
  and _33142_ (_01692_, _01691_, _01688_);
  and _33143_ (_01693_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33144_ (_01695_, _01693_, _01692_);
  and _33145_ (_26891_[10], _01695_, _22762_);
  not _33146_ (_01697_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _33147_ (_01698_, _01681_, _01697_);
  and _33148_ (_01699_, _01698_, _01577_);
  nor _33149_ (_01700_, _01682_, _01697_);
  nor _33150_ (_01701_, _01700_, _01699_);
  not _33151_ (_01702_, _01701_);
  and _33152_ (_01703_, _01702_, _01685_);
  or _33153_ (_01704_, _01702_, _01685_);
  nand _33154_ (_01705_, _01704_, _25728_);
  nor _33155_ (_01706_, _01705_, _01703_);
  nor _33156_ (_01707_, _25728_, _23270_);
  or _33157_ (_01708_, _01707_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33158_ (_01709_, _01708_, _01706_);
  or _33159_ (_01710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _01532_);
  and _33160_ (_01711_, _01710_, _22762_);
  and _33161_ (_26891_[11], _01711_, _01709_);
  not _33162_ (_01712_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _33163_ (_01713_, _01699_, _01712_);
  and _33164_ (_01714_, _01698_, _01712_);
  and _33165_ (_01715_, _01714_, _01577_);
  nor _33166_ (_01717_, _01715_, _01713_);
  not _33167_ (_01718_, _01717_);
  or _33168_ (_01719_, _01718_, _01703_);
  and _33169_ (_01720_, _01718_, _01703_);
  nor _33170_ (_01721_, _01720_, _25729_);
  and _33171_ (_01722_, _01721_, _01719_);
  nor _33172_ (_01723_, _25728_, _23222_);
  or _33173_ (_01724_, _01723_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _33174_ (_01725_, _01724_, _01722_);
  or _33175_ (_01726_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _01532_);
  and _33176_ (_01727_, _01726_, _22762_);
  and _33177_ (_26891_[12], _01727_, _01725_);
  not _33178_ (_01728_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _33179_ (_01729_, _01715_, _01728_);
  and _33180_ (_01730_, _01715_, _01728_);
  nor _33181_ (_01731_, _01730_, _01729_);
  not _33182_ (_01732_, _01731_);
  and _33183_ (_01733_, _01732_, _01720_);
  nor _33184_ (_01734_, _01732_, _01720_);
  nor _33185_ (_01735_, _01734_, _01733_);
  or _33186_ (_01736_, _01735_, _25729_);
  or _33187_ (_01737_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _33188_ (_01738_, _01737_, _01532_);
  and _33189_ (_01739_, _01738_, _01736_);
  and _33190_ (_01740_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _33191_ (_01741_, _01740_, _01739_);
  and _33192_ (_26891_[13], _01741_, _22762_);
  not _33193_ (_01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _33194_ (_01743_, _01730_, _01742_);
  and _33195_ (_01744_, _01730_, _01742_);
  nor _33196_ (_01745_, _01744_, _01743_);
  not _33197_ (_01746_, _01745_);
  and _33198_ (_01747_, _01746_, _01733_);
  nor _33199_ (_01748_, _01746_, _01733_);
  nor _33200_ (_01749_, _01748_, _01747_);
  or _33201_ (_01751_, _01749_, _25729_);
  or _33202_ (_01752_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _33203_ (_01753_, _01752_, _01532_);
  and _33204_ (_01754_, _01753_, _01751_);
  and _33205_ (_01755_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _33206_ (_01756_, _01755_, _01754_);
  and _33207_ (_26891_[14], _01756_, _22762_);
  nand _33208_ (_01757_, _23074_, _22946_);
  and _33209_ (_01758_, _23661_, _01757_);
  and _33210_ (_01759_, _01758_, _24275_);
  and _33211_ (_01760_, _01759_, _23946_);
  not _33212_ (_01762_, _01759_);
  and _33213_ (_01763_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or _33214_ (_22631_, _01763_, _01760_);
  and _33215_ (_01764_, _01759_, _23649_);
  and _33216_ (_01765_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or _33217_ (_22632_, _01765_, _01764_);
  nor _33218_ (_01766_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _33219_ (_01767_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _33220_ (_01768_, _01767_, _01766_);
  nor _33221_ (_01769_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor _33222_ (_01770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _33223_ (_01771_, _01770_, _01769_);
  and _33224_ (_01772_, _01771_, _01768_);
  and _33225_ (_01773_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _33226_ (_01774_, _01773_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _33227_ (_26895_[0], _01774_, _22762_);
  and _33228_ (_01775_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _33229_ (_01776_, _01775_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _33230_ (_26895_[1], _01776_, _22762_);
  and _33231_ (_01777_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or _33232_ (_01778_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _33233_ (_26895_[2], _01778_, _22762_);
  and _33234_ (_01779_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _33235_ (_01781_, _01779_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _33236_ (_26895_[3], _01781_, _22762_);
  and _33237_ (_01782_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _33238_ (_01783_, _01782_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _33239_ (_26895_[4], _01783_, _22762_);
  and _33240_ (_01785_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _33241_ (_01786_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _33242_ (_26895_[5], _01786_, _22762_);
  and _33243_ (_01787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22762_);
  and _33244_ (_01788_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _22762_);
  and _33245_ (_01790_, _01788_, _01772_);
  or _33246_ (_26895_[6], _01790_, _01787_);
  nor _33247_ (_01791_, _01518_, _23950_);
  nand _33248_ (_01792_, _01791_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _33249_ (_01793_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  or _33250_ (_01794_, _01791_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _33251_ (_01795_, _01794_, _01793_);
  and _33252_ (_26896_[0], _01795_, _01792_);
  not _33253_ (_01796_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _33254_ (_01797_, _01518_, _01796_);
  or _33255_ (_01798_, _01505_, _23855_);
  nand _33256_ (_01799_, _01505_, _23855_);
  and _33257_ (_01800_, _01799_, _01798_);
  nand _33258_ (_01801_, _01800_, _01797_);
  or _33259_ (_01802_, _01800_, _01797_);
  and _33260_ (_01803_, _01802_, _01801_);
  or _33261_ (_01804_, _01803_, _23950_);
  or _33262_ (_01805_, _22768_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _33263_ (_01807_, _01805_, _01793_);
  and _33264_ (_26896_[1], _01807_, _01804_);
  and _33265_ (_01808_, _23901_, _23068_);
  and _33266_ (_01809_, _23905_, _23662_);
  and _33267_ (_01810_, _01809_, _01808_);
  and _33268_ (_01811_, _01810_, _23747_);
  not _33269_ (_01812_, _01810_);
  and _33270_ (_01813_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or _33271_ (_22633_, _01813_, _01811_);
  and _33272_ (_22634_, t0_i, _22762_);
  and _33273_ (_01814_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _23978_);
  and _33274_ (_01815_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33275_ (_01816_, _01815_, _01814_);
  and _33276_ (_26899_[0], _01816_, _22762_);
  and _33277_ (_01817_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _23978_);
  and _33278_ (_01818_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33279_ (_01819_, _01818_, _01817_);
  and _33280_ (_26899_[1], _01819_, _22762_);
  and _33281_ (_01821_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _23978_);
  and _33282_ (_01822_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33283_ (_01823_, _01822_, _01821_);
  and _33284_ (_26899_[2], _01823_, _22762_);
  and _33285_ (_01824_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _23978_);
  and _33286_ (_01825_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33287_ (_01826_, _01825_, _01824_);
  and _33288_ (_26899_[3], _01826_, _22762_);
  and _33289_ (_01827_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _23978_);
  and _33290_ (_01828_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33291_ (_01829_, _01828_, _01827_);
  and _33292_ (_26899_[4], _01829_, _22762_);
  and _33293_ (_01830_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _23978_);
  and _33294_ (_01831_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33295_ (_01832_, _01831_, _01830_);
  and _33296_ (_26899_[5], _01832_, _22762_);
  and _33297_ (_01834_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _23978_);
  and _33298_ (_01835_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _33299_ (_01836_, _01835_, _01834_);
  and _33300_ (_26899_[6], _01836_, _22762_);
  and _33301_ (_26902_[0], _23968_, _22762_);
  nor _33302_ (_26902_[1], _23973_, rst);
  and _33303_ (_26902_[2], _23976_, _22762_);
  and _33304_ (_01838_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor _33305_ (_01839_, _23953_, _25783_);
  or _33306_ (_01840_, _01839_, _01838_);
  and _33307_ (_26904_[0], _01840_, _22762_);
  and _33308_ (_01841_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor _33309_ (_01842_, _23953_, _25788_);
  or _33310_ (_01843_, _01842_, _01841_);
  and _33311_ (_26904_[1], _01843_, _22762_);
  and _33312_ (_01844_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor _33313_ (_01845_, _23953_, _25793_);
  or _33314_ (_01846_, _01845_, _01844_);
  and _33315_ (_26904_[2], _01846_, _22762_);
  and _33316_ (_01847_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor _33317_ (_01848_, _23953_, _25798_);
  or _33318_ (_01849_, _01848_, _01847_);
  and _33319_ (_26904_[3], _01849_, _22762_);
  and _33320_ (_01850_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor _33321_ (_01851_, _23953_, _25803_);
  or _33322_ (_01852_, _01851_, _01850_);
  and _33323_ (_26904_[4], _01852_, _22762_);
  and _33324_ (_01853_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor _33325_ (_01854_, _23953_, _25807_);
  or _33326_ (_01855_, _01854_, _01853_);
  and _33327_ (_26904_[5], _01855_, _22762_);
  and _33328_ (_01856_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor _33329_ (_01857_, _23953_, _25811_);
  or _33330_ (_01858_, _01857_, _01856_);
  and _33331_ (_26904_[6], _01858_, _22762_);
  and _33332_ (_01859_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor _33333_ (_01861_, _23953_, _25817_);
  or _33334_ (_01862_, _01861_, _01859_);
  and _33335_ (_26904_[7], _01862_, _22762_);
  and _33336_ (_01863_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _33337_ (_01864_, _23953_, _25822_);
  or _33338_ (_01865_, _01864_, _01863_);
  and _33339_ (_26904_[8], _01865_, _22762_);
  and _33340_ (_01867_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _33341_ (_01868_, _23953_, _25826_);
  or _33342_ (_01869_, _01868_, _01867_);
  and _33343_ (_26904_[9], _01869_, _22762_);
  and _33344_ (_01870_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _33345_ (_01871_, _23953_, _25830_);
  or _33346_ (_01872_, _01871_, _01870_);
  and _33347_ (_26904_[10], _01872_, _22762_);
  and _33348_ (_01873_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _33349_ (_01874_, _23953_, _25834_);
  or _33350_ (_01875_, _01874_, _01873_);
  and _33351_ (_26904_[11], _01875_, _22762_);
  and _33352_ (_01876_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _33353_ (_01877_, _23953_, _25838_);
  or _33354_ (_01879_, _01877_, _01876_);
  and _33355_ (_26904_[12], _01879_, _22762_);
  and _33356_ (_01880_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _33357_ (_01882_, _23953_, _25842_);
  or _33358_ (_01883_, _01882_, _01880_);
  and _33359_ (_26904_[13], _01883_, _22762_);
  and _33360_ (_01884_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _33361_ (_01886_, _23953_, _25846_);
  or _33362_ (_01887_, _01886_, _01884_);
  and _33363_ (_26904_[14], _01887_, _22762_);
  and _33364_ (_01888_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _33365_ (_01889_, _23953_, _25850_);
  or _33366_ (_01890_, _01889_, _01888_);
  and _33367_ (_26904_[15], _01890_, _22762_);
  and _33368_ (_01891_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _33369_ (_01892_, _23953_, _25854_);
  or _33370_ (_01893_, _01892_, _01891_);
  and _33371_ (_26904_[16], _01893_, _22762_);
  and _33372_ (_01894_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _33373_ (_01895_, _23953_, _25858_);
  or _33374_ (_01896_, _01895_, _01894_);
  and _33375_ (_26904_[17], _01896_, _22762_);
  and _33376_ (_01897_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _33377_ (_01898_, _23953_, _25862_);
  or _33378_ (_01899_, _01898_, _01897_);
  and _33379_ (_26904_[18], _01899_, _22762_);
  and _33380_ (_01900_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _33381_ (_01902_, _23953_, _25866_);
  or _33382_ (_01903_, _01902_, _01900_);
  and _33383_ (_26904_[19], _01903_, _22762_);
  and _33384_ (_01904_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _33385_ (_01905_, _23953_, _25870_);
  or _33386_ (_01906_, _01905_, _01904_);
  and _33387_ (_26904_[20], _01906_, _22762_);
  and _33388_ (_01907_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _33389_ (_01908_, _23953_, _25876_);
  or _33390_ (_01909_, _01908_, _01907_);
  and _33391_ (_26904_[21], _01909_, _22762_);
  and _33392_ (_01910_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _33393_ (_01911_, _23953_, _25880_);
  or _33394_ (_01912_, _01911_, _01910_);
  and _33395_ (_26904_[22], _01912_, _22762_);
  and _33396_ (_01913_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _33397_ (_01914_, _23953_, _25884_);
  or _33398_ (_01915_, _01914_, _01913_);
  and _33399_ (_26904_[23], _01915_, _22762_);
  and _33400_ (_01916_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and _33401_ (_01917_, _25888_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or _33402_ (_01918_, _01917_, _01916_);
  and _33403_ (_26904_[24], _01918_, _22762_);
  and _33404_ (_01919_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _33405_ (_01920_, _23953_, _25892_);
  or _33406_ (_01921_, _01920_, _01919_);
  and _33407_ (_26904_[25], _01921_, _22762_);
  and _33408_ (_01922_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _33409_ (_01923_, _23953_, _25896_);
  or _33410_ (_01924_, _01923_, _01922_);
  and _33411_ (_26904_[26], _01924_, _22762_);
  and _33412_ (_01925_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _33413_ (_01926_, _23953_, _25900_);
  or _33414_ (_01927_, _01926_, _01925_);
  and _33415_ (_26904_[27], _01927_, _22762_);
  and _33416_ (_01929_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _33417_ (_01930_, _23953_, _25904_);
  or _33418_ (_01931_, _01930_, _01929_);
  and _33419_ (_26904_[28], _01931_, _22762_);
  and _33420_ (_01932_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _33421_ (_01934_, _23953_, _25908_);
  or _33422_ (_01935_, _01934_, _01932_);
  and _33423_ (_26904_[29], _01935_, _22762_);
  and _33424_ (_01936_, _23953_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _33425_ (_01937_, _23953_, _25912_);
  or _33426_ (_01938_, _01937_, _01936_);
  and _33427_ (_26904_[30], _01938_, _22762_);
  and _33428_ (_01939_, _01759_, _23707_);
  and _33429_ (_01940_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or _33430_ (_22635_, _01940_, _01939_);
  and _33431_ (_01941_, _25733_, _23946_);
  and _33432_ (_01942_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or _33433_ (_22636_, _01942_, _01941_);
  and _33434_ (_01944_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and _33435_ (_01945_, _25763_, _23898_);
  or _33436_ (_22637_, _01945_, _01944_);
  and _33437_ (_01947_, _25733_, _24050_);
  and _33438_ (_01948_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or _33439_ (_22638_, _01948_, _01947_);
  and _33440_ (_01949_, _25733_, _23747_);
  and _33441_ (_01950_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or _33442_ (_22639_, _01950_, _01949_);
  and _33443_ (_01951_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and _33444_ (_01952_, _25763_, _23778_);
  or _33445_ (_22640_, _01952_, _01951_);
  not _33446_ (_01954_, _24096_);
  or _33447_ (_01955_, _26565_, _01954_);
  or _33448_ (_01956_, _24096_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _33449_ (_01957_, _01956_, _22762_);
  and _33450_ (_26908_[0], _01957_, _01955_);
  nand _33451_ (_01958_, _00372_, _24096_);
  or _33452_ (_01959_, _24096_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _33453_ (_01960_, _01959_, _22762_);
  and _33454_ (_26908_[1], _01960_, _01958_);
  or _33455_ (_01961_, _00451_, _01954_);
  or _33456_ (_01962_, _24096_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _33457_ (_01963_, _01962_, _22762_);
  and _33458_ (_26908_[2], _01963_, _01961_);
  or _33459_ (_01964_, _00545_, _01954_);
  or _33460_ (_01965_, _24096_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _33461_ (_01966_, _01965_, _22762_);
  and _33462_ (_26908_[3], _01966_, _01964_);
  and _33463_ (_01967_, _25078_, _24201_);
  not _33464_ (_01968_, _01967_);
  and _33465_ (_01969_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and _33466_ (_01970_, _01967_, _24050_);
  or _33467_ (_22641_, _01970_, _01969_);
  and _33468_ (_01971_, _24329_, _23664_);
  and _33469_ (_01972_, _01971_, _23778_);
  not _33470_ (_01973_, _01971_);
  and _33471_ (_01974_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or _33472_ (_22642_, _01974_, _01972_);
  and _33473_ (_01975_, _24063_, _23662_);
  and _33474_ (_01977_, _01975_, _24297_);
  and _33475_ (_01978_, _01975_, _24126_);
  nor _33476_ (_01979_, _01978_, _01977_);
  or _33477_ (_01980_, _01979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _33478_ (_01981_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _33479_ (_01982_, _01981_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _33480_ (_01983_, _01982_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _33481_ (_01984_, _01983_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _33482_ (_01985_, _01984_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _33483_ (_01986_, _01985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _33484_ (_01987_, _01986_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _33485_ (_01988_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _33486_ (_01989_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _33487_ (_01990_, _01989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _33488_ (_01992_, _01990_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _33489_ (_01993_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _33490_ (_01994_, _01993_, _01992_);
  and _33491_ (_01995_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _33492_ (_01996_, _01995_, _01994_);
  not _33493_ (_01997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nor _33494_ (_01998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _33495_ (_01999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _33496_ (_02000_, _01999_, _01998_);
  and _33497_ (_02001_, _02000_, _01997_);
  not _33498_ (_02002_, _02001_);
  or _33499_ (_02004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _33500_ (_02005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _33501_ (_02006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _02005_);
  and _33502_ (_02007_, _02006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _33503_ (_02009_, _02007_, _02004_);
  and _33504_ (_02010_, _02009_, _01998_);
  and _33505_ (_02011_, _02010_, _02002_);
  nand _33506_ (_02012_, _02011_, _01996_);
  nand _33507_ (_02014_, _02012_, _01979_);
  and _33508_ (_02015_, _02014_, _22762_);
  and _33509_ (_22644_, _02015_, _01980_);
  nand _33510_ (_02016_, _01978_, _23702_);
  not _33511_ (_02017_, _01977_);
  and _33512_ (_02018_, _02009_, _01994_);
  and _33513_ (_02019_, _02018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _33514_ (_02020_, _02019_, _02001_);
  and _33515_ (_02021_, _02020_, _02017_);
  or _33516_ (_02022_, _02021_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _33517_ (_02023_, _02019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _33518_ (_02024_, _02023_, _02002_);
  and _33519_ (_02025_, _01998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not _33520_ (_02026_, _02025_);
  and _33521_ (_02027_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or _33522_ (_02028_, _02027_, _01977_);
  or _33523_ (_02029_, _02028_, _02024_);
  and _33524_ (_02030_, _02029_, _02022_);
  or _33525_ (_02031_, _02030_, _01978_);
  and _33526_ (_02032_, _02031_, _22762_);
  and _33527_ (_22645_, _02032_, _02016_);
  and _33528_ (_02034_, _24655_, _24064_);
  or _33529_ (_02035_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _33530_ (_02036_, _02035_, _22762_);
  not _33531_ (_02037_, _02034_);
  or _33532_ (_02038_, _02037_, _23816_);
  and _33533_ (_22646_, _02038_, _02036_);
  nor _33534_ (_02039_, _02017_, _23702_);
  and _33535_ (_02040_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _33536_ (_02041_, _02009_, _01996_);
  and _33537_ (_02042_, _02041_, _02040_);
  and _33538_ (_02043_, _02009_, _01986_);
  or _33539_ (_02044_, _02043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand _33540_ (_02045_, _02043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _33541_ (_02046_, _02045_, _02044_);
  or _33542_ (_02047_, _02046_, _02001_);
  or _33543_ (_02048_, _02047_, _02042_);
  or _33544_ (_02049_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _33545_ (_02050_, _02049_, _01979_);
  and _33546_ (_02051_, _02050_, _02048_);
  and _33547_ (_02052_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _33548_ (_02053_, _02052_, _02051_);
  or _33549_ (_02054_, _02053_, _02039_);
  and _33550_ (_22647_, _02054_, _22762_);
  not _33551_ (_02055_, _01998_);
  and _33552_ (_02056_, _02009_, _02055_);
  and _33553_ (_02057_, _02056_, _01979_);
  or _33554_ (_02058_, _02057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _33555_ (_02059_, _01996_);
  nand _33556_ (_02061_, _02057_, _02059_);
  and _33557_ (_02063_, _02061_, _22762_);
  and _33558_ (_22648_, _02063_, _02058_);
  nor _33559_ (_02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and _33560_ (_02065_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and _33561_ (_02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _22762_);
  and _33562_ (_02067_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or _33563_ (_22649_, _02067_, _02065_);
  and _33564_ (_02069_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and _33565_ (_02070_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or _33566_ (_22650_, _02070_, _02069_);
  and _33567_ (_02071_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _33568_ (_02072_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _33569_ (_22651_, _02072_, _02071_);
  and _33570_ (_02073_, _01975_, _24119_);
  nand _33571_ (_02074_, _02073_, _23702_);
  and _33572_ (_02075_, _02025_, _01999_);
  not _33573_ (_02076_, _02075_);
  and _33574_ (_02077_, _01975_, _24292_);
  nor _33575_ (_02078_, _02077_, _02076_);
  not _33576_ (_02079_, _02078_);
  and _33577_ (_02080_, _02079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _33578_ (_02081_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _33579_ (_02082_, _02081_, _02080_);
  or _33580_ (_02083_, _02082_, _02073_);
  and _33581_ (_02084_, _02083_, _22762_);
  and _33582_ (_22652_, _02084_, _02074_);
  and _33583_ (_22653_, t2ex_i, _22762_);
  nand _33584_ (_02086_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _22762_);
  nor _33585_ (_22654_, _02086_, t2_i);
  and _33586_ (_22655_, t2_i, _22762_);
  and _33587_ (_02087_, _01758_, _23991_);
  and _33588_ (_02088_, _02087_, _23707_);
  not _33589_ (_02089_, _02087_);
  and _33590_ (_02090_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or _33591_ (_22656_, _02090_, _02088_);
  and _33592_ (_02091_, _24173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and _33593_ (_02092_, _24177_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or _33594_ (_02093_, _02092_, _24257_);
  and _33595_ (_02094_, _02093_, _24255_);
  or _33596_ (_02095_, _02092_, _24243_);
  and _33597_ (_02096_, _02095_, _24132_);
  and _33598_ (_02097_, _25584_, _24145_);
  or _33599_ (_02099_, _02097_, _02092_);
  and _33600_ (_02100_, _02099_, _24184_);
  or _33601_ (_02101_, _02100_, _02096_);
  or _33602_ (_02102_, _02101_, _02094_);
  or _33603_ (_02103_, _02102_, _02091_);
  and _33604_ (_02104_, _02103_, _24128_);
  and _33605_ (_22657_, _02104_, _24166_);
  and _33606_ (_02105_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and _33607_ (_02106_, _25763_, _23824_);
  or _33608_ (_22658_, _02106_, _02105_);
  and _33609_ (_02107_, _24356_, _23069_);
  and _33610_ (_02108_, _02107_, _23649_);
  not _33611_ (_02109_, _02107_);
  and _33612_ (_02110_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  or _33613_ (_22659_, _02110_, _02108_);
  and _33614_ (_02111_, _23790_, _23707_);
  and _33615_ (_02112_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or _33616_ (_22660_, _02112_, _02111_);
  and _33617_ (_02113_, _01759_, _23778_);
  and _33618_ (_02114_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or _33619_ (_22661_, _02114_, _02113_);
  and _33620_ (_02115_, _01759_, _23824_);
  and _33621_ (_02116_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or _33622_ (_22662_, _02116_, _02115_);
  and _33623_ (_22663_, _01787_, _24862_);
  and _33624_ (_02117_, _24862_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _33625_ (_02118_, _02117_, _24951_);
  and _33626_ (_22664_, _02118_, _22762_);
  or _33627_ (_02119_, _25057_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _33628_ (_02120_, _02119_, _25056_);
  and _33629_ (_02121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _24865_);
  nand _33630_ (_02122_, _02121_, _24904_);
  nand _33631_ (_02123_, _02122_, _24913_);
  or _33632_ (_02124_, _02123_, _02120_);
  or _33633_ (_02125_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _33634_ (_02126_, _02125_, _24913_);
  and _33635_ (_02127_, _02126_, _24908_);
  and _33636_ (_02128_, _02127_, _02124_);
  and _33637_ (_02129_, _02121_, _24907_);
  or _33638_ (_02130_, _02129_, _02128_);
  and _33639_ (_02131_, _02130_, _24949_);
  nand _33640_ (_02132_, _24917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nand _33641_ (_02133_, _02132_, _25004_);
  or _33642_ (_02134_, _02133_, _02131_);
  or _33643_ (_02135_, _24954_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _33644_ (_02136_, _02135_, _22762_);
  not _33645_ (_02137_, _24895_);
  nor _33646_ (_02138_, _02121_, _02137_);
  nor _33647_ (_02139_, _02138_, _25136_);
  or _33648_ (_02140_, _25041_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _33649_ (_02141_, _02140_, _25044_);
  nand _33650_ (_02142_, _02121_, _24891_);
  nand _33651_ (_02143_, _02142_, _24888_);
  or _33652_ (_02144_, _02143_, _02141_);
  or _33653_ (_02145_, _02125_, _24888_);
  and _33654_ (_02146_, _02145_, _24883_);
  and _33655_ (_02147_, _02146_, _02144_);
  or _33656_ (_02148_, _02147_, _24862_);
  or _33657_ (_02149_, _02148_, _02139_);
  and _33658_ (_02150_, _02149_, _02136_);
  and _33659_ (_22665_, _02150_, _02134_);
  or _33660_ (_02151_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _24865_);
  or _33661_ (_02152_, _02151_, _24913_);
  and _33662_ (_02153_, _02152_, _24908_);
  or _33663_ (_02154_, _24980_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _33664_ (_02155_, _02154_, _24979_);
  and _33665_ (_02156_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _33666_ (_02157_, _02156_, _24904_);
  nand _33667_ (_02158_, _02157_, _24913_);
  or _33668_ (_02159_, _02158_, _02155_);
  and _33669_ (_02160_, _02159_, _02153_);
  and _33670_ (_02161_, _02156_, _24907_);
  or _33671_ (_02162_, _02161_, _02160_);
  and _33672_ (_02163_, _02162_, _24949_);
  nand _33673_ (_02164_, _24917_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nand _33674_ (_02165_, _02164_, _25004_);
  or _33675_ (_02166_, _02165_, _02163_);
  or _33676_ (_02167_, _24954_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _33677_ (_02168_, _02167_, _22762_);
  nor _33678_ (_02169_, _02156_, _02137_);
  nor _33679_ (_02170_, _02169_, _25136_);
  or _33680_ (_02171_, _24958_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _33681_ (_02172_, _02171_, _24956_);
  nand _33682_ (_02173_, _02156_, _24891_);
  nand _33683_ (_02174_, _02173_, _24888_);
  or _33684_ (_02175_, _02174_, _02172_);
  or _33685_ (_02176_, _02151_, _24888_);
  and _33686_ (_02177_, _02176_, _24883_);
  and _33687_ (_02178_, _02177_, _02175_);
  or _33688_ (_02179_, _02178_, _24862_);
  or _33689_ (_02180_, _02179_, _02170_);
  and _33690_ (_02181_, _02180_, _02168_);
  and _33691_ (_22666_, _02181_, _02166_);
  and _33692_ (_02182_, _24730_, _24125_);
  nand _33693_ (_02183_, _02182_, _23594_);
  or _33694_ (_02184_, _02182_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _33695_ (_02185_, _02184_, _24737_);
  and _33696_ (_02186_, _02185_, _02183_);
  and _33697_ (_02187_, _24736_, _23939_);
  or _33698_ (_02188_, _02187_, _02186_);
  and _33699_ (_22667_, _02188_, _22762_);
  and _33700_ (_02189_, _24648_, _24296_);
  nand _33701_ (_02190_, _02189_, _23594_);
  or _33702_ (_02191_, _02189_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _33703_ (_02192_, _02191_, _24659_);
  and _33704_ (_02193_, _02192_, _02190_);
  and _33705_ (_02194_, _24658_, _23642_);
  or _33706_ (_02195_, _02194_, _02193_);
  and _33707_ (_22668_, _02195_, _22762_);
  and _33708_ (_02196_, _01759_, _23898_);
  and _33709_ (_02197_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or _33710_ (_22669_, _02197_, _02196_);
  and _33711_ (_02198_, _23707_, _23077_);
  and _33712_ (_02199_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  or _33713_ (_22670_, _02199_, _02198_);
  and _33714_ (_02200_, _24356_, _23986_);
  and _33715_ (_02201_, _02200_, _23898_);
  not _33716_ (_02202_, _02200_);
  and _33717_ (_02203_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or _33718_ (_22671_, _02203_, _02201_);
  and _33719_ (_02204_, _24766_, _23986_);
  not _33720_ (_02205_, _02204_);
  and _33721_ (_02206_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and _33722_ (_02207_, _02204_, _23747_);
  or _33723_ (_22672_, _02207_, _02206_);
  and _33724_ (_02208_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and _33725_ (_02209_, _02204_, _23649_);
  or _33726_ (_27039_, _02209_, _02208_);
  and _33727_ (_02211_, _02087_, _23778_);
  and _33728_ (_02212_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or _33729_ (_27008_, _02212_, _02211_);
  and _33730_ (_02213_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and _33731_ (_02214_, _02204_, _23824_);
  or _33732_ (_27038_, _02214_, _02213_);
  and _33733_ (_02215_, _01758_, _23903_);
  and _33734_ (_02216_, _02215_, _23707_);
  not _33735_ (_02217_, _02215_);
  and _33736_ (_02218_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or _33737_ (_22673_, _02218_, _02216_);
  nor _33738_ (_26897_[2], _00470_, rst);
  nor _33739_ (_26887_[5], _00006_, rst);
  and _33740_ (_02219_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and _33741_ (_02220_, _02204_, _24050_);
  or _33742_ (_22674_, _02220_, _02219_);
  and _33743_ (_02221_, _02087_, _23898_);
  and _33744_ (_02222_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or _33745_ (_22675_, _02222_, _02221_);
  and _33746_ (_02223_, _02087_, _23747_);
  and _33747_ (_02224_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or _33748_ (_22676_, _02224_, _02223_);
  and _33749_ (_02225_, _02087_, _23824_);
  and _33750_ (_02226_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or _33751_ (_22677_, _02226_, _02225_);
  and _33752_ (_02227_, _24331_, _23707_);
  and _33753_ (_02228_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or _33754_ (_22678_, _02228_, _02227_);
  and _33755_ (_02229_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and _33756_ (_02230_, _02204_, _23946_);
  or _33757_ (_27040_, _02230_, _02229_);
  nor _33758_ (_26860_[0], _24402_, rst);
  nor _33759_ (_26860_[6], _24486_, rst);
  and _33760_ (_02231_, _24852_, _23707_);
  and _33761_ (_02232_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  or _33762_ (_22679_, _02232_, _02231_);
  and _33763_ (_02233_, _24006_, _23946_);
  and _33764_ (_02234_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or _33765_ (_22680_, _02234_, _02233_);
  and _33766_ (_02235_, _02215_, _23778_);
  and _33767_ (_02236_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or _33768_ (_22681_, _02236_, _02235_);
  and _33769_ (_02237_, _02215_, _23824_);
  and _33770_ (_02238_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or _33771_ (_22682_, _02238_, _02237_);
  and _33772_ (_02239_, _02215_, _23898_);
  and _33773_ (_02240_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or _33774_ (_22683_, _02240_, _02239_);
  and _33775_ (_02241_, _24275_, _23789_);
  and _33776_ (_02242_, _02241_, _23747_);
  not _33777_ (_02243_, _02241_);
  and _33778_ (_02244_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or _33779_ (_27293_, _02244_, _02242_);
  and _33780_ (_02245_, _24766_, _23069_);
  not _33781_ (_02246_, _02245_);
  and _33782_ (_02247_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  and _33783_ (_02248_, _02245_, _23707_);
  or _33784_ (_27037_, _02248_, _02247_);
  and _33785_ (_02249_, _24050_, _23077_);
  and _33786_ (_02250_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  or _33787_ (_22684_, _02250_, _02249_);
  and _33788_ (_02251_, _23946_, _23077_);
  and _33789_ (_02252_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  or _33790_ (_22685_, _02252_, _02251_);
  and _33791_ (_02253_, _25618_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _33792_ (_02254_, _24596_, _24539_);
  or _33793_ (_02255_, _02254_, _24585_);
  and _33794_ (_02256_, _24556_, _24546_);
  or _33795_ (_02257_, _02256_, _25640_);
  and _33796_ (_02258_, _24613_, _26650_);
  or _33797_ (_02259_, _02258_, _26666_);
  and _33798_ (_02260_, _24613_, _24604_);
  and _33799_ (_02261_, _26625_, _24582_);
  and _33800_ (_02262_, _26625_, _24540_);
  or _33801_ (_02263_, _02262_, _02261_);
  or _33802_ (_02264_, _02263_, _02260_);
  or _33803_ (_02265_, _02264_, _26591_);
  or _33804_ (_02266_, _02265_, _02259_);
  and _33805_ (_02267_, _26650_, _26582_);
  and _33806_ (_02268_, _24567_, _24546_);
  or _33807_ (_02269_, _02268_, _02267_);
  and _33808_ (_02270_, _24604_, _24556_);
  and _33809_ (_02271_, _24593_, _24556_);
  or _33810_ (_02272_, _02271_, _02270_);
  and _33811_ (_02273_, _24606_, _24556_);
  and _33812_ (_02274_, _24589_, _24556_);
  or _33813_ (_02275_, _02274_, _02273_);
  or _33814_ (_02276_, _02275_, _02272_);
  or _33815_ (_02277_, _02276_, _02269_);
  or _33816_ (_02278_, _02277_, _02266_);
  or _33817_ (_02279_, _02278_, _02257_);
  or _33818_ (_02280_, _02279_, _02255_);
  and _33819_ (_02281_, _02280_, _25644_);
  or _33820_ (_26867_[0], _02281_, _02253_);
  and _33821_ (_02282_, _24283_, _23898_);
  and _33822_ (_02283_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  or _33823_ (_22686_, _02283_, _02282_);
  and _33824_ (_02284_, _01809_, _24329_);
  and _33825_ (_02285_, _02284_, _24050_);
  not _33826_ (_02286_, _02284_);
  and _33827_ (_02287_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  or _33828_ (_22687_, _02287_, _02285_);
  and _33829_ (_02288_, _02284_, _23649_);
  and _33830_ (_02289_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  or _33831_ (_22688_, _02289_, _02288_);
  and _33832_ (_02290_, _02284_, _23747_);
  and _33833_ (_02291_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  or _33834_ (_22689_, _02291_, _02290_);
  and _33835_ (_02292_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and _33836_ (_02293_, _24692_, _24050_);
  or _33837_ (_22690_, _02293_, _02292_);
  and _33838_ (_02294_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and _33839_ (_02295_, _24692_, _23707_);
  or _33840_ (_27236_, _02295_, _02294_);
  and _33841_ (_02296_, _02284_, _23778_);
  and _33842_ (_02297_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  or _33843_ (_27115_, _02297_, _02296_);
  and _33844_ (_02298_, _24201_, _23752_);
  not _33845_ (_02299_, _02298_);
  and _33846_ (_02300_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  and _33847_ (_02301_, _02298_, _23778_);
  or _33848_ (_22691_, _02301_, _02300_);
  and _33849_ (_02302_, _01809_, _23752_);
  and _33850_ (_02303_, _02302_, _23707_);
  not _33851_ (_02304_, _02302_);
  and _33852_ (_02305_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or _33853_ (_22692_, _02305_, _02303_);
  and _33854_ (_02306_, _24201_, _23069_);
  not _33855_ (_02307_, _02306_);
  and _33856_ (_02308_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  and _33857_ (_02309_, _02306_, _23824_);
  or _33858_ (_22693_, _02309_, _02308_);
  and _33859_ (_02310_, _24678_, _23003_);
  and _33860_ (_02311_, _25769_, _23073_);
  and _33861_ (_02312_, _02311_, _02310_);
  and _33862_ (_02313_, _02312_, _25926_);
  and _33863_ (_02314_, _02313_, _24043_);
  not _33864_ (_02315_, _02313_);
  and _33865_ (_02316_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or _33866_ (_22694_, _02316_, _02314_);
  and _33867_ (_02317_, _02302_, _23946_);
  and _33868_ (_02318_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or _33869_ (_22695_, _02318_, _02317_);
  and _33870_ (_02319_, _02302_, _23747_);
  and _33871_ (_02320_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or _33872_ (_22696_, _02320_, _02319_);
  and _33873_ (_02321_, _24356_, _23752_);
  and _33874_ (_02322_, _02321_, _23649_);
  not _33875_ (_02323_, _02321_);
  and _33876_ (_02324_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  or _33877_ (_22697_, _02324_, _02322_);
  and _33878_ (_02325_, _23662_, _23072_);
  and _33879_ (_02326_, _02325_, _24329_);
  and _33880_ (_02327_, _02326_, _23778_);
  not _33881_ (_02328_, _02326_);
  and _33882_ (_02329_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or _33883_ (_22698_, _02329_, _02327_);
  and _33884_ (_02330_, _02302_, _23898_);
  and _33885_ (_02331_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or _33886_ (_22699_, _02331_, _02330_);
  and _33887_ (_02332_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and _33888_ (_02333_, _24692_, _23649_);
  or _33889_ (_27235_, _02333_, _02332_);
  and _33890_ (_02334_, _02215_, _23946_);
  and _33891_ (_02335_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or _33892_ (_26992_, _02335_, _02334_);
  and _33893_ (_02336_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and _33894_ (_02337_, _02204_, _23778_);
  or _33895_ (_22700_, _02337_, _02336_);
  and _33896_ (_02339_, _02215_, _23649_);
  and _33897_ (_02340_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or _33898_ (_22701_, _02340_, _02339_);
  nor _33899_ (_26887_[0], _00129_, rst);
  and _33900_ (_02341_, _25748_, _23824_);
  and _33901_ (_02342_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or _33902_ (_22702_, _02342_, _02341_);
  and _33903_ (_02343_, _02215_, _23747_);
  and _33904_ (_02344_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or _33905_ (_22703_, _02344_, _02343_);
  and _33906_ (_02345_, _01808_, _24370_);
  and _33907_ (_02346_, _02345_, _23778_);
  not _33908_ (_02347_, _02345_);
  and _33909_ (_02349_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or _33910_ (_22704_, _02349_, _02346_);
  and _33911_ (_02350_, _01758_, _24005_);
  and _33912_ (_02351_, _02350_, _23649_);
  not _33913_ (_02352_, _02350_);
  and _33914_ (_02353_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or _33915_ (_22705_, _02353_, _02351_);
  nor _33916_ (_02354_, _23596_, _26379_);
  and _33917_ (_02355_, _26385_, _23596_);
  or _33918_ (_02356_, _02355_, _02354_);
  and _33919_ (_22706_, _02356_, _22762_);
  and _33920_ (_02357_, _02200_, _23649_);
  and _33921_ (_02358_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or _33922_ (_27166_, _02358_, _02357_);
  and _33923_ (_02359_, _02325_, _01808_);
  and _33924_ (_02360_, _02359_, _24050_);
  not _33925_ (_02361_, _02359_);
  and _33926_ (_02363_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  or _33927_ (_27155_, _02363_, _02360_);
  and _33928_ (_02364_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and _33929_ (_02365_, _24692_, _23946_);
  or _33930_ (_22707_, _02365_, _02364_);
  and _33931_ (_02366_, _01971_, _23898_);
  and _33932_ (_02367_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  or _33933_ (_22708_, _02367_, _02366_);
  and _33934_ (_02368_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and _33935_ (_02369_, _24692_, _23747_);
  or _33936_ (_22709_, _02369_, _02368_);
  and _33937_ (_02370_, _24005_, _23754_);
  and _33938_ (_02371_, _02370_, _23898_);
  not _33939_ (_02372_, _02370_);
  and _33940_ (_02373_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or _33941_ (_22710_, _02373_, _02371_);
  and _33942_ (_02374_, _01809_, _23656_);
  and _33943_ (_02375_, _02374_, _24050_);
  not _33944_ (_02376_, _02374_);
  and _33945_ (_02377_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  or _33946_ (_22711_, _02377_, _02375_);
  nor _33947_ (_02378_, _26656_, _26668_);
  nand _33948_ (_02379_, _02378_, _26597_);
  or _33949_ (_02380_, _26644_, _26652_);
  or _33950_ (_02381_, _26660_, _26641_);
  or _33951_ (_02382_, _02381_, _26637_);
  or _33952_ (_02383_, _02382_, _02380_);
  or _33953_ (_02384_, _02383_, _02379_);
  and _33954_ (_02385_, _02384_, _26572_);
  and _33955_ (_02386_, _25629_, _24566_);
  nor _33956_ (_02387_, _02386_, _02385_);
  not _33957_ (_02388_, _02387_);
  nor _33958_ (_02389_, _02388_, _00099_);
  not _33959_ (_02390_, _02389_);
  or _33960_ (_02391_, _02387_, _26777_);
  or _33961_ (_02392_, _02391_, _00058_);
  and _33962_ (_02393_, _02392_, _02390_);
  and _33963_ (_02394_, _02393_, _22985_);
  nor _33964_ (_02395_, _02393_, _22985_);
  or _33965_ (_02396_, _02395_, _02394_);
  not _33966_ (_02397_, _00058_);
  and _33967_ (_02398_, _02391_, _02397_);
  nor _33968_ (_02399_, _02398_, _23904_);
  and _33969_ (_02400_, _02391_, _00014_);
  nor _33970_ (_02401_, _02400_, _23658_);
  nor _33971_ (_02402_, _02401_, _02399_);
  not _33972_ (_02403_, _23786_);
  not _33973_ (_02404_, _26817_);
  and _33974_ (_02405_, _02391_, _02404_);
  nor _33975_ (_02406_, _02405_, _02403_);
  and _33976_ (_02407_, _02405_, _02403_);
  nor _33977_ (_02408_, _02407_, _02406_);
  and _33978_ (_02409_, _02408_, _02402_);
  and _33979_ (_02410_, _02409_, _02396_);
  not _33980_ (_02411_, _02391_);
  and _33981_ (_02412_, _02411_, _26817_);
  and _33982_ (_02413_, _02391_, _00037_);
  nor _33983_ (_02414_, _02413_, _02412_);
  and _33984_ (_02415_, _02414_, _23039_);
  nor _33985_ (_02416_, _02414_, _23039_);
  or _33986_ (_02417_, _02416_, _02415_);
  not _33987_ (_02418_, _23067_);
  nor _33988_ (_02419_, _02388_, _00168_);
  nor _33989_ (_02420_, _02391_, _00014_);
  nor _33990_ (_02421_, _02420_, _02419_);
  nor _33991_ (_02422_, _02421_, _02418_);
  and _33992_ (_02423_, _02421_, _02418_);
  nor _33993_ (_02424_, _02423_, _02422_);
  not _33994_ (_02425_, _02424_);
  nor _33995_ (_02426_, _02425_, _02417_);
  or _33996_ (_02427_, _02388_, _00134_);
  or _33997_ (_02428_, _02391_, _00037_);
  nand _33998_ (_02429_, _02428_, _02427_);
  and _33999_ (_02430_, _02429_, _23020_);
  nor _34000_ (_02431_, _02429_, _23020_);
  nor _34001_ (_02432_, _02431_, _02430_);
  and _34002_ (_02433_, _02400_, _23658_);
  not _34003_ (_02434_, _02433_);
  and _34004_ (_02435_, _02398_, _23904_);
  not _34005_ (_02436_, _02435_);
  nor _34006_ (_02438_, _26781_, _22947_);
  and _34007_ (_02439_, _02438_, _02436_);
  and _34008_ (_02440_, _02439_, _02434_);
  and _34009_ (_02441_, _02440_, _02432_);
  and _34010_ (_02442_, _02441_, _02426_);
  and _34011_ (_02443_, _02442_, _02410_);
  not _34012_ (_02444_, _26777_);
  not _34013_ (_02445_, _02393_);
  and _34014_ (_02447_, _02428_, _02427_);
  and _34015_ (_02448_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and _34016_ (_02449_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or _34017_ (_02450_, _02449_, _02448_);
  and _34018_ (_02451_, _02450_, _02445_);
  and _34019_ (_02452_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and _34020_ (_02453_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or _34021_ (_02454_, _02453_, _02452_);
  and _34022_ (_02455_, _02454_, _02393_);
  or _34023_ (_02456_, _02455_, _02451_);
  or _34024_ (_02457_, _02456_, _02421_);
  not _34025_ (_02458_, _02414_);
  not _34026_ (_02459_, _02421_);
  and _34027_ (_02460_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and _34028_ (_02461_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or _34029_ (_02462_, _02461_, _02460_);
  and _34030_ (_02463_, _02462_, _02445_);
  and _34031_ (_02464_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and _34032_ (_02465_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or _34033_ (_02466_, _02465_, _02464_);
  and _34034_ (_02467_, _02466_, _02393_);
  or _34035_ (_02468_, _02467_, _02463_);
  or _34036_ (_02469_, _02468_, _02459_);
  and _34037_ (_02470_, _02469_, _02458_);
  and _34038_ (_02471_, _02470_, _02457_);
  or _34039_ (_02472_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or _34040_ (_02473_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and _34041_ (_02474_, _02473_, _02393_);
  and _34042_ (_02475_, _02474_, _02472_);
  or _34043_ (_02476_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or _34044_ (_02477_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and _34045_ (_02478_, _02477_, _02445_);
  and _34046_ (_02479_, _02478_, _02476_);
  or _34047_ (_02480_, _02479_, _02475_);
  or _34048_ (_02481_, _02480_, _02459_);
  or _34049_ (_02482_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or _34050_ (_02483_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and _34051_ (_02484_, _02483_, _02393_);
  and _34052_ (_02485_, _02484_, _02482_);
  or _34053_ (_02486_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or _34054_ (_02487_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and _34055_ (_02488_, _02487_, _02445_);
  and _34056_ (_02489_, _02488_, _02486_);
  or _34057_ (_02490_, _02489_, _02485_);
  or _34058_ (_02491_, _02490_, _02421_);
  and _34059_ (_02492_, _02491_, _02414_);
  and _34060_ (_02493_, _02492_, _02481_);
  or _34061_ (_02494_, _02493_, _02471_);
  or _34062_ (_02495_, _02494_, _02398_);
  not _34063_ (_02496_, _02398_);
  and _34064_ (_02497_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and _34065_ (_02498_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or _34066_ (_02499_, _02498_, _02393_);
  or _34067_ (_02500_, _02499_, _02497_);
  and _34068_ (_02501_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  and _34069_ (_02502_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or _34070_ (_02503_, _02502_, _02445_);
  or _34071_ (_02504_, _02503_, _02501_);
  and _34072_ (_02505_, _02504_, _02500_);
  or _34073_ (_02506_, _02505_, _02459_);
  and _34074_ (_02507_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and _34075_ (_02508_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or _34076_ (_02509_, _02508_, _02393_);
  or _34077_ (_02510_, _02509_, _02507_);
  and _34078_ (_02511_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and _34079_ (_02512_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or _34080_ (_02513_, _02512_, _02445_);
  or _34081_ (_02514_, _02513_, _02511_);
  and _34082_ (_02515_, _02514_, _02510_);
  or _34083_ (_02516_, _02515_, _02421_);
  and _34084_ (_02517_, _02516_, _02458_);
  and _34085_ (_02518_, _02517_, _02506_);
  or _34086_ (_02519_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or _34087_ (_02520_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  and _34088_ (_02521_, _02520_, _02519_);
  or _34089_ (_02522_, _02521_, _02445_);
  or _34090_ (_02523_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or _34091_ (_02524_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and _34092_ (_02525_, _02524_, _02523_);
  or _34093_ (_02526_, _02525_, _02393_);
  and _34094_ (_02527_, _02526_, _02522_);
  or _34095_ (_02528_, _02527_, _02459_);
  or _34096_ (_02529_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or _34097_ (_02530_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and _34098_ (_02531_, _02530_, _02529_);
  or _34099_ (_02532_, _02531_, _02445_);
  or _34100_ (_02533_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or _34101_ (_02534_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and _34102_ (_02535_, _02534_, _02533_);
  or _34103_ (_02536_, _02535_, _02393_);
  and _34104_ (_02537_, _02536_, _02532_);
  or _34105_ (_02538_, _02537_, _02421_);
  and _34106_ (_02540_, _02538_, _02414_);
  and _34107_ (_02541_, _02540_, _02528_);
  or _34108_ (_02542_, _02541_, _02518_);
  or _34109_ (_02543_, _02542_, _02496_);
  and _34110_ (_02544_, _02543_, _02400_);
  and _34111_ (_02545_, _02544_, _02495_);
  not _34112_ (_02546_, _02400_);
  and _34113_ (_02547_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and _34114_ (_02548_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or _34115_ (_02549_, _02548_, _02547_);
  and _34116_ (_02550_, _02549_, _02393_);
  and _34117_ (_02551_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and _34118_ (_02552_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or _34119_ (_02553_, _02552_, _02551_);
  and _34120_ (_02554_, _02553_, _02445_);
  or _34121_ (_02556_, _02554_, _02550_);
  or _34122_ (_02557_, _02556_, _02459_);
  and _34123_ (_02558_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  and _34124_ (_02559_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or _34125_ (_02560_, _02559_, _02558_);
  and _34126_ (_02561_, _02560_, _02393_);
  and _34127_ (_02562_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and _34128_ (_02563_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or _34129_ (_02564_, _02563_, _02562_);
  and _34130_ (_02565_, _02564_, _02445_);
  or _34131_ (_02566_, _02565_, _02561_);
  or _34132_ (_02567_, _02566_, _02421_);
  and _34133_ (_02568_, _02567_, _02458_);
  and _34134_ (_02569_, _02568_, _02557_);
  or _34135_ (_02570_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or _34136_ (_02572_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  and _34137_ (_02573_, _02572_, _02445_);
  and _34138_ (_02574_, _02573_, _02570_);
  or _34139_ (_02575_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or _34140_ (_02576_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and _34141_ (_02577_, _02576_, _02393_);
  and _34142_ (_02578_, _02577_, _02575_);
  or _34143_ (_02579_, _02578_, _02574_);
  or _34144_ (_02580_, _02579_, _02459_);
  or _34145_ (_02581_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or _34146_ (_02583_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  and _34147_ (_02584_, _02583_, _02445_);
  and _34148_ (_02585_, _02584_, _02581_);
  or _34149_ (_02586_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or _34150_ (_02587_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and _34151_ (_02588_, _02587_, _02393_);
  and _34152_ (_02589_, _02588_, _02586_);
  or _34153_ (_02590_, _02589_, _02585_);
  or _34154_ (_02591_, _02590_, _02421_);
  and _34155_ (_02592_, _02591_, _02414_);
  and _34156_ (_02593_, _02592_, _02580_);
  or _34157_ (_02594_, _02593_, _02569_);
  and _34158_ (_02595_, _02594_, _02496_);
  and _34159_ (_02596_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and _34160_ (_02597_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or _34161_ (_02598_, _02597_, _02596_);
  and _34162_ (_02599_, _02598_, _02393_);
  and _34163_ (_02600_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and _34164_ (_02601_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or _34165_ (_02602_, _02601_, _02600_);
  and _34166_ (_02603_, _02602_, _02445_);
  or _34167_ (_02604_, _02603_, _02599_);
  or _34168_ (_02605_, _02604_, _02459_);
  and _34169_ (_02606_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and _34170_ (_02607_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or _34171_ (_02608_, _02607_, _02606_);
  and _34172_ (_02609_, _02608_, _02393_);
  and _34173_ (_02610_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  and _34174_ (_02611_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or _34175_ (_02612_, _02611_, _02610_);
  and _34176_ (_02613_, _02612_, _02445_);
  or _34177_ (_02614_, _02613_, _02609_);
  or _34178_ (_02615_, _02614_, _02421_);
  and _34179_ (_02616_, _02615_, _02458_);
  and _34180_ (_02617_, _02616_, _02605_);
  or _34181_ (_02618_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or _34182_ (_02619_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and _34183_ (_02620_, _02619_, _02618_);
  and _34184_ (_02621_, _02620_, _02393_);
  or _34185_ (_02622_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or _34186_ (_02623_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and _34187_ (_02624_, _02623_, _02622_);
  and _34188_ (_02625_, _02624_, _02445_);
  or _34189_ (_02626_, _02625_, _02621_);
  or _34190_ (_02627_, _02626_, _02459_);
  or _34191_ (_02628_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or _34192_ (_02629_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  and _34193_ (_02630_, _02629_, _02628_);
  and _34194_ (_02631_, _02630_, _02393_);
  or _34195_ (_02632_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or _34196_ (_02633_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and _34197_ (_02634_, _02633_, _02632_);
  and _34198_ (_02635_, _02634_, _02445_);
  or _34199_ (_02636_, _02635_, _02631_);
  or _34200_ (_02637_, _02636_, _02421_);
  and _34201_ (_02638_, _02637_, _02414_);
  and _34202_ (_02639_, _02638_, _02627_);
  or _34203_ (_02640_, _02639_, _02617_);
  and _34204_ (_02641_, _02640_, _02398_);
  or _34205_ (_02642_, _02641_, _02595_);
  and _34206_ (_02643_, _02642_, _02546_);
  or _34207_ (_02644_, _02643_, _02545_);
  or _34208_ (_02645_, _02644_, _02405_);
  not _34209_ (_02646_, _02405_);
  and _34210_ (_02647_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  and _34211_ (_02648_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or _34212_ (_02649_, _02648_, _02647_);
  and _34213_ (_02650_, _02649_, _02393_);
  and _34214_ (_02651_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  and _34215_ (_02652_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or _34216_ (_02653_, _02652_, _02651_);
  and _34217_ (_02654_, _02653_, _02445_);
  or _34218_ (_02655_, _02654_, _02650_);
  and _34219_ (_02656_, _02655_, _02421_);
  and _34220_ (_02657_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  and _34221_ (_02658_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or _34222_ (_02659_, _02658_, _02657_);
  and _34223_ (_02660_, _02659_, _02393_);
  and _34224_ (_02661_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  and _34225_ (_02662_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or _34226_ (_02664_, _02662_, _02661_);
  and _34227_ (_02665_, _02664_, _02445_);
  or _34228_ (_02666_, _02665_, _02660_);
  and _34229_ (_02667_, _02666_, _02459_);
  or _34230_ (_02668_, _02667_, _02414_);
  or _34231_ (_02669_, _02668_, _02656_);
  or _34232_ (_02670_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or _34233_ (_02671_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  and _34234_ (_02672_, _02671_, _02670_);
  and _34235_ (_02673_, _02672_, _02393_);
  or _34236_ (_02674_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or _34237_ (_02675_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  and _34238_ (_02676_, _02675_, _02674_);
  and _34239_ (_02677_, _02676_, _02445_);
  or _34240_ (_02678_, _02677_, _02673_);
  and _34241_ (_02679_, _02678_, _02421_);
  or _34242_ (_02680_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or _34243_ (_02681_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  and _34244_ (_02682_, _02681_, _02680_);
  and _34245_ (_02683_, _02682_, _02393_);
  or _34246_ (_02684_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or _34247_ (_02685_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  and _34248_ (_02686_, _02685_, _02684_);
  and _34249_ (_02687_, _02686_, _02445_);
  or _34250_ (_02688_, _02687_, _02683_);
  and _34251_ (_02689_, _02688_, _02459_);
  or _34252_ (_02690_, _02689_, _02458_);
  or _34253_ (_02691_, _02690_, _02679_);
  and _34254_ (_02692_, _02691_, _02669_);
  or _34255_ (_02693_, _02692_, _02398_);
  and _34256_ (_02694_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and _34257_ (_02695_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or _34258_ (_02696_, _02695_, _02694_);
  and _34259_ (_02697_, _02696_, _02393_);
  and _34260_ (_02698_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  and _34261_ (_02699_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or _34262_ (_02700_, _02699_, _02698_);
  and _34263_ (_02701_, _02700_, _02445_);
  or _34264_ (_02702_, _02701_, _02697_);
  and _34265_ (_02703_, _02702_, _02421_);
  and _34266_ (_02704_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and _34267_ (_02705_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or _34268_ (_02706_, _02705_, _02704_);
  and _34269_ (_02707_, _02706_, _02393_);
  and _34270_ (_02708_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  and _34271_ (_02709_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or _34272_ (_02710_, _02709_, _02708_);
  and _34273_ (_02711_, _02710_, _02445_);
  or _34274_ (_02712_, _02711_, _02707_);
  and _34275_ (_02713_, _02712_, _02459_);
  or _34276_ (_02715_, _02713_, _02414_);
  or _34277_ (_02716_, _02715_, _02703_);
  or _34278_ (_02717_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or _34279_ (_02718_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and _34280_ (_02719_, _02718_, _02717_);
  and _34281_ (_02720_, _02719_, _02393_);
  or _34282_ (_02721_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or _34283_ (_02722_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  and _34284_ (_02723_, _02722_, _02721_);
  and _34285_ (_02724_, _02723_, _02445_);
  or _34286_ (_02725_, _02724_, _02720_);
  and _34287_ (_02726_, _02725_, _02421_);
  or _34288_ (_02727_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or _34289_ (_02728_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and _34290_ (_02729_, _02728_, _02727_);
  and _34291_ (_02730_, _02729_, _02393_);
  or _34292_ (_02731_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or _34293_ (_02732_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  and _34294_ (_02733_, _02732_, _02731_);
  and _34295_ (_02734_, _02733_, _02445_);
  or _34296_ (_02735_, _02734_, _02730_);
  and _34297_ (_02736_, _02735_, _02459_);
  or _34298_ (_02737_, _02736_, _02458_);
  or _34299_ (_02738_, _02737_, _02726_);
  and _34300_ (_02739_, _02738_, _02716_);
  or _34301_ (_02740_, _02739_, _02496_);
  and _34302_ (_02741_, _02740_, _02400_);
  and _34303_ (_02742_, _02741_, _02693_);
  and _34304_ (_02743_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and _34305_ (_02744_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or _34306_ (_02745_, _02744_, _02743_);
  and _34307_ (_02746_, _02745_, _02445_);
  and _34308_ (_02747_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  and _34309_ (_02748_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or _34310_ (_02749_, _02748_, _02747_);
  and _34311_ (_02750_, _02749_, _02393_);
  or _34312_ (_02751_, _02750_, _02746_);
  or _34313_ (_02752_, _02751_, _02459_);
  and _34314_ (_02753_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and _34315_ (_02754_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or _34316_ (_02755_, _02754_, _02753_);
  and _34317_ (_02756_, _02755_, _02445_);
  and _34318_ (_02757_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  and _34319_ (_02758_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or _34320_ (_02759_, _02758_, _02757_);
  and _34321_ (_02760_, _02759_, _02393_);
  or _34322_ (_02761_, _02760_, _02756_);
  or _34323_ (_02762_, _02761_, _02421_);
  and _34324_ (_02763_, _02762_, _02458_);
  and _34325_ (_02764_, _02763_, _02752_);
  or _34326_ (_02765_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or _34327_ (_02766_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and _34328_ (_02767_, _02766_, _02393_);
  and _34329_ (_02768_, _02767_, _02765_);
  or _34330_ (_02769_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or _34331_ (_02770_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and _34332_ (_02771_, _02770_, _02445_);
  and _34333_ (_02772_, _02771_, _02769_);
  or _34334_ (_02773_, _02772_, _02768_);
  or _34335_ (_02774_, _02773_, _02459_);
  or _34336_ (_02775_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or _34337_ (_02776_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  and _34338_ (_02777_, _02776_, _02393_);
  and _34339_ (_02778_, _02777_, _02775_);
  or _34340_ (_02779_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or _34341_ (_02780_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and _34342_ (_02781_, _02780_, _02445_);
  and _34343_ (_02782_, _02781_, _02779_);
  or _34344_ (_02783_, _02782_, _02778_);
  or _34345_ (_02784_, _02783_, _02421_);
  and _34346_ (_02785_, _02784_, _02414_);
  and _34347_ (_02786_, _02785_, _02774_);
  or _34348_ (_02787_, _02786_, _02764_);
  and _34349_ (_02788_, _02787_, _02496_);
  and _34350_ (_02789_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and _34351_ (_02790_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or _34352_ (_02791_, _02790_, _02393_);
  or _34353_ (_02792_, _02791_, _02789_);
  and _34354_ (_02793_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and _34355_ (_02794_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or _34356_ (_02795_, _02794_, _02445_);
  or _34357_ (_02796_, _02795_, _02793_);
  and _34358_ (_02797_, _02796_, _02792_);
  or _34359_ (_02798_, _02797_, _02459_);
  and _34360_ (_02799_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and _34361_ (_02800_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or _34362_ (_02801_, _02800_, _02393_);
  or _34363_ (_02802_, _02801_, _02799_);
  and _34364_ (_02803_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and _34365_ (_02804_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or _34366_ (_02805_, _02804_, _02445_);
  or _34367_ (_02806_, _02805_, _02803_);
  and _34368_ (_02807_, _02806_, _02802_);
  or _34369_ (_02808_, _02807_, _02421_);
  and _34370_ (_02809_, _02808_, _02458_);
  and _34371_ (_02810_, _02809_, _02798_);
  or _34372_ (_02811_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or _34373_ (_02812_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and _34374_ (_02813_, _02812_, _02811_);
  or _34375_ (_02814_, _02813_, _02445_);
  or _34376_ (_02815_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or _34377_ (_02816_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and _34378_ (_02817_, _02816_, _02815_);
  or _34379_ (_02818_, _02817_, _02393_);
  and _34380_ (_02819_, _02818_, _02814_);
  or _34381_ (_02820_, _02819_, _02459_);
  or _34382_ (_02821_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or _34383_ (_02822_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and _34384_ (_02823_, _02822_, _02821_);
  or _34385_ (_02824_, _02823_, _02445_);
  or _34386_ (_02825_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or _34387_ (_02827_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and _34388_ (_02828_, _02827_, _02825_);
  or _34389_ (_02829_, _02828_, _02393_);
  and _34390_ (_02830_, _02829_, _02824_);
  or _34391_ (_02831_, _02830_, _02421_);
  and _34392_ (_02832_, _02831_, _02414_);
  and _34393_ (_02833_, _02832_, _02820_);
  or _34394_ (_02834_, _02833_, _02810_);
  and _34395_ (_02835_, _02834_, _02398_);
  or _34396_ (_02836_, _02835_, _02788_);
  and _34397_ (_02837_, _02836_, _02546_);
  or _34398_ (_02838_, _02837_, _02742_);
  or _34399_ (_02839_, _02838_, _02646_);
  and _34400_ (_02840_, _02839_, _02645_);
  and _34401_ (_02841_, _02840_, _02444_);
  and _34402_ (_02842_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and _34403_ (_02843_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or _34404_ (_02845_, _02843_, _02842_);
  and _34405_ (_02846_, _02845_, _02393_);
  and _34406_ (_02847_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and _34407_ (_02848_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or _34408_ (_02849_, _02848_, _02847_);
  and _34409_ (_02850_, _02849_, _02445_);
  or _34410_ (_02851_, _02850_, _02846_);
  or _34411_ (_02852_, _02851_, _02459_);
  and _34412_ (_02853_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and _34413_ (_02854_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or _34414_ (_02855_, _02854_, _02853_);
  and _34415_ (_02856_, _02855_, _02393_);
  and _34416_ (_02857_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and _34417_ (_02858_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or _34418_ (_02859_, _02858_, _02857_);
  and _34419_ (_02860_, _02859_, _02445_);
  or _34420_ (_02861_, _02860_, _02856_);
  or _34421_ (_02862_, _02861_, _02421_);
  and _34422_ (_02863_, _02862_, _02458_);
  and _34423_ (_02864_, _02863_, _02852_);
  or _34424_ (_02865_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or _34425_ (_02866_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and _34426_ (_02868_, _02866_, _02865_);
  and _34427_ (_02869_, _02868_, _02393_);
  or _34428_ (_02870_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or _34429_ (_02871_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and _34430_ (_02872_, _02871_, _02870_);
  and _34431_ (_02873_, _02872_, _02445_);
  or _34432_ (_02875_, _02873_, _02869_);
  or _34433_ (_02877_, _02875_, _02459_);
  or _34434_ (_02878_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or _34435_ (_02879_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and _34436_ (_02881_, _02879_, _02878_);
  and _34437_ (_02883_, _02881_, _02393_);
  or _34438_ (_02884_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or _34439_ (_02885_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and _34440_ (_02886_, _02885_, _02884_);
  and _34441_ (_02887_, _02886_, _02445_);
  or _34442_ (_02888_, _02887_, _02883_);
  or _34443_ (_02889_, _02888_, _02421_);
  and _34444_ (_02890_, _02889_, _02414_);
  and _34445_ (_02891_, _02890_, _02877_);
  or _34446_ (_02892_, _02891_, _02864_);
  and _34447_ (_02894_, _02892_, _02398_);
  and _34448_ (_02895_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and _34449_ (_02896_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or _34450_ (_02897_, _02896_, _02895_);
  and _34451_ (_02898_, _02897_, _02393_);
  and _34452_ (_02899_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and _34453_ (_02900_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or _34454_ (_02901_, _02900_, _02899_);
  and _34455_ (_02902_, _02901_, _02445_);
  or _34456_ (_02904_, _02902_, _02898_);
  or _34457_ (_02905_, _02904_, _02459_);
  and _34458_ (_02907_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and _34459_ (_02909_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or _34460_ (_02910_, _02909_, _02907_);
  and _34461_ (_02912_, _02910_, _02393_);
  and _34462_ (_02913_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and _34463_ (_02914_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or _34464_ (_02915_, _02914_, _02913_);
  and _34465_ (_02916_, _02915_, _02445_);
  or _34466_ (_02917_, _02916_, _02912_);
  or _34467_ (_02918_, _02917_, _02421_);
  and _34468_ (_02919_, _02918_, _02458_);
  and _34469_ (_02920_, _02919_, _02905_);
  or _34470_ (_02921_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or _34471_ (_02922_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and _34472_ (_02924_, _02922_, _02445_);
  and _34473_ (_02925_, _02924_, _02921_);
  or _34474_ (_02926_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or _34475_ (_02927_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and _34476_ (_02928_, _02927_, _02393_);
  and _34477_ (_02929_, _02928_, _02926_);
  or _34478_ (_02930_, _02929_, _02925_);
  or _34479_ (_02931_, _02930_, _02459_);
  or _34480_ (_02932_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or _34481_ (_02933_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and _34482_ (_02934_, _02933_, _02445_);
  and _34483_ (_02935_, _02934_, _02932_);
  or _34484_ (_02936_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or _34485_ (_02937_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and _34486_ (_02938_, _02937_, _02393_);
  and _34487_ (_02939_, _02938_, _02936_);
  or _34488_ (_02940_, _02939_, _02935_);
  or _34489_ (_02941_, _02940_, _02421_);
  and _34490_ (_02942_, _02941_, _02414_);
  and _34491_ (_02943_, _02942_, _02931_);
  or _34492_ (_02944_, _02943_, _02920_);
  and _34493_ (_02945_, _02944_, _02496_);
  or _34494_ (_02946_, _02945_, _02894_);
  and _34495_ (_02947_, _02946_, _02546_);
  and _34496_ (_02948_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and _34497_ (_02949_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or _34498_ (_02950_, _02949_, _02948_);
  and _34499_ (_02951_, _02950_, _02393_);
  and _34500_ (_02952_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and _34501_ (_02953_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or _34502_ (_02954_, _02953_, _02952_);
  and _34503_ (_02955_, _02954_, _02445_);
  or _34504_ (_02956_, _02955_, _02951_);
  and _34505_ (_02957_, _02956_, _02421_);
  and _34506_ (_02958_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and _34507_ (_02959_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or _34508_ (_02960_, _02959_, _02958_);
  and _34509_ (_02961_, _02960_, _02393_);
  and _34510_ (_02962_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and _34511_ (_02963_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or _34512_ (_02964_, _02963_, _02962_);
  and _34513_ (_02965_, _02964_, _02445_);
  or _34514_ (_02966_, _02965_, _02961_);
  and _34515_ (_02967_, _02966_, _02459_);
  or _34516_ (_02968_, _02967_, _02957_);
  and _34517_ (_02969_, _02968_, _02458_);
  or _34518_ (_02970_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or _34519_ (_02971_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and _34520_ (_02973_, _02971_, _02445_);
  and _34521_ (_02974_, _02973_, _02970_);
  or _34522_ (_02975_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or _34523_ (_02976_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and _34524_ (_02977_, _02976_, _02393_);
  and _34525_ (_02978_, _02977_, _02975_);
  or _34526_ (_02979_, _02978_, _02974_);
  and _34527_ (_02980_, _02979_, _02421_);
  or _34528_ (_02981_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or _34529_ (_02982_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and _34530_ (_02983_, _02982_, _02445_);
  and _34531_ (_02984_, _02983_, _02981_);
  or _34532_ (_02985_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or _34533_ (_02986_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and _34534_ (_02987_, _02986_, _02393_);
  and _34535_ (_02988_, _02987_, _02985_);
  or _34536_ (_02989_, _02988_, _02984_);
  and _34537_ (_02990_, _02989_, _02459_);
  or _34538_ (_02991_, _02990_, _02980_);
  and _34539_ (_02992_, _02991_, _02414_);
  or _34540_ (_02993_, _02992_, _02969_);
  and _34541_ (_02994_, _02993_, _02496_);
  and _34542_ (_02995_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and _34543_ (_02997_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or _34544_ (_02998_, _02997_, _02995_);
  and _34545_ (_02999_, _02998_, _02393_);
  and _34546_ (_03000_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and _34547_ (_03001_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or _34548_ (_03002_, _03001_, _03000_);
  and _34549_ (_03003_, _03002_, _02445_);
  or _34550_ (_03004_, _03003_, _02999_);
  and _34551_ (_03005_, _03004_, _02421_);
  and _34552_ (_03006_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and _34553_ (_03007_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or _34554_ (_03008_, _03007_, _03006_);
  and _34555_ (_03009_, _03008_, _02393_);
  and _34556_ (_03010_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and _34557_ (_03011_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or _34558_ (_03012_, _03011_, _03010_);
  and _34559_ (_03013_, _03012_, _02445_);
  or _34560_ (_03014_, _03013_, _03009_);
  and _34561_ (_03015_, _03014_, _02459_);
  or _34562_ (_03016_, _03015_, _03005_);
  and _34563_ (_03017_, _03016_, _02458_);
  or _34564_ (_03018_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or _34565_ (_03019_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and _34566_ (_03020_, _03019_, _03018_);
  and _34567_ (_03021_, _03020_, _02393_);
  or _34568_ (_03022_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or _34569_ (_03023_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and _34570_ (_03024_, _03023_, _03022_);
  and _34571_ (_03025_, _03024_, _02445_);
  or _34572_ (_03026_, _03025_, _03021_);
  and _34573_ (_03027_, _03026_, _02421_);
  or _34574_ (_03028_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or _34575_ (_03029_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and _34576_ (_03030_, _03029_, _03028_);
  and _34577_ (_03031_, _03030_, _02393_);
  or _34578_ (_03032_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or _34579_ (_03033_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and _34580_ (_03034_, _03033_, _03032_);
  and _34581_ (_03035_, _03034_, _02445_);
  or _34582_ (_03036_, _03035_, _03031_);
  and _34583_ (_03037_, _03036_, _02459_);
  or _34584_ (_03038_, _03037_, _03027_);
  and _34585_ (_03039_, _03038_, _02414_);
  or _34586_ (_03040_, _03039_, _03017_);
  and _34587_ (_03041_, _03040_, _02398_);
  or _34588_ (_03042_, _03041_, _02994_);
  and _34589_ (_03043_, _03042_, _02400_);
  or _34590_ (_03044_, _03043_, _02947_);
  or _34591_ (_03045_, _03044_, _02405_);
  and _34592_ (_03047_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and _34593_ (_03048_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or _34594_ (_03049_, _03048_, _03047_);
  and _34595_ (_03050_, _03049_, _02393_);
  and _34596_ (_03051_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and _34597_ (_03053_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or _34598_ (_03054_, _03053_, _03051_);
  and _34599_ (_03055_, _03054_, _02445_);
  or _34600_ (_03056_, _03055_, _03050_);
  or _34601_ (_03057_, _03056_, _02459_);
  and _34602_ (_03058_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and _34603_ (_03059_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or _34604_ (_03060_, _03059_, _03058_);
  and _34605_ (_03061_, _03060_, _02393_);
  and _34606_ (_03062_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and _34607_ (_03063_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or _34608_ (_03064_, _03063_, _03062_);
  and _34609_ (_03065_, _03064_, _02445_);
  or _34610_ (_03066_, _03065_, _03061_);
  or _34611_ (_03067_, _03066_, _02421_);
  and _34612_ (_03068_, _03067_, _02458_);
  and _34613_ (_03070_, _03068_, _03057_);
  or _34614_ (_03071_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or _34615_ (_03072_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and _34616_ (_03073_, _03072_, _02445_);
  and _34617_ (_03074_, _03073_, _03071_);
  or _34618_ (_03075_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or _34619_ (_03076_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and _34620_ (_03077_, _03076_, _02393_);
  and _34621_ (_03078_, _03077_, _03075_);
  or _34622_ (_03079_, _03078_, _03074_);
  or _34623_ (_03080_, _03079_, _02459_);
  or _34624_ (_03081_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or _34625_ (_03082_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and _34626_ (_03084_, _03082_, _02445_);
  and _34627_ (_03085_, _03084_, _03081_);
  or _34628_ (_03086_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or _34629_ (_03087_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and _34630_ (_03088_, _03087_, _02393_);
  and _34631_ (_03089_, _03088_, _03086_);
  or _34632_ (_03090_, _03089_, _03085_);
  or _34633_ (_03091_, _03090_, _02421_);
  and _34634_ (_03092_, _03091_, _02414_);
  and _34635_ (_03093_, _03092_, _03080_);
  or _34636_ (_03094_, _03093_, _03070_);
  and _34637_ (_03095_, _03094_, _02496_);
  and _34638_ (_03096_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and _34639_ (_03097_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or _34640_ (_03098_, _03097_, _03096_);
  and _34641_ (_03099_, _03098_, _02393_);
  and _34642_ (_03100_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and _34643_ (_03101_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or _34644_ (_03102_, _03101_, _03100_);
  and _34645_ (_03103_, _03102_, _02445_);
  or _34646_ (_03104_, _03103_, _03099_);
  or _34647_ (_03105_, _03104_, _02459_);
  and _34648_ (_03106_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and _34649_ (_03107_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or _34650_ (_03109_, _03107_, _03106_);
  and _34651_ (_03110_, _03109_, _02393_);
  and _34652_ (_03111_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and _34653_ (_03112_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or _34654_ (_03113_, _03112_, _03111_);
  and _34655_ (_03115_, _03113_, _02445_);
  or _34656_ (_03116_, _03115_, _03110_);
  or _34657_ (_03118_, _03116_, _02421_);
  and _34658_ (_03119_, _03118_, _02458_);
  and _34659_ (_03120_, _03119_, _03105_);
  or _34660_ (_03121_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or _34661_ (_03122_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and _34662_ (_03124_, _03122_, _03121_);
  and _34663_ (_03126_, _03124_, _02393_);
  or _34664_ (_03127_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or _34665_ (_03128_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and _34666_ (_03130_, _03128_, _03127_);
  and _34667_ (_03131_, _03130_, _02445_);
  or _34668_ (_03132_, _03131_, _03126_);
  or _34669_ (_03133_, _03132_, _02459_);
  or _34670_ (_03134_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or _34671_ (_03135_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and _34672_ (_03136_, _03135_, _03134_);
  and _34673_ (_03137_, _03136_, _02393_);
  or _34674_ (_03138_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or _34675_ (_03140_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and _34676_ (_03141_, _03140_, _03138_);
  and _34677_ (_03142_, _03141_, _02445_);
  or _34678_ (_03143_, _03142_, _03137_);
  or _34679_ (_03145_, _03143_, _02421_);
  and _34680_ (_03146_, _03145_, _02414_);
  and _34681_ (_03147_, _03146_, _03133_);
  or _34682_ (_03148_, _03147_, _03120_);
  and _34683_ (_03149_, _03148_, _02398_);
  or _34684_ (_03150_, _03149_, _03095_);
  and _34685_ (_03151_, _03150_, _02546_);
  or _34686_ (_03152_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or _34687_ (_03153_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and _34688_ (_03154_, _03153_, _03152_);
  and _34689_ (_03155_, _03154_, _02393_);
  or _34690_ (_03156_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or _34691_ (_03157_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and _34692_ (_03158_, _03157_, _03156_);
  and _34693_ (_03159_, _03158_, _02445_);
  or _34694_ (_03161_, _03159_, _03155_);
  and _34695_ (_03162_, _03161_, _02459_);
  or _34696_ (_03163_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or _34697_ (_03165_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and _34698_ (_03166_, _03165_, _03163_);
  and _34699_ (_03167_, _03166_, _02393_);
  or _34700_ (_03169_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or _34701_ (_03170_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and _34702_ (_03171_, _03170_, _03169_);
  and _34703_ (_03172_, _03171_, _02445_);
  or _34704_ (_03173_, _03172_, _03167_);
  and _34705_ (_03174_, _03173_, _02421_);
  or _34706_ (_03176_, _03174_, _03162_);
  and _34707_ (_03178_, _03176_, _02414_);
  and _34708_ (_03179_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and _34709_ (_03180_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or _34710_ (_03181_, _03180_, _03179_);
  and _34711_ (_03182_, _03181_, _02393_);
  and _34712_ (_03183_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and _34713_ (_03184_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or _34714_ (_03185_, _03184_, _03183_);
  and _34715_ (_03186_, _03185_, _02445_);
  or _34716_ (_03187_, _03186_, _03182_);
  and _34717_ (_03188_, _03187_, _02459_);
  and _34718_ (_03189_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and _34719_ (_03190_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or _34720_ (_03191_, _03190_, _03189_);
  and _34721_ (_03192_, _03191_, _02393_);
  and _34722_ (_03193_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and _34723_ (_03195_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or _34724_ (_03196_, _03195_, _03193_);
  and _34725_ (_03197_, _03196_, _02445_);
  or _34726_ (_03198_, _03197_, _03192_);
  and _34727_ (_03200_, _03198_, _02421_);
  or _34728_ (_03201_, _03200_, _03188_);
  and _34729_ (_03202_, _03201_, _02458_);
  or _34730_ (_03203_, _03202_, _03178_);
  and _34731_ (_03204_, _03203_, _02398_);
  or _34732_ (_03205_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or _34733_ (_03206_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and _34734_ (_03207_, _03206_, _02445_);
  and _34735_ (_03208_, _03207_, _03205_);
  or _34736_ (_03210_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or _34737_ (_03212_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and _34738_ (_03213_, _03212_, _02393_);
  and _34739_ (_03214_, _03213_, _03210_);
  or _34740_ (_03215_, _03214_, _03208_);
  and _34741_ (_03216_, _03215_, _02459_);
  or _34742_ (_03217_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or _34743_ (_03218_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and _34744_ (_03219_, _03218_, _02445_);
  and _34745_ (_03220_, _03219_, _03217_);
  or _34746_ (_03221_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or _34747_ (_03223_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and _34748_ (_03224_, _03223_, _02393_);
  and _34749_ (_03226_, _03224_, _03221_);
  or _34750_ (_03228_, _03226_, _03220_);
  and _34751_ (_03229_, _03228_, _02421_);
  or _34752_ (_03230_, _03229_, _03216_);
  and _34753_ (_03232_, _03230_, _02414_);
  and _34754_ (_03234_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and _34755_ (_03235_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or _34756_ (_03236_, _03235_, _03234_);
  and _34757_ (_03237_, _03236_, _02393_);
  and _34758_ (_03238_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and _34759_ (_03239_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or _34760_ (_03240_, _03239_, _03238_);
  and _34761_ (_03241_, _03240_, _02445_);
  or _34762_ (_03242_, _03241_, _03237_);
  and _34763_ (_03243_, _03242_, _02459_);
  and _34764_ (_03245_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and _34765_ (_03246_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or _34766_ (_03247_, _03246_, _03245_);
  and _34767_ (_03248_, _03247_, _02393_);
  and _34768_ (_03249_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and _34769_ (_03250_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or _34770_ (_03251_, _03250_, _03249_);
  and _34771_ (_03252_, _03251_, _02445_);
  or _34772_ (_03253_, _03252_, _03248_);
  and _34773_ (_03254_, _03253_, _02421_);
  or _34774_ (_03255_, _03254_, _03243_);
  and _34775_ (_03256_, _03255_, _02458_);
  or _34776_ (_03257_, _03256_, _03232_);
  and _34777_ (_03258_, _03257_, _02496_);
  or _34778_ (_03259_, _03258_, _03204_);
  and _34779_ (_03260_, _03259_, _02400_);
  or _34780_ (_03261_, _03260_, _03151_);
  or _34781_ (_03262_, _03261_, _02646_);
  and _34782_ (_03263_, _03262_, _03045_);
  and _34783_ (_03264_, _03263_, _26777_);
  or _34784_ (_03265_, _03264_, _02841_);
  or _34785_ (_03266_, _03265_, _02443_);
  not _34786_ (_03267_, _02443_);
  or _34787_ (_03268_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and _34788_ (_03269_, _03268_, _22762_);
  and _34789_ (_22712_, _03269_, _03266_);
  and _34790_ (_03271_, _02374_, _23649_);
  and _34791_ (_03272_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  or _34792_ (_22713_, _03272_, _03271_);
  or _34793_ (_03273_, _02268_, _24537_);
  and _34794_ (_03274_, _26625_, _24584_);
  and _34795_ (_03275_, _25621_, _26582_);
  or _34796_ (_03276_, _03275_, _24585_);
  or _34797_ (_03277_, _03276_, _03274_);
  or _34798_ (_03278_, _03277_, _03273_);
  and _34799_ (_03279_, _03278_, _22768_);
  and _34800_ (_03280_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  or _34801_ (_03281_, _03280_, _25664_);
  or _34802_ (_03283_, _03281_, _03279_);
  and _34803_ (_26866_[1], _03283_, _22762_);
  and _34804_ (_03284_, _25656_, _23898_);
  and _34805_ (_03285_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or _34806_ (_22714_, _03285_, _03284_);
  and _34807_ (_03286_, _25142_, _23946_);
  and _34808_ (_03288_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or _34809_ (_22715_, _03288_, _03286_);
  and _34810_ (_03290_, _02350_, _23747_);
  and _34811_ (_03292_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or _34812_ (_26978_, _03292_, _03290_);
  and _34813_ (_03293_, _25649_, _23747_);
  and _34814_ (_03295_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or _34815_ (_22716_, _03295_, _03293_);
  and _34816_ (_03296_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  and _34817_ (_03297_, _02245_, _23747_);
  or _34818_ (_22717_, _03297_, _03296_);
  and _34819_ (_03298_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  and _34820_ (_03299_, _02245_, _23824_);
  or _34821_ (_22718_, _03299_, _03298_);
  and _34822_ (_03300_, _23752_, _23664_);
  and _34823_ (_03301_, _03300_, _23747_);
  not _34824_ (_03302_, _03300_);
  and _34825_ (_03303_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or _34826_ (_22719_, _03303_, _03301_);
  and _34827_ (_03305_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _22762_);
  and _34828_ (_03306_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _22762_);
  and _34829_ (_03307_, _03306_, _01772_);
  or _34830_ (_26895_[7], _03307_, _03305_);
  or _34831_ (_03308_, _26622_, _26646_);
  and _34832_ (_03309_, _26645_, _24613_);
  and _34833_ (_03311_, _24597_, _24538_);
  and _34834_ (_03312_, _03311_, _25667_);
  or _34835_ (_03313_, _03312_, _03309_);
  or _34836_ (_03314_, _03313_, _03308_);
  or _34837_ (_03315_, _26669_, _26657_);
  or _34838_ (_03316_, _26581_, _26615_);
  or _34839_ (_03317_, _26636_, _26665_);
  or _34840_ (_03318_, _03317_, _03316_);
  or _34841_ (_03319_, _03318_, _03315_);
  or _34842_ (_03320_, _03319_, _03314_);
  and _34843_ (_03321_, _26568_, _24538_);
  and _34844_ (_03322_, _24552_, _24445_);
  or _34845_ (_03323_, _03322_, _03321_);
  or _34846_ (_03324_, _26661_, _24608_);
  or _34847_ (_03325_, _03324_, _03323_);
  or _34848_ (_03327_, _03325_, _03320_);
  and _34849_ (_03328_, _03327_, _22768_);
  and _34850_ (_03329_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _34851_ (_03330_, _03321_, _03309_);
  and _34852_ (_03331_, _03330_, _24566_);
  or _34853_ (_03332_, _03331_, _25664_);
  and _34854_ (_03334_, _26645_, _24567_);
  and _34855_ (_03335_, _03334_, _24566_);
  or _34856_ (_03336_, _03335_, _03332_);
  or _34857_ (_03337_, _03336_, _03329_);
  or _34858_ (_03338_, _03337_, _03328_);
  and _34859_ (_26868_[0], _03338_, _22762_);
  and _34860_ (_03339_, _01809_, _24282_);
  and _34861_ (_03340_, _03339_, _23649_);
  not _34862_ (_03342_, _03339_);
  and _34863_ (_03343_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or _34864_ (_22720_, _03343_, _03340_);
  and _34865_ (_03344_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and _34866_ (_03345_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or _34867_ (_03347_, _03345_, _03344_);
  and _34868_ (_03348_, _03347_, _02393_);
  and _34869_ (_03349_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and _34870_ (_03350_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or _34871_ (_03351_, _03350_, _03349_);
  and _34872_ (_03352_, _03351_, _02445_);
  or _34873_ (_03353_, _03352_, _03348_);
  and _34874_ (_03354_, _03353_, _02421_);
  and _34875_ (_03355_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and _34876_ (_03356_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or _34877_ (_03358_, _03356_, _03355_);
  and _34878_ (_03359_, _03358_, _02393_);
  and _34879_ (_03360_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and _34880_ (_03361_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or _34881_ (_03363_, _03361_, _03360_);
  and _34882_ (_03364_, _03363_, _02445_);
  or _34883_ (_03366_, _03364_, _03359_);
  and _34884_ (_03367_, _03366_, _02459_);
  or _34885_ (_03368_, _03367_, _03354_);
  and _34886_ (_03369_, _03368_, _02458_);
  or _34887_ (_03370_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or _34888_ (_03372_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and _34889_ (_03373_, _03372_, _03370_);
  and _34890_ (_03374_, _03373_, _02393_);
  or _34891_ (_03375_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or _34892_ (_03376_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and _34893_ (_03377_, _03376_, _03375_);
  and _34894_ (_03378_, _03377_, _02445_);
  or _34895_ (_03379_, _03378_, _03374_);
  and _34896_ (_03380_, _03379_, _02421_);
  or _34897_ (_03381_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or _34898_ (_03382_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and _34899_ (_03383_, _03382_, _03381_);
  and _34900_ (_03384_, _03383_, _02393_);
  or _34901_ (_03385_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or _34902_ (_03386_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and _34903_ (_03387_, _03386_, _03385_);
  and _34904_ (_03388_, _03387_, _02445_);
  or _34905_ (_03389_, _03388_, _03384_);
  and _34906_ (_03390_, _03389_, _02459_);
  or _34907_ (_03392_, _03390_, _03380_);
  and _34908_ (_03393_, _03392_, _02414_);
  or _34909_ (_03394_, _03393_, _03369_);
  and _34910_ (_03395_, _03394_, _02398_);
  and _34911_ (_03396_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and _34912_ (_03397_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or _34913_ (_03399_, _03397_, _03396_);
  and _34914_ (_03401_, _03399_, _02393_);
  and _34915_ (_03402_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and _34916_ (_03403_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or _34917_ (_03404_, _03403_, _03402_);
  and _34918_ (_03405_, _03404_, _02445_);
  or _34919_ (_03407_, _03405_, _03401_);
  and _34920_ (_03408_, _03407_, _02421_);
  and _34921_ (_03410_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and _34922_ (_03411_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or _34923_ (_03412_, _03411_, _03410_);
  and _34924_ (_03413_, _03412_, _02393_);
  and _34925_ (_03414_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and _34926_ (_03415_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or _34927_ (_03416_, _03415_, _03414_);
  and _34928_ (_03417_, _03416_, _02445_);
  or _34929_ (_03419_, _03417_, _03413_);
  and _34930_ (_03420_, _03419_, _02459_);
  or _34931_ (_03421_, _03420_, _03408_);
  and _34932_ (_03422_, _03421_, _02458_);
  or _34933_ (_03423_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or _34934_ (_03424_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and _34935_ (_03425_, _03424_, _02445_);
  and _34936_ (_03426_, _03425_, _03423_);
  or _34937_ (_03427_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or _34938_ (_03428_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and _34939_ (_03429_, _03428_, _02393_);
  and _34940_ (_03430_, _03429_, _03427_);
  or _34941_ (_03431_, _03430_, _03426_);
  and _34942_ (_03432_, _03431_, _02421_);
  or _34943_ (_03434_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or _34944_ (_03435_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and _34945_ (_03437_, _03435_, _02445_);
  and _34946_ (_03438_, _03437_, _03434_);
  or _34947_ (_03440_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or _34948_ (_03442_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and _34949_ (_03443_, _03442_, _02393_);
  and _34950_ (_03445_, _03443_, _03440_);
  or _34951_ (_03446_, _03445_, _03438_);
  and _34952_ (_03447_, _03446_, _02459_);
  or _34953_ (_03449_, _03447_, _03432_);
  and _34954_ (_03450_, _03449_, _02414_);
  or _34955_ (_03451_, _03450_, _03422_);
  and _34956_ (_03452_, _03451_, _02496_);
  or _34957_ (_03454_, _03452_, _03395_);
  and _34958_ (_03455_, _03454_, _02400_);
  and _34959_ (_03456_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and _34960_ (_03457_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or _34961_ (_03458_, _03457_, _03456_);
  and _34962_ (_03459_, _03458_, _02393_);
  and _34963_ (_03460_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and _34964_ (_03461_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or _34965_ (_03462_, _03461_, _03460_);
  and _34966_ (_03464_, _03462_, _02445_);
  or _34967_ (_03465_, _03464_, _03459_);
  or _34968_ (_03466_, _03465_, _02459_);
  and _34969_ (_03467_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and _34970_ (_03468_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or _34971_ (_03469_, _03468_, _03467_);
  and _34972_ (_03470_, _03469_, _02393_);
  and _34973_ (_03471_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and _34974_ (_03472_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or _34975_ (_03473_, _03472_, _03471_);
  and _34976_ (_03474_, _03473_, _02445_);
  or _34977_ (_03475_, _03474_, _03470_);
  or _34978_ (_03476_, _03475_, _02421_);
  and _34979_ (_03478_, _03476_, _02458_);
  and _34980_ (_03479_, _03478_, _03466_);
  or _34981_ (_03480_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or _34982_ (_03481_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and _34983_ (_03482_, _03481_, _02445_);
  and _34984_ (_03483_, _03482_, _03480_);
  or _34985_ (_03484_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or _34986_ (_03485_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and _34987_ (_03487_, _03485_, _02393_);
  and _34988_ (_03488_, _03487_, _03484_);
  or _34989_ (_03489_, _03488_, _03483_);
  or _34990_ (_03490_, _03489_, _02459_);
  or _34991_ (_03491_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or _34992_ (_03492_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and _34993_ (_03493_, _03492_, _02445_);
  and _34994_ (_03494_, _03493_, _03491_);
  or _34995_ (_03495_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or _34996_ (_03496_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and _34997_ (_03497_, _03496_, _02393_);
  and _34998_ (_03498_, _03497_, _03495_);
  or _34999_ (_03499_, _03498_, _03494_);
  or _35000_ (_03501_, _03499_, _02421_);
  and _35001_ (_03502_, _03501_, _02414_);
  and _35002_ (_03503_, _03502_, _03490_);
  or _35003_ (_03504_, _03503_, _03479_);
  and _35004_ (_03506_, _03504_, _02496_);
  and _35005_ (_03507_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and _35006_ (_03508_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or _35007_ (_03510_, _03508_, _03507_);
  and _35008_ (_03511_, _03510_, _02393_);
  and _35009_ (_03512_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and _35010_ (_03513_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or _35011_ (_03514_, _03513_, _03512_);
  and _35012_ (_03515_, _03514_, _02445_);
  or _35013_ (_03516_, _03515_, _03511_);
  or _35014_ (_03517_, _03516_, _02459_);
  and _35015_ (_03519_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and _35016_ (_03520_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or _35017_ (_03521_, _03520_, _03519_);
  and _35018_ (_03522_, _03521_, _02393_);
  and _35019_ (_03523_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and _35020_ (_03525_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or _35021_ (_03526_, _03525_, _03523_);
  and _35022_ (_03527_, _03526_, _02445_);
  or _35023_ (_03528_, _03527_, _03522_);
  or _35024_ (_03529_, _03528_, _02421_);
  and _35025_ (_03530_, _03529_, _02458_);
  and _35026_ (_03531_, _03530_, _03517_);
  or _35027_ (_03532_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or _35028_ (_03533_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and _35029_ (_03534_, _03533_, _03532_);
  and _35030_ (_03535_, _03534_, _02393_);
  or _35031_ (_03536_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or _35032_ (_03537_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and _35033_ (_03538_, _03537_, _03536_);
  and _35034_ (_03540_, _03538_, _02445_);
  or _35035_ (_03541_, _03540_, _03535_);
  or _35036_ (_03543_, _03541_, _02459_);
  or _35037_ (_03544_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or _35038_ (_03545_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and _35039_ (_03546_, _03545_, _03544_);
  and _35040_ (_03547_, _03546_, _02393_);
  or _35041_ (_03548_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or _35042_ (_03549_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and _35043_ (_03550_, _03549_, _03548_);
  and _35044_ (_03551_, _03550_, _02445_);
  or _35045_ (_03552_, _03551_, _03547_);
  or _35046_ (_03553_, _03552_, _02421_);
  and _35047_ (_03554_, _03553_, _02414_);
  and _35048_ (_03555_, _03554_, _03543_);
  or _35049_ (_03556_, _03555_, _03531_);
  and _35050_ (_03558_, _03556_, _02398_);
  or _35051_ (_03559_, _03558_, _03506_);
  and _35052_ (_03560_, _03559_, _02546_);
  or _35053_ (_03561_, _03560_, _03455_);
  and _35054_ (_03562_, _03561_, _02646_);
  or _35055_ (_03563_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or _35056_ (_03564_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and _35057_ (_03565_, _03564_, _02445_);
  and _35058_ (_03566_, _03565_, _03563_);
  or _35059_ (_03567_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or _35060_ (_03568_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and _35061_ (_03569_, _03568_, _02393_);
  and _35062_ (_03570_, _03569_, _03567_);
  or _35063_ (_03571_, _03570_, _03566_);
  and _35064_ (_03572_, _03571_, _02459_);
  or _35065_ (_03573_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or _35066_ (_03575_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and _35067_ (_03576_, _03575_, _02445_);
  and _35068_ (_03578_, _03576_, _03573_);
  or _35069_ (_03579_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or _35070_ (_03580_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and _35071_ (_03581_, _03580_, _02393_);
  and _35072_ (_03582_, _03581_, _03579_);
  or _35073_ (_03583_, _03582_, _03578_);
  and _35074_ (_03584_, _03583_, _02421_);
  or _35075_ (_03585_, _03584_, _03572_);
  and _35076_ (_03586_, _03585_, _02414_);
  and _35077_ (_03587_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and _35078_ (_03588_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or _35079_ (_03589_, _03588_, _03587_);
  and _35080_ (_03590_, _03589_, _02393_);
  and _35081_ (_03591_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and _35082_ (_03592_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or _35083_ (_03593_, _03592_, _03591_);
  and _35084_ (_03594_, _03593_, _02445_);
  or _35085_ (_03595_, _03594_, _03590_);
  and _35086_ (_03596_, _03595_, _02459_);
  and _35087_ (_03597_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and _35088_ (_03598_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or _35089_ (_03599_, _03598_, _03597_);
  and _35090_ (_03600_, _03599_, _02393_);
  and _35091_ (_03601_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and _35092_ (_03602_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or _35093_ (_03603_, _03602_, _03601_);
  and _35094_ (_03604_, _03603_, _02445_);
  or _35095_ (_03606_, _03604_, _03600_);
  and _35096_ (_03607_, _03606_, _02421_);
  or _35097_ (_03609_, _03607_, _03596_);
  and _35098_ (_03610_, _03609_, _02458_);
  or _35099_ (_03611_, _03610_, _03586_);
  and _35100_ (_03612_, _03611_, _02496_);
  or _35101_ (_03614_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or _35102_ (_03615_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and _35103_ (_03616_, _03615_, _03614_);
  and _35104_ (_03617_, _03616_, _02393_);
  or _35105_ (_03618_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or _35106_ (_03619_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and _35107_ (_03620_, _03619_, _03618_);
  and _35108_ (_03621_, _03620_, _02445_);
  or _35109_ (_03622_, _03621_, _03617_);
  and _35110_ (_03623_, _03622_, _02459_);
  or _35111_ (_03624_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or _35112_ (_03625_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and _35113_ (_03626_, _03625_, _03624_);
  and _35114_ (_03627_, _03626_, _02393_);
  or _35115_ (_03629_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or _35116_ (_03630_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and _35117_ (_03631_, _03630_, _03629_);
  and _35118_ (_03632_, _03631_, _02445_);
  or _35119_ (_03633_, _03632_, _03627_);
  and _35120_ (_03634_, _03633_, _02421_);
  or _35121_ (_03635_, _03634_, _03623_);
  and _35122_ (_03636_, _03635_, _02414_);
  and _35123_ (_03637_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and _35124_ (_03639_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or _35125_ (_03640_, _03639_, _03637_);
  and _35126_ (_03641_, _03640_, _02393_);
  and _35127_ (_03642_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and _35128_ (_03643_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or _35129_ (_03644_, _03643_, _03642_);
  and _35130_ (_03645_, _03644_, _02445_);
  or _35131_ (_03646_, _03645_, _03641_);
  and _35132_ (_03647_, _03646_, _02459_);
  and _35133_ (_03648_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and _35134_ (_03649_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or _35135_ (_03650_, _03649_, _03648_);
  and _35136_ (_03651_, _03650_, _02393_);
  and _35137_ (_03652_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and _35138_ (_03653_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or _35139_ (_03654_, _03653_, _03652_);
  and _35140_ (_03655_, _03654_, _02445_);
  or _35141_ (_03657_, _03655_, _03651_);
  and _35142_ (_03658_, _03657_, _02421_);
  or _35143_ (_03659_, _03658_, _03647_);
  and _35144_ (_03660_, _03659_, _02458_);
  or _35145_ (_03661_, _03660_, _03636_);
  and _35146_ (_03662_, _03661_, _02398_);
  or _35147_ (_03663_, _03662_, _03612_);
  and _35148_ (_03665_, _03663_, _02400_);
  and _35149_ (_03666_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and _35150_ (_03667_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or _35151_ (_03668_, _03667_, _03666_);
  and _35152_ (_03669_, _03668_, _02393_);
  and _35153_ (_03670_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and _35154_ (_03671_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or _35155_ (_03672_, _03671_, _03670_);
  and _35156_ (_03673_, _03672_, _02445_);
  or _35157_ (_03674_, _03673_, _03669_);
  or _35158_ (_03675_, _03674_, _02459_);
  and _35159_ (_03677_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and _35160_ (_03678_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or _35161_ (_03679_, _03678_, _03677_);
  and _35162_ (_03681_, _03679_, _02393_);
  and _35163_ (_03682_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and _35164_ (_03684_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or _35165_ (_03685_, _03684_, _03682_);
  and _35166_ (_03686_, _03685_, _02445_);
  or _35167_ (_03687_, _03686_, _03681_);
  or _35168_ (_03688_, _03687_, _02421_);
  and _35169_ (_03689_, _03688_, _02458_);
  and _35170_ (_03690_, _03689_, _03675_);
  or _35171_ (_03691_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or _35172_ (_03692_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and _35173_ (_03693_, _03692_, _03691_);
  and _35174_ (_03694_, _03693_, _02393_);
  or _35175_ (_03695_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or _35176_ (_03696_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and _35177_ (_03697_, _03696_, _03695_);
  and _35178_ (_03698_, _03697_, _02445_);
  or _35179_ (_03699_, _03698_, _03694_);
  or _35180_ (_03700_, _03699_, _02459_);
  or _35181_ (_03702_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or _35182_ (_03704_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and _35183_ (_03705_, _03704_, _03702_);
  and _35184_ (_03706_, _03705_, _02393_);
  or _35185_ (_03707_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or _35186_ (_03708_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and _35187_ (_03709_, _03708_, _03707_);
  and _35188_ (_03711_, _03709_, _02445_);
  or _35189_ (_03712_, _03711_, _03706_);
  or _35190_ (_03714_, _03712_, _02421_);
  and _35191_ (_03715_, _03714_, _02414_);
  and _35192_ (_03716_, _03715_, _03700_);
  or _35193_ (_03717_, _03716_, _03690_);
  and _35194_ (_03718_, _03717_, _02398_);
  and _35195_ (_03719_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and _35196_ (_03720_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or _35197_ (_03721_, _03720_, _03719_);
  and _35198_ (_03722_, _03721_, _02393_);
  and _35199_ (_03723_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and _35200_ (_03725_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or _35201_ (_03726_, _03725_, _03723_);
  and _35202_ (_03727_, _03726_, _02445_);
  or _35203_ (_03728_, _03727_, _03722_);
  or _35204_ (_03729_, _03728_, _02459_);
  and _35205_ (_03730_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and _35206_ (_03731_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or _35207_ (_03732_, _03731_, _03730_);
  and _35208_ (_03733_, _03732_, _02393_);
  and _35209_ (_03734_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and _35210_ (_03735_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or _35211_ (_03736_, _03735_, _03734_);
  and _35212_ (_03737_, _03736_, _02445_);
  or _35213_ (_03738_, _03737_, _03733_);
  or _35214_ (_03739_, _03738_, _02421_);
  and _35215_ (_03740_, _03739_, _02458_);
  and _35216_ (_03741_, _03740_, _03729_);
  or _35217_ (_03743_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or _35218_ (_03744_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and _35219_ (_03745_, _03744_, _02445_);
  and _35220_ (_03746_, _03745_, _03743_);
  or _35221_ (_03747_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or _35222_ (_03749_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and _35223_ (_03750_, _03749_, _02393_);
  and _35224_ (_03752_, _03750_, _03747_);
  or _35225_ (_03753_, _03752_, _03746_);
  or _35226_ (_03754_, _03753_, _02459_);
  or _35227_ (_03755_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or _35228_ (_03756_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and _35229_ (_03757_, _03756_, _02445_);
  and _35230_ (_03758_, _03757_, _03755_);
  or _35231_ (_03759_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or _35232_ (_03760_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and _35233_ (_03761_, _03760_, _02393_);
  and _35234_ (_03762_, _03761_, _03759_);
  or _35235_ (_03764_, _03762_, _03758_);
  or _35236_ (_03766_, _03764_, _02421_);
  and _35237_ (_03767_, _03766_, _02414_);
  and _35238_ (_03769_, _03767_, _03754_);
  or _35239_ (_03770_, _03769_, _03741_);
  and _35240_ (_03771_, _03770_, _02496_);
  or _35241_ (_03772_, _03771_, _03718_);
  and _35242_ (_03773_, _03772_, _02546_);
  or _35243_ (_03774_, _03773_, _03665_);
  and _35244_ (_03776_, _03774_, _02405_);
  or _35245_ (_03777_, _03776_, _03562_);
  and _35246_ (_03778_, _03777_, _26777_);
  and _35247_ (_03779_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  and _35248_ (_03780_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or _35249_ (_03781_, _03780_, _03779_);
  and _35250_ (_03782_, _03781_, _02393_);
  and _35251_ (_03783_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and _35252_ (_03784_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or _35253_ (_03785_, _03784_, _03783_);
  and _35254_ (_03786_, _03785_, _02445_);
  or _35255_ (_03787_, _03786_, _03782_);
  and _35256_ (_03789_, _03787_, _02421_);
  and _35257_ (_03790_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  and _35258_ (_03791_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or _35259_ (_03793_, _03791_, _03790_);
  and _35260_ (_03794_, _03793_, _02393_);
  and _35261_ (_03795_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  and _35262_ (_03796_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or _35263_ (_03797_, _03796_, _03795_);
  and _35264_ (_03798_, _03797_, _02445_);
  or _35265_ (_03799_, _03798_, _03794_);
  and _35266_ (_03800_, _03799_, _02459_);
  or _35267_ (_03801_, _03800_, _03789_);
  and _35268_ (_03803_, _03801_, _02458_);
  or _35269_ (_03804_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or _35270_ (_03805_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  and _35271_ (_03806_, _03805_, _03804_);
  and _35272_ (_03807_, _03806_, _02393_);
  or _35273_ (_03808_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or _35274_ (_03810_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and _35275_ (_03811_, _03810_, _03808_);
  and _35276_ (_03812_, _03811_, _02445_);
  or _35277_ (_03813_, _03812_, _03807_);
  and _35278_ (_03814_, _03813_, _02421_);
  or _35279_ (_03815_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or _35280_ (_03816_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  and _35281_ (_03817_, _03816_, _03815_);
  and _35282_ (_03818_, _03817_, _02393_);
  or _35283_ (_03819_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or _35284_ (_03820_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and _35285_ (_03821_, _03820_, _03819_);
  and _35286_ (_03823_, _03821_, _02445_);
  or _35287_ (_03824_, _03823_, _03818_);
  and _35288_ (_03825_, _03824_, _02459_);
  or _35289_ (_03826_, _03825_, _03814_);
  and _35290_ (_03827_, _03826_, _02414_);
  or _35291_ (_03828_, _03827_, _03803_);
  and _35292_ (_03829_, _03828_, _02398_);
  and _35293_ (_03830_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and _35294_ (_03831_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or _35295_ (_03832_, _03831_, _03830_);
  and _35296_ (_03833_, _03832_, _02393_);
  and _35297_ (_03834_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and _35298_ (_03835_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or _35299_ (_03836_, _03835_, _03834_);
  and _35300_ (_03837_, _03836_, _02445_);
  or _35301_ (_03838_, _03837_, _03833_);
  and _35302_ (_03839_, _03838_, _02421_);
  and _35303_ (_03840_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and _35304_ (_03841_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _35305_ (_03842_, _03841_, _03840_);
  and _35306_ (_03843_, _03842_, _02393_);
  and _35307_ (_03844_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and _35308_ (_03845_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _35309_ (_03847_, _03845_, _03844_);
  and _35310_ (_03848_, _03847_, _02445_);
  or _35311_ (_03850_, _03848_, _03843_);
  and _35312_ (_03851_, _03850_, _02459_);
  or _35313_ (_03852_, _03851_, _03839_);
  and _35314_ (_03853_, _03852_, _02458_);
  or _35315_ (_03854_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or _35316_ (_03856_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and _35317_ (_03857_, _03856_, _02445_);
  and _35318_ (_03858_, _03857_, _03854_);
  or _35319_ (_03859_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _35320_ (_03860_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and _35321_ (_03861_, _03860_, _02393_);
  and _35322_ (_03862_, _03861_, _03859_);
  or _35323_ (_03863_, _03862_, _03858_);
  and _35324_ (_03864_, _03863_, _02421_);
  or _35325_ (_03866_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or _35326_ (_03867_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and _35327_ (_03868_, _03867_, _02445_);
  and _35328_ (_03869_, _03868_, _03866_);
  or _35329_ (_03870_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or _35330_ (_03872_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and _35331_ (_03873_, _03872_, _02393_);
  and _35332_ (_03874_, _03873_, _03870_);
  or _35333_ (_03875_, _03874_, _03869_);
  and _35334_ (_03876_, _03875_, _02459_);
  or _35335_ (_03877_, _03876_, _03864_);
  and _35336_ (_03879_, _03877_, _02414_);
  or _35337_ (_03881_, _03879_, _03853_);
  and _35338_ (_03882_, _03881_, _02496_);
  or _35339_ (_03884_, _03882_, _03829_);
  and _35340_ (_03885_, _03884_, _02400_);
  and _35341_ (_03886_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and _35342_ (_03887_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or _35343_ (_03888_, _03887_, _03886_);
  and _35344_ (_03889_, _03888_, _02393_);
  and _35345_ (_03890_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and _35346_ (_03891_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or _35347_ (_03892_, _03891_, _03890_);
  and _35348_ (_03893_, _03892_, _02445_);
  or _35349_ (_03895_, _03893_, _03889_);
  or _35350_ (_03896_, _03895_, _02459_);
  and _35351_ (_03897_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and _35352_ (_03898_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or _35353_ (_03899_, _03898_, _03897_);
  and _35354_ (_03900_, _03899_, _02393_);
  and _35355_ (_03901_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and _35356_ (_03902_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or _35357_ (_03903_, _03902_, _03901_);
  and _35358_ (_03904_, _03903_, _02445_);
  or _35359_ (_03905_, _03904_, _03900_);
  or _35360_ (_03906_, _03905_, _02421_);
  and _35361_ (_03907_, _03906_, _02458_);
  and _35362_ (_03908_, _03907_, _03896_);
  or _35363_ (_03909_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or _35364_ (_03910_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and _35365_ (_03911_, _03910_, _02445_);
  and _35366_ (_03912_, _03911_, _03909_);
  or _35367_ (_03913_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or _35368_ (_03914_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and _35369_ (_03915_, _03914_, _02393_);
  and _35370_ (_03916_, _03915_, _03913_);
  or _35371_ (_03917_, _03916_, _03912_);
  or _35372_ (_03918_, _03917_, _02459_);
  or _35373_ (_03919_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or _35374_ (_03920_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and _35375_ (_03921_, _03920_, _02445_);
  and _35376_ (_03922_, _03921_, _03919_);
  or _35377_ (_03923_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or _35378_ (_03924_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and _35379_ (_03925_, _03924_, _02393_);
  and _35380_ (_03926_, _03925_, _03923_);
  or _35381_ (_03927_, _03926_, _03922_);
  or _35382_ (_03928_, _03927_, _02421_);
  and _35383_ (_03929_, _03928_, _02414_);
  and _35384_ (_03930_, _03929_, _03918_);
  or _35385_ (_03931_, _03930_, _03908_);
  and _35386_ (_03932_, _03931_, _02496_);
  and _35387_ (_03933_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and _35388_ (_03934_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or _35389_ (_03935_, _03934_, _03933_);
  and _35390_ (_03937_, _03935_, _02393_);
  and _35391_ (_03938_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and _35392_ (_03939_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or _35393_ (_03940_, _03939_, _03938_);
  and _35394_ (_03941_, _03940_, _02445_);
  or _35395_ (_03942_, _03941_, _03937_);
  or _35396_ (_03943_, _03942_, _02459_);
  and _35397_ (_03944_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and _35398_ (_03945_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or _35399_ (_03946_, _03945_, _03944_);
  and _35400_ (_03947_, _03946_, _02393_);
  and _35401_ (_03948_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and _35402_ (_03949_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or _35403_ (_03950_, _03949_, _03948_);
  and _35404_ (_03951_, _03950_, _02445_);
  or _35405_ (_03952_, _03951_, _03947_);
  or _35406_ (_03953_, _03952_, _02421_);
  and _35407_ (_03954_, _03953_, _02458_);
  and _35408_ (_03955_, _03954_, _03943_);
  or _35409_ (_03956_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or _35410_ (_03957_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and _35411_ (_03958_, _03957_, _03956_);
  and _35412_ (_03959_, _03958_, _02393_);
  or _35413_ (_03960_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or _35414_ (_03961_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and _35415_ (_03962_, _03961_, _03960_);
  and _35416_ (_03963_, _03962_, _02445_);
  or _35417_ (_03964_, _03963_, _03959_);
  or _35418_ (_03965_, _03964_, _02459_);
  or _35419_ (_03966_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or _35420_ (_03967_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  and _35421_ (_03968_, _03967_, _03966_);
  and _35422_ (_03970_, _03968_, _02393_);
  or _35423_ (_03971_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or _35424_ (_03972_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and _35425_ (_03973_, _03972_, _03971_);
  and _35426_ (_03974_, _03973_, _02445_);
  or _35427_ (_03975_, _03974_, _03970_);
  or _35428_ (_03976_, _03975_, _02421_);
  and _35429_ (_03977_, _03976_, _02414_);
  and _35430_ (_03978_, _03977_, _03965_);
  or _35431_ (_03979_, _03978_, _03955_);
  and _35432_ (_03981_, _03979_, _02398_);
  or _35433_ (_03982_, _03981_, _03932_);
  and _35434_ (_03983_, _03982_, _02546_);
  or _35435_ (_03985_, _03983_, _03885_);
  and _35436_ (_03986_, _03985_, _02646_);
  or _35437_ (_03988_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or _35438_ (_03989_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and _35439_ (_03990_, _03989_, _02445_);
  and _35440_ (_03991_, _03990_, _03988_);
  or _35441_ (_03992_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or _35442_ (_03993_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and _35443_ (_03994_, _03993_, _02393_);
  and _35444_ (_03996_, _03994_, _03992_);
  or _35445_ (_03998_, _03996_, _03991_);
  and _35446_ (_03999_, _03998_, _02459_);
  or _35447_ (_04000_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or _35448_ (_04001_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and _35449_ (_04002_, _04001_, _02445_);
  and _35450_ (_04004_, _04002_, _04000_);
  or _35451_ (_04005_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or _35452_ (_04006_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and _35453_ (_04008_, _04006_, _02393_);
  and _35454_ (_04009_, _04008_, _04005_);
  or _35455_ (_04010_, _04009_, _04004_);
  and _35456_ (_04011_, _04010_, _02421_);
  or _35457_ (_04012_, _04011_, _03999_);
  and _35458_ (_04013_, _04012_, _02414_);
  and _35459_ (_04014_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and _35460_ (_04015_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or _35461_ (_04016_, _04015_, _04014_);
  and _35462_ (_04017_, _04016_, _02393_);
  and _35463_ (_04018_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and _35464_ (_04019_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or _35465_ (_04020_, _04019_, _04018_);
  and _35466_ (_04021_, _04020_, _02445_);
  or _35467_ (_04022_, _04021_, _04017_);
  and _35468_ (_04023_, _04022_, _02459_);
  and _35469_ (_04024_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and _35470_ (_04026_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or _35471_ (_04027_, _04026_, _04024_);
  and _35472_ (_04028_, _04027_, _02393_);
  and _35473_ (_04029_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and _35474_ (_04030_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or _35475_ (_04032_, _04030_, _04029_);
  and _35476_ (_04034_, _04032_, _02445_);
  or _35477_ (_04035_, _04034_, _04028_);
  and _35478_ (_04036_, _04035_, _02421_);
  or _35479_ (_04037_, _04036_, _04023_);
  and _35480_ (_04038_, _04037_, _02458_);
  or _35481_ (_04039_, _04038_, _04013_);
  and _35482_ (_04040_, _04039_, _02496_);
  or _35483_ (_04041_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or _35484_ (_04042_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and _35485_ (_04043_, _04042_, _04041_);
  and _35486_ (_04044_, _04043_, _02393_);
  or _35487_ (_04046_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or _35488_ (_04047_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  and _35489_ (_04048_, _04047_, _04046_);
  and _35490_ (_04050_, _04048_, _02445_);
  or _35491_ (_04051_, _04050_, _04044_);
  and _35492_ (_04052_, _04051_, _02459_);
  or _35493_ (_04053_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or _35494_ (_04054_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and _35495_ (_04055_, _04054_, _04053_);
  and _35496_ (_04056_, _04055_, _02393_);
  or _35497_ (_04057_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or _35498_ (_04058_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and _35499_ (_04059_, _04058_, _04057_);
  and _35500_ (_04060_, _04059_, _02445_);
  or _35501_ (_04061_, _04060_, _04056_);
  and _35502_ (_04062_, _04061_, _02421_);
  or _35503_ (_04063_, _04062_, _04052_);
  and _35504_ (_04064_, _04063_, _02414_);
  and _35505_ (_04065_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and _35506_ (_04066_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or _35507_ (_04067_, _04066_, _04065_);
  and _35508_ (_04068_, _04067_, _02393_);
  and _35509_ (_04069_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and _35510_ (_04070_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or _35511_ (_04071_, _04070_, _04069_);
  and _35512_ (_04072_, _04071_, _02445_);
  or _35513_ (_04073_, _04072_, _04068_);
  and _35514_ (_04074_, _04073_, _02459_);
  and _35515_ (_04075_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and _35516_ (_04076_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or _35517_ (_04077_, _04076_, _04075_);
  and _35518_ (_04078_, _04077_, _02393_);
  and _35519_ (_04079_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  and _35520_ (_04081_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or _35521_ (_04082_, _04081_, _04079_);
  and _35522_ (_04083_, _04082_, _02445_);
  or _35523_ (_04084_, _04083_, _04078_);
  and _35524_ (_04085_, _04084_, _02421_);
  or _35525_ (_04086_, _04085_, _04074_);
  and _35526_ (_04087_, _04086_, _02458_);
  or _35527_ (_04088_, _04087_, _04064_);
  and _35528_ (_04089_, _04088_, _02398_);
  or _35529_ (_04091_, _04089_, _04040_);
  and _35530_ (_04092_, _04091_, _02400_);
  and _35531_ (_04093_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and _35532_ (_04094_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or _35533_ (_04095_, _04094_, _04093_);
  and _35534_ (_04096_, _04095_, _02393_);
  and _35535_ (_04097_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and _35536_ (_04099_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or _35537_ (_04100_, _04099_, _04097_);
  and _35538_ (_04101_, _04100_, _02445_);
  or _35539_ (_04102_, _04101_, _04096_);
  or _35540_ (_04103_, _04102_, _02459_);
  and _35541_ (_04104_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and _35542_ (_04105_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or _35543_ (_04106_, _04105_, _04104_);
  and _35544_ (_04107_, _04106_, _02393_);
  and _35545_ (_04108_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and _35546_ (_04109_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or _35547_ (_04110_, _04109_, _04108_);
  and _35548_ (_04112_, _04110_, _02445_);
  or _35549_ (_04113_, _04112_, _04107_);
  or _35550_ (_04115_, _04113_, _02421_);
  and _35551_ (_04116_, _04115_, _02458_);
  and _35552_ (_04118_, _04116_, _04103_);
  or _35553_ (_04119_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or _35554_ (_04121_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and _35555_ (_04122_, _04121_, _04119_);
  and _35556_ (_04123_, _04122_, _02393_);
  or _35557_ (_04124_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or _35558_ (_04126_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and _35559_ (_04127_, _04126_, _04124_);
  and _35560_ (_04128_, _04127_, _02445_);
  or _35561_ (_04129_, _04128_, _04123_);
  or _35562_ (_04130_, _04129_, _02459_);
  or _35563_ (_04131_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or _35564_ (_04132_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and _35565_ (_04134_, _04132_, _04131_);
  and _35566_ (_04135_, _04134_, _02393_);
  or _35567_ (_04136_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or _35568_ (_04137_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and _35569_ (_04138_, _04137_, _04136_);
  and _35570_ (_04139_, _04138_, _02445_);
  or _35571_ (_04141_, _04139_, _04135_);
  or _35572_ (_04142_, _04141_, _02421_);
  and _35573_ (_04143_, _04142_, _02414_);
  and _35574_ (_04144_, _04143_, _04130_);
  or _35575_ (_04145_, _04144_, _04118_);
  and _35576_ (_04146_, _04145_, _02398_);
  and _35577_ (_04147_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  and _35578_ (_04148_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or _35579_ (_04149_, _04148_, _04147_);
  and _35580_ (_04150_, _04149_, _02393_);
  and _35581_ (_04151_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and _35582_ (_04152_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or _35583_ (_04153_, _04152_, _04151_);
  and _35584_ (_04154_, _04153_, _02445_);
  or _35585_ (_04155_, _04154_, _04150_);
  or _35586_ (_04156_, _04155_, _02459_);
  and _35587_ (_04157_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and _35588_ (_04158_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or _35589_ (_04159_, _04158_, _04157_);
  and _35590_ (_04160_, _04159_, _02393_);
  and _35591_ (_04161_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  and _35592_ (_04162_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or _35593_ (_04163_, _04162_, _04161_);
  and _35594_ (_04164_, _04163_, _02445_);
  or _35595_ (_04165_, _04164_, _04160_);
  or _35596_ (_04166_, _04165_, _02421_);
  and _35597_ (_04167_, _04166_, _02458_);
  and _35598_ (_04168_, _04167_, _04156_);
  or _35599_ (_04169_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or _35600_ (_04170_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and _35601_ (_04172_, _04170_, _02445_);
  and _35602_ (_04173_, _04172_, _04169_);
  or _35603_ (_04175_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or _35604_ (_04176_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and _35605_ (_04177_, _04176_, _02393_);
  and _35606_ (_04178_, _04177_, _04175_);
  or _35607_ (_04179_, _04178_, _04173_);
  or _35608_ (_04180_, _04179_, _02459_);
  or _35609_ (_04181_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or _35610_ (_04182_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and _35611_ (_04183_, _04182_, _02445_);
  and _35612_ (_04184_, _04183_, _04181_);
  or _35613_ (_04185_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or _35614_ (_04186_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and _35615_ (_04187_, _04186_, _02393_);
  and _35616_ (_04188_, _04187_, _04185_);
  or _35617_ (_04189_, _04188_, _04184_);
  or _35618_ (_04190_, _04189_, _02421_);
  and _35619_ (_04191_, _04190_, _02414_);
  and _35620_ (_04192_, _04191_, _04180_);
  or _35621_ (_04194_, _04192_, _04168_);
  and _35622_ (_04196_, _04194_, _02496_);
  or _35623_ (_04197_, _04196_, _04146_);
  and _35624_ (_04198_, _04197_, _02546_);
  or _35625_ (_04200_, _04198_, _04092_);
  and _35626_ (_04201_, _04200_, _02405_);
  or _35627_ (_04202_, _04201_, _03986_);
  and _35628_ (_04204_, _04202_, _02444_);
  or _35629_ (_04205_, _04204_, _03778_);
  or _35630_ (_04206_, _04205_, _02443_);
  or _35631_ (_04207_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and _35632_ (_04208_, _04207_, _22762_);
  and _35633_ (_22721_, _04208_, _04206_);
  nor _35634_ (_04210_, _01772_, rst);
  nand _35635_ (_04211_, _22768_, _01532_);
  and _35636_ (_26893_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _22762_);
  and _35637_ (_04213_, _26893_, _04211_);
  or _35638_ (_26894_, _04213_, _04210_);
  and _35639_ (_04215_, _03339_, _23824_);
  and _35640_ (_04216_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or _35641_ (_27112_, _04216_, _04215_);
  and _35642_ (_04218_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  and _35643_ (_04219_, _02298_, _24050_);
  or _35644_ (_27237_, _04219_, _04218_);
  and _35645_ (_04220_, _25656_, _23824_);
  and _35646_ (_04221_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or _35647_ (_22723_, _04221_, _04220_);
  and _35648_ (_04222_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _22762_);
  and _35649_ (_04223_, _04222_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _35650_ (_04224_, _01744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _35651_ (_04226_, _01744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _35652_ (_04227_, _04226_, _04224_);
  not _35653_ (_04228_, _04227_);
  nor _35654_ (_04229_, _04228_, _01747_);
  and _35655_ (_04230_, _04228_, _01747_);
  or _35656_ (_04231_, _04230_, _04229_);
  or _35657_ (_04232_, _04231_, _25729_);
  or _35658_ (_04233_, _25728_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _35659_ (_04234_, _04233_, _01793_);
  and _35660_ (_04235_, _04234_, _04232_);
  or _35661_ (_26891_[15], _04235_, _04223_);
  and _35662_ (_04236_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  and _35663_ (_04237_, _02306_, _23898_);
  or _35664_ (_22724_, _04237_, _04236_);
  and _35665_ (_04239_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _35666_ (_04240_, _04239_, _03332_);
  and _35667_ (_04241_, _04240_, _22762_);
  and _35668_ (_04242_, _03311_, _24581_);
  or _35669_ (_04243_, _04242_, _24617_);
  or _35670_ (_04244_, _04243_, _26616_);
  and _35671_ (_04245_, _26621_, _24471_);
  or _35672_ (_04247_, _04245_, _24585_);
  or _35673_ (_04248_, _04247_, _03330_);
  or _35674_ (_04249_, _04248_, _04244_);
  and _35675_ (_04250_, _04249_, _25644_);
  or _35676_ (_26868_[1], _04250_, _04241_);
  and _35677_ (_26889_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _22762_);
  and _35678_ (_04251_, _03339_, _23778_);
  and _35679_ (_04252_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or _35680_ (_22725_, _04252_, _04251_);
  and _35681_ (_04253_, _02350_, _23707_);
  and _35682_ (_04254_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or _35683_ (_22726_, _04254_, _04253_);
  and _35684_ (_04255_, _02350_, _24050_);
  and _35685_ (_04256_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or _35686_ (_22727_, _04256_, _04255_);
  nand _35687_ (_04257_, _00886_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _35688_ (_04259_, _04257_, _01213_);
  and _35689_ (_04260_, _04259_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _35690_ (_04261_, _01216_, _23185_);
  and _35691_ (_04262_, _04261_, _23149_);
  or _35692_ (_04263_, _04262_, _04260_);
  nand _35693_ (_04264_, _04263_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or _35694_ (_04265_, _04263_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _35695_ (_04266_, _04265_, _00401_);
  and _35696_ (_04267_, _04266_, _04264_);
  and _35697_ (_04268_, _00875_, _24628_);
  nor _35698_ (_04269_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _35699_ (_04271_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23095_);
  nor _35700_ (_04272_, _04271_, _04269_);
  nor _35701_ (_04273_, _04272_, _01283_);
  and _35702_ (_04274_, _04272_, _01283_);
  or _35703_ (_04276_, _04274_, _04273_);
  and _35704_ (_04277_, _04276_, _23480_);
  or _35705_ (_04278_, _26521_, _26481_);
  and _35706_ (_04279_, _04278_, _26522_);
  and _35707_ (_04280_, _04279_, _23596_);
  and _35708_ (_04281_, _01294_, _23179_);
  nor _35709_ (_04282_, _04281_, _01293_);
  nor _35710_ (_04283_, _04282_, _01302_);
  nand _35711_ (_04284_, _04283_, _23142_);
  or _35712_ (_04285_, _04283_, _23142_);
  and _35713_ (_04286_, _04285_, _23609_);
  and _35714_ (_04287_, _04286_, _04284_);
  and _35715_ (_04288_, _23521_, _23142_);
  or _35716_ (_04289_, _04288_, _23537_);
  and _35717_ (_04290_, _04289_, _23627_);
  and _35718_ (_04291_, _00611_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _35719_ (_04292_, _23579_, _23142_);
  and _35720_ (_04293_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  or _35721_ (_04294_, _04293_, _04292_);
  or _35722_ (_04295_, _04294_, _04291_);
  or _35723_ (_04296_, _04295_, _04290_);
  or _35724_ (_04297_, _04296_, _04287_);
  or _35725_ (_04298_, _04297_, _04280_);
  or _35726_ (_04299_, _04298_, _04277_);
  and _35727_ (_04300_, _04299_, _26566_);
  nor _35728_ (_04301_, _01343_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _35729_ (_04302_, _01343_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _35730_ (_04303_, _04302_, _04301_);
  nand _35731_ (_04304_, _04303_, _01349_);
  or _35732_ (_04305_, _04303_, _01349_);
  and _35733_ (_04306_, _04305_, _04304_);
  and _35734_ (_04307_, _04306_, _00405_);
  and _35735_ (_04308_, _26573_, _26772_);
  or _35736_ (_04309_, _04308_, _04307_);
  and _35737_ (_04310_, _26611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _35738_ (_04311_, _04310_, _04309_);
  nor _35739_ (_04312_, _04311_, _04300_);
  nand _35740_ (_04313_, _04312_, _00289_);
  or _35741_ (_04314_, _04313_, _04268_);
  or _35742_ (_04315_, _04314_, _04267_);
  or _35743_ (_04316_, _04303_, _00289_);
  and _35744_ (_04317_, _04316_, _22762_);
  and _35745_ (_26890_[15], _04317_, _04315_);
  nor _35746_ (_04318_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _35747_ (_26892_, _04318_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  nor _35748_ (_04319_, _23953_, _23950_);
  and _35749_ (_04320_, _01801_, _01798_);
  nor _35750_ (_04321_, _04320_, _23950_);
  and _35751_ (_04322_, _04321_, _23840_);
  nor _35752_ (_04323_, _04321_, _23840_);
  nor _35753_ (_04324_, _04323_, _04322_);
  nor _35754_ (_04325_, _04324_, _04319_);
  and _35755_ (_04326_, _23856_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _35756_ (_04327_, _04326_, _04319_);
  and _35757_ (_04328_, _04327_, _01517_);
  or _35758_ (_04329_, _04328_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _35759_ (_04331_, _04329_, _04325_);
  and _35760_ (_26896_[2], _04331_, _22762_);
  and _35761_ (_04333_, _24812_, _24647_);
  and _35762_ (_04334_, _04333_, _24705_);
  nand _35763_ (_04335_, _04334_, _23594_);
  and _35764_ (_04336_, _25769_, _23753_);
  and _35765_ (_04337_, _04336_, _24735_);
  not _35766_ (_04339_, _04337_);
  or _35767_ (_04340_, _04334_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _35768_ (_04341_, _04340_, _04339_);
  and _35769_ (_04342_, _04341_, _04335_);
  and _35770_ (_04343_, _04337_, _24043_);
  or _35771_ (_04344_, _04343_, _04342_);
  and _35772_ (_22728_, _04344_, _22762_);
  and _35773_ (_04346_, _04333_, _24125_);
  nand _35774_ (_04347_, _04346_, _23594_);
  or _35775_ (_04348_, _04346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _35776_ (_04349_, _04348_, _04339_);
  and _35777_ (_04350_, _04349_, _04347_);
  and _35778_ (_04351_, _04337_, _23939_);
  or _35779_ (_04353_, _04351_, _04350_);
  and _35780_ (_22729_, _04353_, _22762_);
  and _35781_ (_04354_, _24746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _35782_ (_04356_, _04354_, _24745_);
  and _35783_ (_04357_, _04356_, _04333_);
  not _35784_ (_04358_, _04333_);
  or _35785_ (_04360_, _04358_, _24752_);
  and _35786_ (_04362_, _04360_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _35787_ (_04363_, _04362_, _04337_);
  or _35788_ (_04365_, _04363_, _04357_);
  or _35789_ (_04366_, _04339_, _23642_);
  and _35790_ (_04367_, _04366_, _22762_);
  and _35791_ (_22730_, _04367_, _04365_);
  and _35792_ (_04368_, _04333_, _24118_);
  nand _35793_ (_04369_, _04368_, _23594_);
  or _35794_ (_04370_, _04368_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _35795_ (_04372_, _04370_, _04339_);
  and _35796_ (_04373_, _04372_, _04369_);
  and _35797_ (_04374_, _04337_, _23738_);
  or _35798_ (_04375_, _04374_, _04373_);
  and _35799_ (_22731_, _04375_, _22762_);
  nor _35800_ (_04376_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _35801_ (_04377_, _04376_);
  nor _35802_ (_04378_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _35803_ (_04380_, _04378_, _04377_);
  and _35804_ (_04381_, _04380_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not _35805_ (_04383_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor _35806_ (_04384_, _04380_, _04383_);
  or _35807_ (_04386_, _04384_, _04381_);
  or _35808_ (_04387_, _04386_, _04333_);
  not _35809_ (_04388_, _24291_);
  nor _35810_ (_04389_, _04388_, _23594_);
  or _35811_ (_04390_, _24291_, _04383_);
  nand _35812_ (_04391_, _04390_, _04333_);
  or _35813_ (_04392_, _04391_, _04389_);
  and _35814_ (_04393_, _04392_, _04387_);
  or _35815_ (_04394_, _04393_, _04337_);
  or _35816_ (_04395_, _04339_, _23816_);
  and _35817_ (_04396_, _04395_, _22762_);
  and _35818_ (_22732_, _04396_, _04394_);
  not _35819_ (_04397_, _24067_);
  nor _35820_ (_04398_, _04397_, _23594_);
  nand _35821_ (_04399_, _04397_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _35822_ (_04401_, _04399_, _04333_);
  or _35823_ (_04402_, _04401_, _04398_);
  or _35824_ (_04403_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _35825_ (_04404_, _04403_, _04333_);
  and _35826_ (_04405_, _04404_, _04402_);
  or _35827_ (_04406_, _04405_, _04337_);
  or _35828_ (_04407_, _04339_, _23892_);
  and _35829_ (_04408_, _04407_, _22762_);
  and _35830_ (_22733_, _04408_, _04406_);
  not _35831_ (_04410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _35832_ (_04411_, _04410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _35833_ (_04413_, _04411_, _04376_);
  and _35834_ (_04414_, _04413_, _04378_);
  or _35835_ (_04415_, _04414_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _35836_ (_04417_, _04415_, _04333_);
  and _35837_ (_04418_, _24678_, _23711_);
  not _35838_ (_04420_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _35839_ (_04421_, _24678_, _04420_);
  nand _35840_ (_04423_, _04421_, _04333_);
  or _35841_ (_04424_, _04423_, _04418_);
  and _35842_ (_04425_, _04424_, _04417_);
  or _35843_ (_04426_, _04425_, _04337_);
  nand _35844_ (_04427_, _04337_, _23772_);
  and _35845_ (_04428_, _04427_, _22762_);
  and _35846_ (_22734_, _04428_, _04426_);
  or _35847_ (_04429_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _35848_ (_04430_, _04429_, _22762_);
  or _35849_ (_04431_, _02037_, _24043_);
  and _35850_ (_22735_, _04431_, _04430_);
  or _35851_ (_04432_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _35852_ (_04433_, _04432_, _22762_);
  or _35853_ (_04434_, _02037_, _23939_);
  and _35854_ (_22736_, _04434_, _04433_);
  or _35855_ (_04435_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _35856_ (_04436_, _04435_, _22762_);
  or _35857_ (_04437_, _02037_, _23738_);
  and _35858_ (_22737_, _04437_, _04436_);
  or _35859_ (_04438_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _35860_ (_04439_, _04438_, _22762_);
  or _35861_ (_04440_, _02037_, _23892_);
  and _35862_ (_22738_, _04440_, _04439_);
  nand _35863_ (_04441_, _02034_, _23772_);
  or _35864_ (_04442_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _35865_ (_04443_, _04442_, _22762_);
  and _35866_ (_22739_, _04443_, _04441_);
  and _35867_ (_04444_, _02350_, _23946_);
  and _35868_ (_04445_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or _35869_ (_22740_, _04445_, _04444_);
  and _35870_ (_04447_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _35871_ (_04448_, _04447_, _04376_);
  and _35872_ (_04449_, _04377_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _35873_ (_04451_, _04449_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _35874_ (_04452_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _35875_ (_04453_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _35876_ (_04454_, _04453_, _04452_);
  and _35877_ (_04455_, _04454_, _04451_);
  nor _35878_ (_04457_, _04455_, _04448_);
  not _35879_ (_04458_, _04457_);
  and _35880_ (_04459_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _35881_ (_04460_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor _35882_ (_04461_, _04460_, _04459_);
  and _35883_ (_04462_, _04336_, _24072_);
  nor _35884_ (_04463_, _04462_, _04461_);
  not _35885_ (_04464_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _35886_ (_04465_, _04464_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _35887_ (_04466_, _04465_, _04377_);
  and _35888_ (_04467_, _04466_, _04462_);
  or _35889_ (_04469_, _04467_, _04463_);
  and _35890_ (_22741_, _04469_, _22762_);
  and _35891_ (_04470_, _04462_, _04377_);
  nand _35892_ (_04471_, _04470_, _23702_);
  and _35893_ (_04473_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _35894_ (_04474_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _35895_ (_04475_, _04474_, _04473_);
  or _35896_ (_04476_, _04475_, _04462_);
  and _35897_ (_04477_, _04476_, _22762_);
  and _35898_ (_22742_, _04477_, _04471_);
  and _35899_ (_04478_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _35900_ (_04479_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor _35901_ (_04480_, _04479_, _04478_);
  nor _35902_ (_04481_, _04480_, _04462_);
  and _35903_ (_04483_, _04470_, _24043_);
  or _35904_ (_04484_, _04483_, _04481_);
  and _35905_ (_04485_, _04462_, _04376_);
  and _35906_ (_04486_, _04485_, _26750_);
  or _35907_ (_04487_, _04486_, _04484_);
  and _35908_ (_22743_, _04487_, _22762_);
  not _35909_ (_04488_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _35910_ (_04490_, _04462_, _04464_);
  and _35911_ (_04491_, _04490_, _04488_);
  and _35912_ (_04493_, _04491_, _24043_);
  and _35913_ (_04494_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _35914_ (_04495_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor _35915_ (_04496_, _04495_, _04494_);
  nor _35916_ (_04497_, _04496_, _04462_);
  and _35917_ (_04498_, _04470_, _23939_);
  or _35918_ (_04500_, _04498_, _04497_);
  or _35919_ (_04501_, _04500_, _04493_);
  and _35920_ (_22744_, _04501_, _22762_);
  and _35921_ (_04504_, _04491_, _23939_);
  and _35922_ (_04505_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _35923_ (_04506_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor _35924_ (_04507_, _04506_, _04505_);
  nor _35925_ (_04508_, _04507_, _04462_);
  and _35926_ (_04509_, _04470_, _23642_);
  or _35927_ (_04510_, _04509_, _04508_);
  or _35928_ (_04511_, _04510_, _04504_);
  and _35929_ (_22745_, _04511_, _22762_);
  and _35930_ (_04513_, _04491_, _23642_);
  and _35931_ (_04514_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _35932_ (_04515_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _35933_ (_04516_, _04515_, _04514_);
  nor _35934_ (_04517_, _04516_, _04462_);
  and _35935_ (_04518_, _04470_, _23738_);
  or _35936_ (_04520_, _04518_, _04517_);
  or _35937_ (_04521_, _04520_, _04513_);
  and _35938_ (_22747_, _04521_, _22762_);
  and _35939_ (_04522_, _04470_, _23816_);
  and _35940_ (_04523_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and _35941_ (_04524_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _35942_ (_04525_, _04524_, _04523_);
  nor _35943_ (_04526_, _04525_, _04462_);
  and _35944_ (_04527_, _04491_, _23738_);
  or _35945_ (_04528_, _04527_, _04526_);
  or _35946_ (_04529_, _04528_, _04522_);
  and _35947_ (_22748_, _04529_, _22762_);
  and _35948_ (_04531_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _35949_ (_04532_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor _35950_ (_04533_, _04532_, _04531_);
  nor _35951_ (_04535_, _04533_, _04462_);
  and _35952_ (_04536_, _04470_, _23892_);
  or _35953_ (_04537_, _04536_, _04535_);
  and _35954_ (_04538_, _04485_, _23816_);
  or _35955_ (_04540_, _04538_, _04537_);
  and _35956_ (_22749_, _04540_, _22762_);
  and _35957_ (_04541_, _04491_, _23892_);
  and _35958_ (_04543_, _04458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _35959_ (_04544_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor _35960_ (_04545_, _04544_, _04543_);
  nor _35961_ (_04547_, _04545_, _04462_);
  and _35962_ (_04549_, _04470_, _24685_);
  or _35963_ (_04551_, _04549_, _04547_);
  or _35964_ (_04552_, _04551_, _04541_);
  and _35965_ (_22750_, _04552_, _22762_);
  or _35966_ (_04554_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _35967_ (_04555_, _04448_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _35968_ (_04556_, _04555_, _04455_);
  and _35969_ (_04557_, _04556_, _04554_);
  nor _35970_ (_04558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nor _35971_ (_04559_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _35972_ (_04560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _35973_ (_04561_, _04560_, _04559_);
  and _35974_ (_04563_, _04561_, _04558_);
  nor _35975_ (_04564_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _35976_ (_04565_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _35977_ (_04567_, _04565_, _04564_);
  and _35978_ (_04568_, _04567_, _04448_);
  and _35979_ (_04569_, _04568_, _04563_);
  and _35980_ (_04570_, _04569_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor _35981_ (_04571_, _04570_, _04557_);
  nor _35982_ (_04572_, _04571_, _04462_);
  and _35983_ (_04574_, _04485_, _24685_);
  or _35984_ (_04575_, _04574_, _04572_);
  and _35985_ (_22751_, _04575_, _22762_);
  not _35986_ (_04576_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor _35987_ (_04578_, _04376_, _04576_);
  and _35988_ (_04579_, _04578_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _35989_ (_04581_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _35990_ (_04582_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _04581_);
  not _35991_ (_04584_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _35992_ (_04586_, _04584_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _35993_ (_04588_, _04586_, _04582_);
  and _35994_ (_04589_, _04588_, _04579_);
  and _35995_ (_04591_, _04576_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _35996_ (_04593_, _04376_, _04420_);
  and _35997_ (_04594_, _04593_, _04591_);
  and _35998_ (_04595_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _35999_ (_04596_, _04595_, _04377_);
  nor _36000_ (_04598_, _04596_, _04594_);
  nor _36001_ (_04599_, _04598_, _04579_);
  or _36002_ (_04600_, _04599_, _04589_);
  and _36003_ (_04601_, _04376_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _36004_ (_04602_, _04601_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or _36005_ (_04603_, _04602_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _36006_ (_04604_, _04603_, _04600_);
  nor _36007_ (_04605_, _04602_, _04589_);
  or _36008_ (_04606_, _04605_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _36009_ (_04607_, _04606_, _02066_);
  and _36010_ (_04608_, _04607_, _04604_);
  or _36011_ (_22752_, _04608_, _02065_);
  not _36012_ (_04609_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  not _36013_ (_04611_, _04605_);
  nor _36014_ (_04612_, _04611_, _04599_);
  nor _36015_ (_04613_, _04612_, _04609_);
  or _36016_ (_04615_, _04613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _36017_ (_04616_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _04609_);
  or _36018_ (_04618_, _04616_, _04605_);
  and _36019_ (_04619_, _04618_, _22762_);
  and _36020_ (_22753_, _04619_, _04615_);
  and _36021_ (_04621_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  and _36022_ (_04623_, _02245_, _23946_);
  or _36023_ (_22754_, _04623_, _04621_);
  and _36024_ (_04625_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _36025_ (_04627_, _04611_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  not _36026_ (_04628_, _04579_);
  nor _36027_ (_04629_, _04588_, _04628_);
  and _36028_ (_04630_, _04629_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _36029_ (_04631_, _04596_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nand _36030_ (_04632_, _04631_, _04628_);
  nor _36031_ (_04633_, _04632_, _04594_);
  nor _36032_ (_04634_, _04633_, _04630_);
  nor _36033_ (_04636_, _04634_, _04602_);
  or _36034_ (_04637_, _04636_, _04627_);
  and _36035_ (_04639_, _04637_, _02066_);
  or _36036_ (_22755_, _04639_, _04625_);
  and _36037_ (_04641_, _01810_, _23946_);
  and _36038_ (_04643_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or _36039_ (_22756_, _04643_, _04641_);
  and _36040_ (_04644_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  and _36041_ (_04646_, _02245_, _23649_);
  or _36042_ (_27036_, _04646_, _04644_);
  and _36043_ (_04648_, _25656_, _23649_);
  and _36044_ (_04650_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or _36045_ (_27192_, _04650_, _04648_);
  and _36046_ (_04652_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  and _36047_ (_04654_, _02298_, _23707_);
  or _36048_ (_27238_, _04654_, _04652_);
  and _36049_ (_04656_, _01758_, _23986_);
  and _36050_ (_04658_, _04656_, _23707_);
  not _36051_ (_04660_, _04656_);
  and _36052_ (_04661_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or _36053_ (_22758_, _04661_, _04658_);
  and _36054_ (_04663_, _01478_, _01377_);
  or _36055_ (_04665_, _04663_, _01474_);
  and _36056_ (_04666_, _01487_, _01383_);
  and _36057_ (_04667_, _01426_, _01362_);
  or _36058_ (_04668_, _04667_, _04666_);
  or _36059_ (_04669_, _04668_, _04665_);
  and _36060_ (_04671_, _01422_, _01357_);
  and _36061_ (_04673_, _01472_, _01425_);
  and _36062_ (_04674_, _01368_, _01362_);
  or _36063_ (_04675_, _04674_, _04673_);
  or _36064_ (_04676_, _04675_, _04671_);
  or _36065_ (_04677_, _01509_, _01491_);
  or _36066_ (_04678_, _04677_, _01380_);
  or _36067_ (_04679_, _04678_, _04676_);
  or _36068_ (_04680_, _04679_, _04669_);
  and _36069_ (_04681_, _01461_, _01401_);
  and _36070_ (_04682_, _01401_, _01395_);
  or _36071_ (_04683_, _01453_, _01376_);
  and _36072_ (_04684_, _04683_, _01426_);
  or _36073_ (_04685_, _04684_, _04682_);
  nor _36074_ (_04686_, _04685_, _04681_);
  nand _36075_ (_04688_, _04686_, _01436_);
  or _36076_ (_04690_, _04688_, _04680_);
  and _36077_ (_04691_, _04690_, _22769_);
  and _36078_ (_04693_, _22765_, _22766_);
  and _36079_ (_04694_, _04693_, _24564_);
  nor _36080_ (_04695_, _04694_, _25661_);
  or _36081_ (_04696_, _04695_, rst);
  or _36082_ (_26863_[1], _04696_, _04691_);
  and _36083_ (_04698_, _04656_, _24050_);
  and _36084_ (_04700_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or _36085_ (_22759_, _04700_, _04698_);
  not _36086_ (_04701_, _04612_);
  or _36087_ (_04702_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _36088_ (_04703_, _04605_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _36089_ (_04704_, _04703_, _02066_);
  and _36090_ (_04705_, _04704_, _04702_);
  or _36091_ (_22760_, _04705_, _02071_);
  and _36092_ (_04706_, _02370_, _23824_);
  and _36093_ (_04707_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or _36094_ (_22761_, _04707_, _04706_);
  and _36095_ (_04708_, _02200_, _23778_);
  and _36096_ (_04709_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or _36097_ (_22774_, _04709_, _04708_);
  and _36098_ (_04711_, _04588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _36099_ (_04712_, _04711_, _04598_);
  or _36100_ (_04714_, _04712_, _04612_);
  and _36101_ (_04715_, _04714_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _36102_ (_04717_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _04609_);
  nand _36103_ (_04718_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _36104_ (_04720_, _04718_, _04605_);
  or _36105_ (_04721_, _04720_, _04717_);
  or _36106_ (_04723_, _04721_, _04715_);
  and _36107_ (_22776_, _04723_, _22762_);
  nor _36108_ (_04724_, _04596_, _04579_);
  or _36109_ (_04725_, _04724_, _04609_);
  or _36110_ (_04726_, _04725_, _04584_);
  and _36111_ (_04727_, _04579_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _36112_ (_04728_, _04727_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _36113_ (_04729_, _04728_, _22762_);
  and _36114_ (_22779_, _04729_, _04726_);
  and _36115_ (_04730_, _24331_, _24050_);
  and _36116_ (_04732_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or _36117_ (_22787_, _04732_, _04730_);
  nand _36118_ (_04734_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22762_);
  nor _36119_ (_04735_, _04734_, _04613_);
  or _36120_ (_04736_, _04712_, _04611_);
  and _36121_ (_04737_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _36122_ (_04738_, _04737_, _04736_);
  or _36123_ (_22790_, _04738_, _04735_);
  and _36124_ (_04740_, _04725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _36125_ (_04741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _36126_ (_04743_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _36127_ (_04744_, _04743_, _04741_);
  and _36128_ (_04745_, _04744_, _04727_);
  or _36129_ (_04746_, _04745_, _04740_);
  and _36130_ (_22792_, _04746_, _22762_);
  and _36131_ (_04748_, _01808_, _24766_);
  not _36132_ (_04749_, _04748_);
  and _36133_ (_04751_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  and _36134_ (_04752_, _04748_, _23707_);
  or _36135_ (_22818_, _04752_, _04751_);
  or _36136_ (_04754_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _36137_ (_04756_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _36138_ (_04757_, _04756_, rst);
  nand _36139_ (_04758_, _04757_, _04754_);
  nor _36140_ (_22831_, _04758_, _04462_);
  and _36141_ (_04760_, _23788_, _23072_);
  and _36142_ (_04761_, _04760_, _01808_);
  not _36143_ (_04762_, _04761_);
  and _36144_ (_04763_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and _36145_ (_04764_, _04761_, _23649_);
  or _36146_ (_22835_, _04764_, _04763_);
  and _36147_ (_04766_, _04741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _36148_ (_04767_, _04766_, _04581_);
  and _36149_ (_04768_, _04727_, _04767_);
  or _36150_ (_04769_, _04768_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not _36151_ (_04770_, rxd_i);
  nand _36152_ (_04771_, _04768_, _04770_);
  and _36153_ (_04772_, _04771_, _22762_);
  and _36154_ (_22851_, _04772_, _04769_);
  or _36155_ (_04773_, _04756_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _36156_ (_04774_, _04756_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _36157_ (_04775_, _04774_, rst);
  nand _36158_ (_04776_, _04775_, _04773_);
  nor _36159_ (_22856_, _04776_, _04462_);
  nor _36160_ (_04778_, _04774_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and _36161_ (_04780_, _04774_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _36162_ (_04781_, _04780_, _04778_);
  nand _36163_ (_04782_, _04781_, _22762_);
  nor _36164_ (_22858_, _04782_, _04462_);
  and _36165_ (_04783_, _02350_, _23898_);
  and _36166_ (_04785_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or _36167_ (_22863_, _04785_, _04783_);
  and _36168_ (_04786_, _24006_, _23747_);
  and _36169_ (_04787_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  or _36170_ (_22866_, _04787_, _04786_);
  or _36171_ (_04788_, _04613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _36172_ (_04789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _04609_);
  or _36173_ (_04790_, _04789_, _04605_);
  and _36174_ (_04791_, _04790_, _22762_);
  and _36175_ (_22873_, _04791_, _04788_);
  and _36176_ (_04792_, _02350_, _23778_);
  and _36177_ (_04793_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or _36178_ (_22880_, _04793_, _04792_);
  and _36179_ (_04794_, _01971_, _23824_);
  and _36180_ (_04795_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  or _36181_ (_22898_, _04795_, _04794_);
  and _36182_ (_04797_, _01809_, _23069_);
  and _36183_ (_04799_, _04797_, _23824_);
  not _36184_ (_04800_, _04797_);
  and _36185_ (_04801_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or _36186_ (_22902_, _04801_, _04799_);
  and _36187_ (_04804_, _04725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor _36188_ (_04805_, _04766_, _04628_);
  or _36189_ (_04806_, _04805_, _04804_);
  and _36190_ (_04807_, _04741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _36191_ (_04809_, _04807_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _36192_ (_04810_, _04809_, _22762_);
  and _36193_ (_22911_, _04810_, _04806_);
  and _36194_ (_04811_, _23754_, _23069_);
  and _36195_ (_04812_, _04811_, _23946_);
  not _36196_ (_04813_, _04811_);
  and _36197_ (_04814_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  or _36198_ (_22916_, _04814_, _04812_);
  and _36199_ (_04816_, _24699_, _23649_);
  and _36200_ (_04817_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  or _36201_ (_22925_, _04817_, _04816_);
  and _36202_ (_04819_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _36203_ (_22933_, _04819_, _04625_);
  and _36204_ (_04820_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and _36205_ (_04821_, _02245_, _23778_);
  or _36206_ (_22936_, _04821_, _04820_);
  and _36207_ (_04822_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _36208_ (_04823_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _36209_ (_22955_, _04823_, _04822_);
  and _36210_ (_04825_, _04656_, _23778_);
  and _36211_ (_04826_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or _36212_ (_22959_, _04826_, _04825_);
  and _36213_ (_04828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _36214_ (_04829_, _04828_, _04717_);
  and _36215_ (_22965_, _04829_, _22762_);
  and _36216_ (_04830_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _36217_ (_04831_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or _36218_ (_22988_, _04831_, _04830_);
  and _36219_ (_04832_, _01758_, _23069_);
  and _36220_ (_04833_, _04832_, _23707_);
  not _36221_ (_04834_, _04832_);
  and _36222_ (_04835_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or _36223_ (_22993_, _04835_, _04833_);
  and _36224_ (_04836_, _03300_, _23824_);
  and _36225_ (_04838_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or _36226_ (_22998_, _04838_, _04836_);
  or _36227_ (_04839_, _04613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _36228_ (_04840_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _04609_);
  or _36229_ (_04842_, _04840_, _04605_);
  and _36230_ (_04843_, _04842_, _22762_);
  and _36231_ (_23001_, _04843_, _04839_);
  or _36232_ (_04845_, _04701_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _36233_ (_04846_, _04605_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _36234_ (_04848_, _04846_, _02066_);
  and _36235_ (_04850_, _04848_, _04845_);
  or _36236_ (_23007_, _04850_, _02069_);
  or _36237_ (_04852_, _04613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _36238_ (_04853_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _04609_);
  or _36239_ (_04854_, _04853_, _04605_);
  and _36240_ (_04855_, _04854_, _22762_);
  and _36241_ (_23010_, _04855_, _04852_);
  or _36242_ (_04856_, _04613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _36243_ (_04857_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _04609_);
  or _36244_ (_04858_, _04857_, _04605_);
  and _36245_ (_04859_, _04858_, _22762_);
  and _36246_ (_23013_, _04859_, _04856_);
  and _36247_ (_04860_, _26099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _36248_ (_04861_, _04860_, _26100_);
  not _36249_ (_04862_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _36250_ (_04863_, _26117_, _26114_);
  and _36251_ (_04864_, _04863_, _26110_);
  and _36252_ (_04866_, _04864_, _24308_);
  and _36253_ (_04867_, _04866_, _26099_);
  nor _36254_ (_04869_, _04867_, _04862_);
  and _36255_ (_04871_, _04867_, _04862_);
  or _36256_ (_04872_, _04871_, _04869_);
  and _36257_ (_04873_, _04872_, _04861_);
  and _36258_ (_04874_, _24308_, _24300_);
  and _36259_ (_04876_, _04874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _36260_ (_04877_, _04874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _36261_ (_04878_, _04877_, _24302_);
  nor _36262_ (_04879_, _04878_, _04876_);
  and _36263_ (_04880_, _26115_, _24307_);
  and _36264_ (_04881_, _04880_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _36265_ (_04882_, _04881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _36266_ (_04883_, _04881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _36267_ (_04885_, _04883_, _26097_);
  nor _36268_ (_04886_, _04885_, _04882_);
  or _36269_ (_04887_, _04886_, _04879_);
  or _36270_ (_04888_, _04887_, _04873_);
  or _36271_ (_04890_, _04888_, _24299_);
  not _36272_ (_04891_, _24299_);
  or _36273_ (_04892_, _04891_, _23738_);
  and _36274_ (_04894_, _04892_, _04890_);
  or _36275_ (_04895_, _04894_, _24293_);
  nand _36276_ (_04896_, _24293_, _04862_);
  and _36277_ (_04897_, _04896_, _22762_);
  and _36278_ (_23032_, _04897_, _04895_);
  and _36279_ (_04898_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  and _36280_ (_04900_, _04748_, _23747_);
  or _36281_ (_23037_, _04900_, _04898_);
  and _36282_ (_04901_, _04656_, _23747_);
  and _36283_ (_04903_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or _36284_ (_23119_, _04903_, _04901_);
  and _36285_ (_04905_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  and _36286_ (_04907_, _04748_, _23946_);
  or _36287_ (_27031_, _04907_, _04905_);
  and _36288_ (_04908_, _04656_, _23824_);
  and _36289_ (_04909_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or _36290_ (_23125_, _04909_, _04908_);
  and _36291_ (_04911_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  and _36292_ (_04913_, _04748_, _23649_);
  or _36293_ (_23136_, _04913_, _04911_);
  and _36294_ (_04914_, _25142_, _24050_);
  and _36295_ (_04915_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  or _36296_ (_23162_, _04915_, _04914_);
  and _36297_ (_04917_, _01809_, _23911_);
  and _36298_ (_04918_, _04917_, _23707_);
  not _36299_ (_04919_, _04917_);
  and _36300_ (_04920_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or _36301_ (_23176_, _04920_, _04918_);
  and _36302_ (_04922_, _23991_, _23754_);
  and _36303_ (_04924_, _04922_, _23898_);
  not _36304_ (_04925_, _04922_);
  and _36305_ (_04926_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  or _36306_ (_23189_, _04926_, _04924_);
  and _36307_ (_04927_, _03300_, _23898_);
  and _36308_ (_04928_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or _36309_ (_23207_, _04928_, _04927_);
  and _36310_ (_04929_, _04832_, _23747_);
  and _36311_ (_04931_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or _36312_ (_23210_, _04931_, _04929_);
  and _36313_ (_04934_, _04832_, _23824_);
  and _36314_ (_04935_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or _36315_ (_26942_, _04935_, _04934_);
  and _36316_ (_04936_, _04797_, _23946_);
  and _36317_ (_04937_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or _36318_ (_23234_, _04937_, _04936_);
  and _36319_ (_04938_, _26589_, _24597_);
  or _36320_ (_04939_, _04938_, _24586_);
  or _36321_ (_04940_, _04939_, _04242_);
  or _36322_ (_04941_, _04940_, _03330_);
  and _36323_ (_04942_, _24546_, _24445_);
  or _36324_ (_04943_, _04942_, _24594_);
  or _36325_ (_04944_, _04943_, _24591_);
  and _36326_ (_04945_, _26582_, _24546_);
  and _36327_ (_04946_, _03275_, _24612_);
  or _36328_ (_04947_, _04946_, _04945_);
  or _36329_ (_04948_, _04947_, _04944_);
  or _36330_ (_04949_, _04948_, _04941_);
  and _36331_ (_04950_, _24613_, _24589_);
  and _36332_ (_04952_, _26650_, _24556_);
  and _36333_ (_04953_, _24598_, _24538_);
  and _36334_ (_04955_, _04953_, _25667_);
  or _36335_ (_04956_, _04955_, _04952_);
  or _36336_ (_04957_, _04956_, _04950_);
  and _36337_ (_04958_, _24593_, _26582_);
  and _36338_ (_04959_, _04958_, _24471_);
  or _36339_ (_04961_, _04959_, _24542_);
  and _36340_ (_04962_, _24592_, _24448_);
  and _36341_ (_04964_, _24556_, _24540_);
  or _36342_ (_04965_, _04964_, _04962_);
  or _36343_ (_04966_, _04965_, _04961_);
  or _36344_ (_04967_, _04966_, _04957_);
  or _36345_ (_04968_, _04967_, _04949_);
  or _36346_ (_04969_, _26583_, _25639_);
  and _36347_ (_04970_, _04953_, _24556_);
  or _36348_ (_04972_, _04970_, _24558_);
  or _36349_ (_04973_, _24618_, _24616_);
  and _36350_ (_04974_, _04973_, _24556_);
  or _36351_ (_04976_, _04974_, _04972_);
  or _36352_ (_04977_, _04976_, _04969_);
  and _36353_ (_04978_, _26589_, _24588_);
  and _36354_ (_04979_, _24593_, _24445_);
  or _36355_ (_04980_, _04979_, _04978_);
  and _36356_ (_04981_, _24545_, _24448_);
  and _36357_ (_04982_, _24589_, _26582_);
  or _36358_ (_04983_, _04982_, _04981_);
  and _36359_ (_04984_, _00234_, _26582_);
  or _36360_ (_04985_, _04984_, _24559_);
  or _36361_ (_04987_, _04985_, _04983_);
  or _36362_ (_04989_, _04987_, _04980_);
  or _36363_ (_04991_, _04989_, _04977_);
  or _36364_ (_04992_, _04991_, _04968_);
  and _36365_ (_04993_, _04992_, _22768_);
  and _36366_ (_04994_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _36367_ (_04995_, _25638_);
  nor _36368_ (_04996_, _24567_, _24447_);
  nor _36369_ (_04998_, _04996_, _04995_);
  nor _36370_ (_05000_, _04998_, _04981_);
  not _36371_ (_05001_, _05000_);
  and _36372_ (_05003_, _05001_, _25662_);
  or _36373_ (_05005_, _05003_, _24572_);
  or _36374_ (_05006_, _05005_, _04994_);
  or _36375_ (_05007_, _05006_, _04993_);
  and _36376_ (_26869_[0], _05007_, _22762_);
  and _36377_ (_05008_, _25078_, _23754_);
  and _36378_ (_05009_, _05008_, _23946_);
  not _36379_ (_05011_, _05008_);
  and _36380_ (_05012_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or _36381_ (_23248_, _05012_, _05009_);
  and _36382_ (_05013_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  and _36383_ (_05014_, _01967_, _23707_);
  or _36384_ (_23255_, _05014_, _05013_);
  or _36385_ (_05016_, _04980_, _04962_);
  or _36386_ (_05017_, _26654_, _26620_);
  and _36387_ (_05018_, _05017_, _24408_);
  or _36388_ (_05019_, _05018_, _05016_);
  or _36389_ (_05020_, _05019_, _04948_);
  or _36390_ (_05022_, _24559_, _24548_);
  or _36391_ (_05023_, _03312_, _26629_);
  or _36392_ (_05024_, _05023_, _05022_);
  and _36393_ (_05025_, _04953_, _24581_);
  or _36394_ (_05026_, _02268_, _26661_);
  or _36395_ (_05027_, _05026_, _05025_);
  and _36396_ (_05028_, _26589_, _24598_);
  or _36397_ (_05029_, _05028_, _24586_);
  or _36398_ (_05030_, _05029_, _24542_);
  or _36399_ (_05031_, _05030_, _05027_);
  or _36400_ (_05032_, _05031_, _05024_);
  or _36401_ (_05033_, _05032_, _05020_);
  or _36402_ (_05034_, _05033_, _04977_);
  and _36403_ (_05035_, _05034_, _22768_);
  and _36404_ (_05036_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _36405_ (_05037_, _05036_, _05005_);
  or _36406_ (_05038_, _05037_, _05035_);
  and _36407_ (_26869_[1], _05038_, _22762_);
  and _36408_ (_05039_, _04832_, _23946_);
  and _36409_ (_05041_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or _36410_ (_23297_, _05041_, _05039_);
  and _36411_ (_05042_, _01809_, _23991_);
  and _36412_ (_05044_, _05042_, _23778_);
  not _36413_ (_05045_, _05042_);
  and _36414_ (_05047_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or _36415_ (_23300_, _05047_, _05044_);
  and _36416_ (_05049_, _24639_, _23649_);
  and _36417_ (_05050_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or _36418_ (_23319_, _05050_, _05049_);
  and _36419_ (_05052_, _02326_, _23707_);
  and _36420_ (_05053_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or _36421_ (_23328_, _05053_, _05052_);
  and _36422_ (_05054_, _25618_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _36423_ (_05055_, _26645_, _24618_);
  and _36424_ (_05057_, _05055_, _24448_);
  or _36425_ (_05058_, _05057_, _04945_);
  or _36426_ (_05060_, _05058_, _02381_);
  or _36427_ (_05061_, _24616_, _24584_);
  and _36428_ (_05063_, _05061_, _26589_);
  or _36429_ (_05064_, _05063_, _24537_);
  or _36430_ (_05065_, _05064_, _26581_);
  or _36431_ (_05066_, _05065_, _05060_);
  or _36432_ (_05067_, _04942_, _03274_);
  or _36433_ (_05068_, _05067_, _04984_);
  and _36434_ (_05070_, _24606_, _24448_);
  and _36435_ (_05072_, _00234_, _24445_);
  or _36436_ (_05073_, _05072_, _05070_);
  or _36437_ (_05074_, _03317_, _02380_);
  and _36438_ (_05075_, _24596_, _24584_);
  and _36439_ (_05077_, _24616_, _26587_);
  or _36440_ (_05079_, _05077_, _05075_);
  and _36441_ (_05080_, _26587_, _24545_);
  and _36442_ (_05081_, _24594_, _24538_);
  or _36443_ (_05083_, _05081_, _05080_);
  or _36444_ (_05085_, _05083_, _05079_);
  or _36445_ (_05086_, _05085_, _05074_);
  and _36446_ (_05087_, _24618_, _24556_);
  and _36447_ (_05088_, _26645_, _26582_);
  or _36448_ (_05089_, _05088_, _05087_);
  and _36449_ (_05090_, _00234_, _24448_);
  or _36450_ (_05091_, _05090_, _26668_);
  or _36451_ (_05093_, _05091_, _05089_);
  or _36452_ (_05095_, _05093_, _05086_);
  or _36453_ (_05096_, _05095_, _05073_);
  or _36454_ (_05097_, _05096_, _05068_);
  or _36455_ (_05098_, _05097_, _05066_);
  and _36456_ (_05099_, _05098_, _25644_);
  or _36457_ (_26870_[0], _05099_, _05054_);
  and _36458_ (_05100_, _05008_, _23824_);
  and _36459_ (_05101_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or _36460_ (_27060_, _05101_, _05100_);
  and _36461_ (_05102_, _01808_, _01758_);
  and _36462_ (_05104_, _05102_, _23707_);
  not _36463_ (_05105_, _05102_);
  and _36464_ (_05107_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or _36465_ (_23388_, _05107_, _05104_);
  and _36466_ (_05109_, _05102_, _24050_);
  and _36467_ (_05110_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _36468_ (_27302_, _05110_, _05109_);
  and _36469_ (_05111_, _05102_, _23946_);
  and _36470_ (_05113_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or _36471_ (_23406_, _05113_, _05111_);
  and _36472_ (_05114_, _24356_, _23656_);
  and _36473_ (_05116_, _05114_, _23898_);
  not _36474_ (_05117_, _05114_);
  and _36475_ (_05118_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or _36476_ (_23410_, _05118_, _05116_);
  and _36477_ (_05119_, _24370_, _24005_);
  and _36478_ (_05120_, _05119_, _23946_);
  not _36479_ (_05121_, _05119_);
  and _36480_ (_05122_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  or _36481_ (_23426_, _05122_, _05120_);
  and _36482_ (_05125_, _24282_, _23754_);
  and _36483_ (_05126_, _05125_, _24050_);
  not _36484_ (_05127_, _05125_);
  and _36485_ (_05128_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  or _36486_ (_23477_, _05128_, _05126_);
  and _36487_ (_05129_, _05008_, _23778_);
  and _36488_ (_05130_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or _36489_ (_23504_, _05130_, _05129_);
  and _36490_ (_05131_, _05102_, _23778_);
  and _36491_ (_05132_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or _36492_ (_23507_, _05132_, _05131_);
  and _36493_ (_05133_, _05102_, _23898_);
  and _36494_ (_05134_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or _36495_ (_23513_, _05134_, _05133_);
  and _36496_ (_05135_, _05125_, _23707_);
  and _36497_ (_05137_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  or _36498_ (_23517_, _05137_, _05135_);
  and _36499_ (_05138_, _24852_, _23898_);
  and _36500_ (_05139_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  or _36501_ (_23554_, _05139_, _05138_);
  and _36502_ (_05140_, _05102_, _23747_);
  and _36503_ (_05141_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or _36504_ (_23566_, _05141_, _05140_);
  nand _36505_ (_05142_, _24299_, _23702_);
  not _36506_ (_05143_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _36507_ (_05144_, _04864_, _24313_);
  nor _36508_ (_05145_, _05144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _36509_ (_05146_, _05145_, _05143_);
  and _36510_ (_05147_, _05145_, _05143_);
  or _36511_ (_05148_, _05147_, _05146_);
  and _36512_ (_05149_, _05148_, _04861_);
  and _36513_ (_05151_, _04876_, _24310_);
  and _36514_ (_05152_, _05151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _36515_ (_05153_, _05152_, _05143_);
  and _36516_ (_05154_, _05152_, _05143_);
  or _36517_ (_05156_, _05154_, _05153_);
  and _36518_ (_05157_, _05156_, _24302_);
  and _36519_ (_05158_, _24309_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _36520_ (_05159_, _05158_, _26114_);
  and _36521_ (_05160_, _05159_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _36522_ (_05161_, _05160_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _36523_ (_05162_, _05161_, _26110_);
  or _36524_ (_05163_, _05162_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _36525_ (_05164_, _05158_, _26115_);
  and _36526_ (_05165_, _05164_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _36527_ (_05166_, _05165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _36528_ (_05167_, _05166_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _36529_ (_05168_, _05167_, _26097_);
  and _36530_ (_05169_, _05168_, _05163_);
  or _36531_ (_05170_, _05169_, _05157_);
  or _36532_ (_05171_, _05170_, _05149_);
  or _36533_ (_05172_, _05171_, _24299_);
  and _36534_ (_05173_, _05172_, _24294_);
  and _36535_ (_05174_, _05173_, _05142_);
  and _36536_ (_05175_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _36537_ (_05176_, _05175_, _05174_);
  and _36538_ (_23573_, _05176_, _22762_);
  and _36539_ (_05177_, _05125_, _23649_);
  and _36540_ (_05178_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  or _36541_ (_23586_, _05178_, _05177_);
  and _36542_ (_05180_, _01809_, _23903_);
  and _36543_ (_05181_, _05180_, _23649_);
  not _36544_ (_05182_, _05180_);
  and _36545_ (_05183_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or _36546_ (_23620_, _05183_, _05181_);
  and _36547_ (_05184_, _05114_, _23707_);
  and _36548_ (_05186_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or _36549_ (_23650_, _05186_, _05184_);
  and _36550_ (_05187_, _25078_, _24356_);
  and _36551_ (_05188_, _05187_, _23824_);
  not _36552_ (_05189_, _05187_);
  and _36553_ (_05190_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or _36554_ (_23659_, _05190_, _05188_);
  and _36555_ (_05191_, _25142_, _23824_);
  and _36556_ (_05192_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  or _36557_ (_23685_, _05192_, _05191_);
  and _36558_ (_05193_, _24201_, _23911_);
  not _36559_ (_05194_, _05193_);
  and _36560_ (_05195_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  and _36561_ (_05197_, _05193_, _23707_);
  or _36562_ (_23698_, _05197_, _05195_);
  and _36563_ (_05199_, _24282_, _24201_);
  not _36564_ (_05200_, _05199_);
  and _36565_ (_05201_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  and _36566_ (_05203_, _05199_, _23898_);
  or _36567_ (_23703_, _05203_, _05201_);
  and _36568_ (_05204_, _02321_, _23778_);
  and _36569_ (_05205_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  or _36570_ (_23723_, _05205_, _05204_);
  nor _36571_ (_26912_, _02387_, rst);
  and _36572_ (_05206_, _24063_, _23073_);
  and _36573_ (_05207_, _05206_, _25171_);
  and _36574_ (_05208_, _05207_, _25926_);
  nand _36575_ (_05209_, _05208_, _23702_);
  or _36576_ (_05210_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _36577_ (_05211_, _05210_, _22762_);
  and _36578_ (_26874_[7], _05211_, _05209_);
  and _36579_ (_05212_, _05206_, _26683_);
  not _36580_ (_05213_, _05212_);
  nor _36581_ (_05214_, _05213_, _23702_);
  not _36582_ (_05215_, _25926_);
  and _36583_ (_05216_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _36584_ (_05217_, _05216_, _05215_);
  or _36585_ (_05218_, _05217_, _05214_);
  or _36586_ (_05219_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _36587_ (_05221_, _05219_, _22762_);
  and _36588_ (_26875_[7], _05221_, _05218_);
  and _36589_ (_05222_, _05206_, _02310_);
  and _36590_ (_05223_, _05222_, _25926_);
  nand _36591_ (_05224_, _05223_, _23702_);
  or _36592_ (_05226_, _05223_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _36593_ (_05227_, _05226_, _22762_);
  and _36594_ (_26876_[7], _05227_, _05224_);
  and _36595_ (_05228_, _05206_, _24076_);
  and _36596_ (_05229_, _05228_, _25926_);
  not _36597_ (_05230_, _05229_);
  nor _36598_ (_05231_, _05230_, _23702_);
  and _36599_ (_05233_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or _36600_ (_05234_, _05233_, _05231_);
  and _36601_ (_26877_[7], _05234_, _22762_);
  and _36602_ (_05235_, _02311_, _25171_);
  and _36603_ (_05236_, _05235_, _25926_);
  and _36604_ (_05237_, _05236_, _26750_);
  or _36605_ (_05238_, _05222_, _05228_);
  or _36606_ (_05239_, _05235_, _05238_);
  nor _36607_ (_05240_, _05239_, _05212_);
  or _36608_ (_05241_, _05240_, _05215_);
  or _36609_ (_05242_, _05238_, _05212_);
  and _36610_ (_05243_, _05242_, _25926_);
  or _36611_ (_05244_, _05243_, _05241_);
  and _36612_ (_05245_, _05244_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or _36613_ (_05246_, _05245_, _05237_);
  and _36614_ (_26878_[7], _05246_, _22762_);
  and _36615_ (_05247_, _02311_, _26683_);
  nor _36616_ (_05248_, _05247_, _05235_);
  not _36617_ (_05249_, _05248_);
  nor _36618_ (_05250_, _05249_, _05238_);
  or _36619_ (_05251_, _05250_, _05215_);
  or _36620_ (_05252_, _05251_, _05239_);
  and _36621_ (_05253_, _05252_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _36622_ (_05254_, _05247_, _25926_);
  not _36623_ (_05255_, _05254_);
  nor _36624_ (_05256_, _05255_, _23702_);
  or _36625_ (_05257_, _05256_, _05253_);
  and _36626_ (_26879_[7], _05257_, _22762_);
  nor _36627_ (_05259_, _02315_, _23702_);
  and _36628_ (_05260_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or _36629_ (_05261_, _05260_, _05259_);
  and _36630_ (_26880_[7], _05261_, _22762_);
  and _36631_ (_05262_, _02311_, _24076_);
  and _36632_ (_05263_, _05262_, _25926_);
  and _36633_ (_05264_, _05263_, _26750_);
  nor _36634_ (_05265_, _05262_, _02312_);
  and _36635_ (_05266_, _05265_, _05248_);
  or _36636_ (_05267_, _05266_, _05215_);
  not _36637_ (_05268_, _02312_);
  nand _36638_ (_05269_, _05248_, _05268_);
  and _36639_ (_05270_, _05269_, _25926_);
  or _36640_ (_05271_, _05270_, _05267_);
  and _36641_ (_05272_, _05271_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or _36642_ (_05273_, _05272_, _05264_);
  and _36643_ (_26881_[7], _05273_, _22762_);
  or _36644_ (_05275_, _05223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  not _36645_ (_05276_, _05223_);
  or _36646_ (_05277_, _05276_, _23816_);
  and _36647_ (_23763_, _05277_, _05275_);
  and _36648_ (_05278_, _05223_, _23898_);
  and _36649_ (_05279_, _05276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or _36650_ (_23815_, _05279_, _05278_);
  and _36651_ (_05281_, _23986_, _23754_);
  and _36652_ (_05282_, _05281_, _23747_);
  not _36653_ (_05283_, _05281_);
  and _36654_ (_05284_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or _36655_ (_23819_, _05284_, _05282_);
  and _36656_ (_05285_, _05223_, _23778_);
  and _36657_ (_05286_, _05276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or _36658_ (_23826_, _05286_, _05285_);
  and _36659_ (_05288_, _23911_, _23754_);
  and _36660_ (_05289_, _05288_, _23649_);
  not _36661_ (_05290_, _05288_);
  and _36662_ (_05291_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  or _36663_ (_23891_, _05291_, _05289_);
  and _36664_ (_05292_, _05223_, _23946_);
  and _36665_ (_05293_, _05276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or _36666_ (_27278_, _05293_, _05292_);
  and _36667_ (_05294_, _05223_, _23649_);
  and _36668_ (_05295_, _05276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or _36669_ (_23928_, _05295_, _05294_);
  and _36670_ (_05296_, _05223_, _23747_);
  and _36671_ (_05297_, _05276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or _36672_ (_23931_, _05297_, _05296_);
  and _36673_ (_05298_, _01758_, _23752_);
  and _36674_ (_05299_, _05298_, _23824_);
  not _36675_ (_05301_, _05298_);
  and _36676_ (_05302_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or _36677_ (_23996_, _05302_, _05299_);
  and _36678_ (_05303_, _05298_, _23649_);
  and _36679_ (_05304_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or _36680_ (_23999_, _05304_, _05303_);
  and _36681_ (_05305_, _05298_, _23747_);
  and _36682_ (_05307_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or _36683_ (_24002_, _05307_, _05305_);
  nor _36684_ (_26897_[5], _00727_, rst);
  and _36685_ (_05308_, _05288_, _23898_);
  and _36686_ (_05309_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  or _36687_ (_24091_, _05309_, _05308_);
  and _36688_ (_05310_, _05298_, _23707_);
  and _36689_ (_05311_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or _36690_ (_24097_, _05311_, _05310_);
  and _36691_ (_05313_, _05298_, _24050_);
  and _36692_ (_05314_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _36693_ (_24099_, _05314_, _05313_);
  and _36694_ (_05315_, _05288_, _23707_);
  and _36695_ (_05316_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or _36696_ (_24106_, _05316_, _05315_);
  and _36697_ (_05317_, _05288_, _24050_);
  and _36698_ (_05318_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  or _36699_ (_27057_, _05318_, _05317_);
  and _36700_ (_05319_, _01758_, _23656_);
  and _36701_ (_05320_, _05319_, _23747_);
  not _36702_ (_05322_, _05319_);
  and _36703_ (_05323_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _36704_ (_24133_, _05323_, _05320_);
  and _36705_ (_05324_, _05319_, _23946_);
  and _36706_ (_05325_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _36707_ (_27234_, _05325_, _05324_);
  and _36708_ (_05326_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  and _36709_ (_05327_, _05199_, _23778_);
  or _36710_ (_27230_, _05327_, _05326_);
  and _36711_ (_05328_, _05319_, _23649_);
  and _36712_ (_05329_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or _36713_ (_24183_, _05329_, _05328_);
  and _36714_ (_05330_, _05125_, _23778_);
  and _36715_ (_05331_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  or _36716_ (_24200_, _05331_, _05330_);
  and _36717_ (_05332_, _05319_, _23707_);
  and _36718_ (_05333_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _36719_ (_24202_, _05333_, _05332_);
  and _36720_ (_05334_, _05298_, _23778_);
  and _36721_ (_05335_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or _36722_ (_24205_, _05335_, _05334_);
  and _36723_ (_05336_, _23785_, _23662_);
  and _36724_ (_05337_, _05336_, _24085_);
  not _36725_ (_05338_, _05337_);
  and _36726_ (_05339_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  and _36727_ (_05340_, _05337_, _23649_);
  or _36728_ (_24227_, _05340_, _05339_);
  and _36729_ (_05342_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  and _36730_ (_05343_, _05337_, _23747_);
  or _36731_ (_24233_, _05343_, _05342_);
  and _36732_ (_05344_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  and _36733_ (_05345_, _05337_, _23824_);
  or _36734_ (_24278_, _05345_, _05344_);
  and _36735_ (_05346_, _01758_, _25078_);
  and _36736_ (_05347_, _05346_, _24050_);
  not _36737_ (_05348_, _05346_);
  and _36738_ (_05349_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or _36739_ (_24281_, _05349_, _05347_);
  and _36740_ (_05350_, _01808_, _23754_);
  and _36741_ (_05351_, _05350_, _23707_);
  not _36742_ (_05352_, _05350_);
  and _36743_ (_05353_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  or _36744_ (_24298_, _05353_, _05351_);
  and _36745_ (_05354_, _05336_, _24010_);
  not _36746_ (_05355_, _05354_);
  and _36747_ (_05356_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  and _36748_ (_05357_, _05354_, _23778_);
  or _36749_ (_24306_, _05357_, _05356_);
  and _36750_ (_05358_, _05336_, _24275_);
  not _36751_ (_05359_, _05358_);
  and _36752_ (_05360_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  and _36753_ (_05361_, _05358_, _23898_);
  or _36754_ (_27105_, _05361_, _05360_);
  and _36755_ (_05362_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  and _36756_ (_05363_, _05358_, _24050_);
  or _36757_ (_24311_, _05363_, _05362_);
  and _36758_ (_05364_, _05319_, _23898_);
  and _36759_ (_05365_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _36760_ (_24314_, _05365_, _05364_);
  and _36761_ (_05366_, _05319_, _23778_);
  and _36762_ (_05367_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _36763_ (_24321_, _05367_, _05366_);
  and _36764_ (_05368_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  and _36765_ (_05369_, _05358_, _23707_);
  or _36766_ (_24327_, _05369_, _05368_);
  and _36767_ (_05371_, _01809_, _23784_);
  and _36768_ (_05372_, _05371_, _23778_);
  not _36769_ (_05373_, _05371_);
  and _36770_ (_05374_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or _36771_ (_24330_, _05374_, _05372_);
  and _36772_ (_05375_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  and _36773_ (_05376_, _05337_, _23707_);
  or _36774_ (_24355_, _05376_, _05375_);
  and _36775_ (_05377_, _04797_, _23747_);
  and _36776_ (_05378_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or _36777_ (_24357_, _05378_, _05377_);
  and _36778_ (_05379_, _01758_, _24282_);
  and _36779_ (_05380_, _05379_, _23707_);
  not _36780_ (_05381_, _05379_);
  and _36781_ (_05382_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or _36782_ (_24387_, _05382_, _05380_);
  and _36783_ (_05384_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  and _36784_ (_05385_, _05337_, _24050_);
  or _36785_ (_24390_, _05385_, _05384_);
  and _36786_ (_05387_, _05379_, _24050_);
  and _36787_ (_05388_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _36788_ (_27204_, _05388_, _05387_);
  and _36789_ (_05390_, _05379_, _23946_);
  and _36790_ (_05391_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _36791_ (_24395_, _05391_, _05390_);
  and _36792_ (_05392_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  and _36793_ (_05393_, _05337_, _23946_);
  or _36794_ (_24398_, _05393_, _05392_);
  and _36795_ (_05394_, _05346_, _23747_);
  and _36796_ (_05395_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or _36797_ (_24410_, _05395_, _05394_);
  and _36798_ (_05396_, _05346_, _23824_);
  and _36799_ (_05397_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or _36800_ (_24413_, _05397_, _05396_);
  and _36801_ (_05398_, _05336_, _23784_);
  not _36802_ (_05399_, _05398_);
  and _36803_ (_05400_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and _36804_ (_05401_, _05398_, _23649_);
  or _36805_ (_24416_, _05401_, _05400_);
  and _36806_ (_05402_, _05346_, _23898_);
  and _36807_ (_05403_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or _36808_ (_24419_, _05403_, _05402_);
  and _36809_ (_05404_, _05346_, _23778_);
  and _36810_ (_05405_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or _36811_ (_24423_, _05405_, _05404_);
  and _36812_ (_05407_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and _36813_ (_05409_, _05398_, _23946_);
  or _36814_ (_24433_, _05409_, _05407_);
  and _36815_ (_05410_, _01808_, _23076_);
  and _36816_ (_05411_, _05410_, _23649_);
  not _36817_ (_05412_, _05410_);
  and _36818_ (_05413_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  or _36819_ (_24449_, _05413_, _05411_);
  and _36820_ (_05414_, _05379_, _23778_);
  and _36821_ (_05415_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or _36822_ (_27203_, _05415_, _05414_);
  and _36823_ (_05416_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and _36824_ (_05417_, _05398_, _23707_);
  or _36825_ (_24465_, _05417_, _05416_);
  and _36826_ (_05419_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  and _36827_ (_05420_, _05337_, _23778_);
  or _36828_ (_24468_, _05420_, _05419_);
  and _36829_ (_05422_, _05379_, _23747_);
  and _36830_ (_05424_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _36831_ (_24496_, _05424_, _05422_);
  and _36832_ (_05425_, _05379_, _23824_);
  and _36833_ (_05426_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _36834_ (_24499_, _05426_, _05425_);
  and _36835_ (_05427_, _05379_, _23898_);
  and _36836_ (_05428_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or _36837_ (_24502_, _05428_, _05427_);
  and _36838_ (_05429_, _01758_, _23911_);
  and _36839_ (_05430_, _05429_, _23824_);
  not _36840_ (_05431_, _05429_);
  and _36841_ (_05432_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or _36842_ (_24547_, _05432_, _05430_);
  and _36843_ (_05433_, _05429_, _23649_);
  and _36844_ (_05434_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or _36845_ (_24551_, _05434_, _05433_);
  and _36846_ (_05435_, _05429_, _23747_);
  and _36847_ (_05436_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or _36848_ (_24557_, _05436_, _05435_);
  and _36849_ (_05437_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  and _36850_ (_05438_, _05358_, _23946_);
  or _36851_ (_24571_, _05438_, _05437_);
  and _36852_ (_05439_, _05371_, _23898_);
  and _36853_ (_05440_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or _36854_ (_24580_, _05440_, _05439_);
  and _36855_ (_05441_, _05371_, _23747_);
  and _36856_ (_05442_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or _36857_ (_24583_, _05442_, _05441_);
  and _36858_ (_05443_, _05429_, _24050_);
  and _36859_ (_05444_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or _36860_ (_24590_, _05444_, _05443_);
  and _36861_ (_05445_, _01809_, _24085_);
  and _36862_ (_05446_, _05445_, _23778_);
  not _36863_ (_05447_, _05445_);
  and _36864_ (_05448_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  or _36865_ (_27106_, _05448_, _05446_);
  and _36866_ (_05449_, _05371_, _24050_);
  and _36867_ (_05450_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or _36868_ (_24603_, _05450_, _05449_);
  and _36869_ (_05452_, _05371_, _23707_);
  and _36870_ (_05453_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or _36871_ (_24609_, _05453_, _05452_);
  and _36872_ (_05454_, _01758_, _24010_);
  and _36873_ (_05455_, _05454_, _24050_);
  not _36874_ (_05457_, _05454_);
  and _36875_ (_05458_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or _36876_ (_24638_, _05458_, _05455_);
  not _36877_ (_05459_, _05208_);
  and _36878_ (_05460_, _05459_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _36879_ (_05461_, _05208_, _24685_);
  or _36880_ (_05462_, _05461_, _05460_);
  and _36881_ (_26874_[0], _05462_, _22762_);
  or _36882_ (_05463_, _05459_, _23892_);
  or _36883_ (_05464_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _36884_ (_05466_, _05464_, _22762_);
  and _36885_ (_26874_[1], _05466_, _05463_);
  or _36886_ (_05467_, _05459_, _23816_);
  or _36887_ (_05468_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _36888_ (_05469_, _05468_, _22762_);
  and _36889_ (_26874_[2], _05469_, _05467_);
  or _36890_ (_05470_, _05459_, _23738_);
  or _36891_ (_05471_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _36892_ (_05472_, _05471_, _22762_);
  and _36893_ (_26874_[3], _05472_, _05470_);
  or _36894_ (_05474_, _05459_, _23642_);
  or _36895_ (_05475_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _36896_ (_05477_, _05475_, _22762_);
  and _36897_ (_26874_[4], _05477_, _05474_);
  or _36898_ (_05478_, _05459_, _23939_);
  or _36899_ (_05480_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _36900_ (_05481_, _05480_, _22762_);
  and _36901_ (_26874_[5], _05481_, _05478_);
  or _36902_ (_05482_, _05459_, _24043_);
  or _36903_ (_05483_, _05208_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _36904_ (_05484_, _05483_, _22762_);
  and _36905_ (_26874_[6], _05484_, _05482_);
  nor _36906_ (_05485_, _05215_, _23772_);
  and _36907_ (_05486_, _05485_, _05212_);
  nand _36908_ (_05487_, _05212_, _25926_);
  and _36909_ (_05488_, _05487_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or _36910_ (_05489_, _05488_, _05486_);
  and _36911_ (_26875_[0], _05489_, _22762_);
  and _36912_ (_05490_, _05212_, _23892_);
  and _36913_ (_05491_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or _36914_ (_05492_, _05491_, _05215_);
  or _36915_ (_05493_, _05492_, _05490_);
  or _36916_ (_05494_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _36917_ (_05495_, _05494_, _22762_);
  and _36918_ (_26875_[1], _05495_, _05493_);
  and _36919_ (_05496_, _05212_, _23816_);
  and _36920_ (_05497_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _36921_ (_05499_, _05497_, _05215_);
  or _36922_ (_05500_, _05499_, _05496_);
  or _36923_ (_05501_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _36924_ (_05502_, _05501_, _22762_);
  and _36925_ (_26875_[2], _05502_, _05500_);
  and _36926_ (_05504_, _05212_, _23738_);
  and _36927_ (_05505_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _36928_ (_05506_, _05505_, _05215_);
  or _36929_ (_05507_, _05506_, _05504_);
  or _36930_ (_05508_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _36931_ (_05509_, _05508_, _22762_);
  and _36932_ (_26875_[3], _05509_, _05507_);
  and _36933_ (_05510_, _05212_, _23642_);
  and _36934_ (_05511_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _36935_ (_05512_, _05511_, _05215_);
  or _36936_ (_05513_, _05512_, _05510_);
  or _36937_ (_05514_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _36938_ (_05515_, _05514_, _22762_);
  and _36939_ (_26875_[4], _05515_, _05513_);
  and _36940_ (_05516_, _05212_, _23939_);
  and _36941_ (_05517_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _36942_ (_05518_, _05517_, _05215_);
  or _36943_ (_05519_, _05518_, _05516_);
  or _36944_ (_05520_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _36945_ (_05521_, _05520_, _22762_);
  and _36946_ (_26875_[5], _05521_, _05519_);
  and _36947_ (_05522_, _05212_, _24043_);
  and _36948_ (_05523_, _05213_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _36949_ (_05524_, _05523_, _05215_);
  or _36950_ (_05525_, _05524_, _05522_);
  or _36951_ (_05526_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _36952_ (_05527_, _05526_, _22762_);
  and _36953_ (_26875_[6], _05527_, _05525_);
  not _36954_ (_05528_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _36955_ (_05529_, _05212_, _05207_);
  not _36956_ (_05530_, _05222_);
  and _36957_ (_05531_, _05530_, _05529_);
  nor _36958_ (_05532_, _05531_, _05215_);
  nor _36959_ (_05533_, _05532_, _05528_);
  nand _36960_ (_05534_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _36961_ (_05535_, _05534_, _05529_);
  and _36962_ (_05536_, _05223_, _24685_);
  or _36963_ (_05537_, _05536_, _05535_);
  or _36964_ (_05538_, _05537_, _05533_);
  and _36965_ (_26876_[0], _05538_, _22762_);
  and _36966_ (_05539_, _05223_, _23892_);
  and _36967_ (_05540_, _05276_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or _36968_ (_05541_, _05540_, _05539_);
  and _36969_ (_26876_[1], _05541_, _22762_);
  or _36970_ (_05544_, _05223_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _36971_ (_05545_, _05544_, _22762_);
  and _36972_ (_26876_[2], _05545_, _05277_);
  or _36973_ (_05547_, _05276_, _23738_);
  or _36974_ (_05548_, _05223_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _36975_ (_05550_, _05548_, _22762_);
  and _36976_ (_26876_[3], _05550_, _05547_);
  or _36977_ (_05551_, _05276_, _23642_);
  or _36978_ (_05552_, _05223_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _36979_ (_05553_, _05552_, _22762_);
  and _36980_ (_26876_[4], _05553_, _05551_);
  and _36981_ (_05554_, _05223_, _23939_);
  and _36982_ (_05555_, _05276_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or _36983_ (_05556_, _05555_, _05554_);
  and _36984_ (_26876_[5], _05556_, _22762_);
  and _36985_ (_05558_, _05223_, _24043_);
  and _36986_ (_05559_, _05276_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or _36987_ (_05560_, _05559_, _05558_);
  and _36988_ (_26876_[6], _05560_, _22762_);
  and _36989_ (_05561_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _36990_ (_05562_, _05485_, _05228_);
  or _36991_ (_05563_, _05562_, _05561_);
  and _36992_ (_26877_[0], _05563_, _22762_);
  and _36993_ (_05564_, _05229_, _23892_);
  or _36994_ (_05565_, _05230_, _05532_);
  and _36995_ (_05566_, _05565_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or _36996_ (_05567_, _05566_, _05564_);
  and _36997_ (_26877_[1], _05567_, _22762_);
  and _36998_ (_05569_, _05229_, _23816_);
  and _36999_ (_05571_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or _37000_ (_05572_, _05571_, _05569_);
  and _37001_ (_26877_[2], _05572_, _22762_);
  and _37002_ (_05574_, _05229_, _23738_);
  and _37003_ (_05575_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or _37004_ (_05576_, _05575_, _05574_);
  and _37005_ (_26877_[3], _05576_, _22762_);
  and _37006_ (_05578_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _37007_ (_05579_, _05229_, _23642_);
  or _37008_ (_05580_, _05579_, _05578_);
  and _37009_ (_26877_[4], _05580_, _22762_);
  and _37010_ (_05581_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and _37011_ (_05582_, _05229_, _23939_);
  or _37012_ (_05583_, _05582_, _05581_);
  and _37013_ (_26877_[5], _05583_, _22762_);
  and _37014_ (_05585_, _05229_, _24043_);
  and _37015_ (_05586_, _05230_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or _37016_ (_05588_, _05586_, _05585_);
  and _37017_ (_26877_[6], _05588_, _22762_);
  and _37018_ (_05590_, _05454_, _23946_);
  and _37019_ (_05591_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or _37020_ (_27172_, _05591_, _05590_);
  or _37021_ (_05592_, _05242_, _05241_);
  and _37022_ (_05593_, _05592_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _37023_ (_05594_, _05485_, _05235_);
  or _37024_ (_05595_, _05594_, _05593_);
  and _37025_ (_26878_[0], _05595_, _22762_);
  and _37026_ (_05596_, _05236_, _23892_);
  and _37027_ (_05597_, _05244_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  or _37028_ (_05599_, _05597_, _05596_);
  and _37029_ (_26878_[1], _05599_, _22762_);
  and _37030_ (_05600_, _05236_, _23816_);
  and _37031_ (_05601_, _05244_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or _37032_ (_05602_, _05601_, _05600_);
  and _37033_ (_26878_[2], _05602_, _22762_);
  and _37034_ (_05603_, _05236_, _23738_);
  and _37035_ (_05604_, _05244_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or _37036_ (_05605_, _05604_, _05603_);
  and _37037_ (_26878_[3], _05605_, _22762_);
  and _37038_ (_05606_, _05592_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _37039_ (_05607_, _05236_, _23642_);
  or _37040_ (_05608_, _05607_, _05606_);
  and _37041_ (_26878_[4], _05608_, _22762_);
  and _37042_ (_05609_, _05236_, _23939_);
  and _37043_ (_05610_, _05244_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or _37044_ (_05611_, _05610_, _05609_);
  and _37045_ (_26878_[5], _05611_, _22762_);
  and _37046_ (_05612_, _05236_, _24043_);
  and _37047_ (_05613_, _05244_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  or _37048_ (_05614_, _05613_, _05612_);
  and _37049_ (_26878_[6], _05614_, _22762_);
  and _37050_ (_05615_, _05252_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _37051_ (_05616_, _05485_, _05247_);
  or _37052_ (_05617_, _05616_, _05615_);
  and _37053_ (_26879_[0], _05617_, _22762_);
  and _37054_ (_05618_, _05251_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _37055_ (_05619_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _37056_ (_05620_, _05619_, _05239_);
  and _37057_ (_05621_, _05254_, _23892_);
  or _37058_ (_05623_, _05621_, _05620_);
  or _37059_ (_05624_, _05623_, _05618_);
  and _37060_ (_26879_[1], _05624_, _22762_);
  and _37061_ (_05626_, _05254_, _23816_);
  and _37062_ (_05627_, _05255_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  or _37063_ (_05628_, _05627_, _05626_);
  and _37064_ (_26879_[2], _05628_, _22762_);
  and _37065_ (_05629_, _05254_, _23738_);
  and _37066_ (_05630_, _05251_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and _37067_ (_05631_, _25926_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and _37068_ (_05632_, _05631_, _05239_);
  or _37069_ (_05634_, _05632_, _05630_);
  or _37070_ (_05635_, _05634_, _05629_);
  and _37071_ (_26879_[3], _05635_, _22762_);
  and _37072_ (_05636_, _05254_, _23642_);
  and _37073_ (_05637_, _05252_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  or _37074_ (_05638_, _05637_, _05636_);
  and _37075_ (_26879_[4], _05638_, _22762_);
  and _37076_ (_05640_, _05255_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _37077_ (_05641_, _05254_, _23939_);
  or _37078_ (_05642_, _05641_, _05640_);
  and _37079_ (_26879_[5], _05642_, _22762_);
  and _37080_ (_05644_, _05254_, _24043_);
  and _37081_ (_05645_, _05252_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or _37082_ (_05646_, _05645_, _05644_);
  and _37083_ (_26879_[6], _05646_, _22762_);
  and _37084_ (_05647_, _05454_, _23649_);
  and _37085_ (_05648_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or _37086_ (_24681_, _05648_, _05647_);
  and _37087_ (_05649_, _05485_, _02312_);
  and _37088_ (_05650_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  or _37089_ (_05651_, _05650_, _05649_);
  and _37090_ (_26880_[0], _05651_, _22762_);
  and _37091_ (_05652_, _02313_, _23892_);
  and _37092_ (_05653_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  or _37093_ (_05654_, _05653_, _05652_);
  and _37094_ (_26880_[1], _05654_, _22762_);
  and _37095_ (_05655_, _02313_, _23816_);
  and _37096_ (_05656_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or _37097_ (_05657_, _05656_, _05655_);
  and _37098_ (_26880_[2], _05657_, _22762_);
  and _37099_ (_05658_, _02313_, _23738_);
  and _37100_ (_05660_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or _37101_ (_05662_, _05660_, _05658_);
  and _37102_ (_26880_[3], _05662_, _22762_);
  and _37103_ (_05663_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _37104_ (_05664_, _02313_, _23642_);
  or _37105_ (_05665_, _05664_, _05663_);
  and _37106_ (_26880_[4], _05665_, _22762_);
  and _37107_ (_05666_, _02313_, _23939_);
  and _37108_ (_05667_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or _37109_ (_05668_, _05667_, _05666_);
  and _37110_ (_26880_[5], _05668_, _22762_);
  and _37111_ (_05669_, _02315_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or _37112_ (_05670_, _05669_, _02314_);
  and _37113_ (_26880_[6], _05670_, _22762_);
  and _37114_ (_05671_, _05485_, _05262_);
  and _37115_ (_05672_, _05271_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or _37116_ (_05674_, _05672_, _05671_);
  and _37117_ (_26881_[0], _05674_, _22762_);
  and _37118_ (_05675_, _05263_, _23892_);
  and _37119_ (_05676_, _05271_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  or _37120_ (_05677_, _05676_, _05675_);
  and _37121_ (_26881_[1], _05677_, _22762_);
  and _37122_ (_05679_, _05263_, _23816_);
  or _37123_ (_05680_, _05267_, _05269_);
  and _37124_ (_05681_, _05680_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or _37125_ (_05682_, _05681_, _05679_);
  and _37126_ (_26881_[2], _05682_, _22762_);
  and _37127_ (_05683_, _05263_, _23738_);
  and _37128_ (_05684_, _05271_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  or _37129_ (_05685_, _05684_, _05683_);
  and _37130_ (_26881_[3], _05685_, _22762_);
  and _37131_ (_05686_, _05263_, _23642_);
  and _37132_ (_05687_, _05271_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or _37133_ (_05688_, _05687_, _05686_);
  and _37134_ (_26881_[4], _05688_, _22762_);
  and _37135_ (_05690_, _05680_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _37136_ (_05691_, _05263_, _23939_);
  or _37137_ (_05692_, _05691_, _05690_);
  and _37138_ (_26881_[5], _05692_, _22762_);
  and _37139_ (_05693_, _05263_, _24043_);
  and _37140_ (_05694_, _05271_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or _37141_ (_05695_, _05694_, _05693_);
  and _37142_ (_26881_[6], _05695_, _22762_);
  and _37143_ (_05696_, _05410_, _23747_);
  and _37144_ (_05697_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  or _37145_ (_24697_, _05697_, _05696_);
  and _37146_ (_05698_, _25142_, _23898_);
  and _37147_ (_05699_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  or _37148_ (_27200_, _05699_, _05698_);
  and _37149_ (_05701_, _23991_, _23664_);
  and _37150_ (_05702_, _05701_, _23898_);
  not _37151_ (_05703_, _05701_);
  and _37152_ (_05704_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or _37153_ (_25107_, _05704_, _05702_);
  and _37154_ (_05705_, _05336_, _23911_);
  not _37155_ (_05706_, _05705_);
  and _37156_ (_05708_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and _37157_ (_05709_, _05705_, _23649_);
  or _37158_ (_25124_, _05709_, _05708_);
  and _37159_ (_05710_, _02325_, _23991_);
  and _37160_ (_05711_, _05710_, _23649_);
  not _37161_ (_05712_, _05710_);
  and _37162_ (_05713_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  or _37163_ (_27162_, _05713_, _05711_);
  and _37164_ (_05714_, _02325_, _23903_);
  and _37165_ (_05715_, _05714_, _23946_);
  not _37166_ (_05716_, _05714_);
  and _37167_ (_05717_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  or _37168_ (_25147_, _05717_, _05715_);
  and _37169_ (_05718_, _05701_, _23778_);
  and _37170_ (_05719_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or _37171_ (_25149_, _05719_, _05718_);
  and _37172_ (_05720_, _05714_, _23778_);
  and _37173_ (_05721_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  or _37174_ (_25152_, _05721_, _05720_);
  and _37175_ (_05722_, _04917_, _23946_);
  and _37176_ (_05723_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or _37177_ (_25177_, _05723_, _05722_);
  and _37178_ (_05724_, _04917_, _23747_);
  and _37179_ (_05725_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or _37180_ (_25180_, _05725_, _05724_);
  not _37181_ (_05726_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _37182_ (_05727_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and _37183_ (_05728_, _05727_, _05726_);
  and _37184_ (_05729_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _22762_);
  and _37185_ (_27303_, _05729_, _05728_);
  nor _37186_ (_05730_, _05728_, rst);
  nand _37187_ (_05731_, _05727_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or _37188_ (_05732_, _05727_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _37189_ (_05733_, _05732_, _05731_);
  and _37190_ (_27304_[3], _05733_, _05730_);
  not _37191_ (_05734_, _00014_);
  nor _37192_ (_05735_, _05734_, _26817_);
  and _37193_ (_05736_, _02397_, _26777_);
  and _37194_ (_05737_, _05736_, _00037_);
  and _37195_ (_05738_, _05737_, _05735_);
  not _37196_ (_05739_, _00263_);
  nand _37197_ (_05740_, _00451_, _05739_);
  and _37198_ (_05741_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _37199_ (_05742_, _00267_, _00264_);
  not _37200_ (_05743_, _05742_);
  nor _37201_ (_05744_, _24291_, _23304_);
  nor _37202_ (_05745_, _05744_, _04389_);
  nor _37203_ (_05746_, _05745_, _05743_);
  nor _37204_ (_05747_, _05746_, _05741_);
  nand _37205_ (_05748_, _05747_, _05740_);
  nand _37206_ (_05749_, _05748_, _00257_);
  nor _37207_ (_05750_, _01061_, _00257_);
  not _37208_ (_05751_, _05750_);
  nand _37209_ (_05752_, _05751_, _05749_);
  nand _37210_ (_05753_, _00545_, _05739_);
  and _37211_ (_05755_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand _37212_ (_05756_, _24118_, _23594_);
  or _37213_ (_05757_, _24118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _37214_ (_05758_, _05757_, _05742_);
  and _37215_ (_05759_, _05758_, _05756_);
  nor _37216_ (_05760_, _05759_, _05755_);
  and _37217_ (_05761_, _05760_, _00257_);
  and _37218_ (_05762_, _05761_, _05753_);
  and _37219_ (_05763_, _01129_, _00256_);
  nor _37220_ (_05764_, _05763_, _05762_);
  nand _37221_ (_05765_, _05764_, _05752_);
  or _37222_ (_05766_, _05764_, _05752_);
  nand _37223_ (_05767_, _05766_, _05765_);
  nand _37224_ (_05768_, _26565_, _05739_);
  nor _37225_ (_05770_, _24678_, _23387_);
  nor _37226_ (_05771_, _05770_, _04418_);
  nor _37227_ (_05772_, _05771_, _05743_);
  and _37228_ (_05773_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _37229_ (_05774_, _05773_, _00256_);
  nor _37230_ (_05775_, _05774_, _05772_);
  nand _37231_ (_05776_, _05775_, _05768_);
  or _37232_ (_05777_, _00930_, _00257_);
  and _37233_ (_05778_, _05777_, _05776_);
  or _37234_ (_05779_, _00372_, _00263_);
  nor _37235_ (_05780_, _24067_, _23355_);
  nor _37236_ (_05781_, _05780_, _04398_);
  nor _37237_ (_05782_, _05781_, _05743_);
  and _37238_ (_05783_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _37239_ (_05785_, _05783_, _00256_);
  nor _37240_ (_05786_, _05785_, _05782_);
  nand _37241_ (_05787_, _05786_, _05779_);
  and _37242_ (_05789_, _00993_, _00256_);
  not _37243_ (_05790_, _05789_);
  nand _37244_ (_05791_, _05790_, _05787_);
  nand _37245_ (_05792_, _05791_, _05778_);
  or _37246_ (_05793_, _05791_, _05778_);
  nand _37247_ (_05794_, _05793_, _05792_);
  nand _37248_ (_05795_, _05794_, _05767_);
  or _37249_ (_05796_, _05794_, _05767_);
  nand _37250_ (_05797_, _05796_, _05795_);
  and _37251_ (_05798_, _00620_, _05739_);
  nor _37252_ (_05799_, _24296_, _23239_);
  or _37253_ (_05800_, _05799_, _24745_);
  and _37254_ (_05801_, _05800_, _05742_);
  and _37255_ (_05802_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _37256_ (_05803_, _05802_, _00256_);
  or _37257_ (_05805_, _05803_, _05801_);
  or _37258_ (_05806_, _05805_, _05798_);
  or _37259_ (_05807_, _01192_, _00257_);
  and _37260_ (_05808_, _05807_, _05806_);
  and _37261_ (_05809_, _00708_, _05739_);
  nand _37262_ (_05810_, _24125_, _23594_);
  or _37263_ (_05811_, _24125_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _37264_ (_05812_, _05811_, _05742_);
  and _37265_ (_05813_, _05812_, _05810_);
  and _37266_ (_05814_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _37267_ (_05816_, _05814_, _00256_);
  or _37268_ (_05817_, _05816_, _05813_);
  or _37269_ (_05818_, _05817_, _05809_);
  or _37270_ (_05819_, _01255_, _00257_);
  and _37271_ (_05820_, _05819_, _05818_);
  or _37272_ (_05821_, _05820_, _05808_);
  nand _37273_ (_05822_, _05820_, _05808_);
  nand _37274_ (_05823_, _05822_, _05821_);
  or _37275_ (_05824_, _00793_, _00263_);
  not _37276_ (_05826_, _24705_);
  nor _37277_ (_05827_, _05826_, _23594_);
  nor _37278_ (_05828_, _24705_, _23166_);
  nor _37279_ (_05829_, _05828_, _05827_);
  nor _37280_ (_05830_, _05829_, _05743_);
  and _37281_ (_05831_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _37282_ (_05832_, _05831_, _00256_);
  nor _37283_ (_05833_, _05832_, _05830_);
  and _37284_ (_05834_, _05833_, _05824_);
  and _37285_ (_05835_, _01318_, _00256_);
  or _37286_ (_05836_, _05835_, _05834_);
  and _37287_ (_05837_, _00875_, _05739_);
  not _37288_ (_05838_, _24654_);
  nor _37289_ (_05839_, _05838_, _23594_);
  nor _37290_ (_05840_, _24654_, _23126_);
  or _37291_ (_05841_, _05840_, _05839_);
  and _37292_ (_05843_, _05841_, _05742_);
  and _37293_ (_05844_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _37294_ (_05845_, _05844_, _00256_);
  or _37295_ (_05846_, _05845_, _05843_);
  or _37296_ (_05847_, _05846_, _05837_);
  or _37297_ (_05848_, _04299_, _00257_);
  and _37298_ (_05850_, _05848_, _05847_);
  or _37299_ (_05851_, _05850_, _05836_);
  nand _37300_ (_05852_, _05850_, _05836_);
  and _37301_ (_05853_, _05852_, _05851_);
  nand _37302_ (_05855_, _05853_, _05823_);
  or _37303_ (_05856_, _05853_, _05823_);
  nand _37304_ (_05857_, _05856_, _05855_);
  nand _37305_ (_05858_, _05857_, _05797_);
  or _37306_ (_05859_, _05857_, _05797_);
  and _37307_ (_05860_, _05859_, _05858_);
  nand _37308_ (_05861_, _05860_, _00168_);
  and _37309_ (_05863_, _00134_, _00099_);
  or _37310_ (_05864_, _00168_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _37311_ (_05865_, _05864_, _05863_);
  and _37312_ (_05866_, _05865_, _05861_);
  not _37313_ (_05867_, _00134_);
  nor _37314_ (_05868_, _05867_, _00099_);
  nor _37315_ (_05869_, _00168_, _00527_);
  and _37316_ (_05870_, _00168_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _37317_ (_05871_, _05870_, _05869_);
  and _37318_ (_05872_, _05871_, _05868_);
  or _37319_ (_05873_, _00168_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _37320_ (_05874_, _00134_, _00099_);
  not _37321_ (_05876_, _00168_);
  or _37322_ (_05877_, _05876_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _37323_ (_05878_, _05877_, _05874_);
  and _37324_ (_05879_, _05878_, _05873_);
  or _37325_ (_05880_, _00168_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _37326_ (_05881_, _05867_, _00099_);
  or _37327_ (_05882_, _05876_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _37328_ (_05883_, _05882_, _05881_);
  and _37329_ (_05884_, _05883_, _05880_);
  or _37330_ (_05885_, _05884_, _05879_);
  or _37331_ (_05886_, _05885_, _05872_);
  or _37332_ (_05887_, _05886_, _05866_);
  and _37333_ (_05888_, _05887_, _05738_);
  and _37334_ (_05889_, _00175_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  not _37335_ (_05890_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not _37336_ (_05891_, _00037_);
  and _37337_ (_05892_, _00058_, _26777_);
  and _37338_ (_05893_, _05892_, _05891_);
  and _37339_ (_05894_, _05893_, _05735_);
  nor _37340_ (_05895_, _05894_, _05890_);
  and _37341_ (_05896_, _05892_, _00037_);
  not _37342_ (_05897_, _05896_);
  nor _37343_ (_05898_, _05897_, _05735_);
  and _37344_ (_05900_, _26817_, _26777_);
  and _37345_ (_05901_, _05900_, _05891_);
  or _37346_ (_05903_, _05901_, _05737_);
  nor _37347_ (_05904_, _05903_, _05898_);
  and _37348_ (_05906_, _05904_, _05895_);
  nor _37349_ (_05908_, _00014_, _26817_);
  and _37350_ (_05909_, _05908_, _05737_);
  and _37351_ (_05910_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _37352_ (_05911_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _37353_ (_05912_, _05911_, _05910_);
  and _37354_ (_05913_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _37355_ (_05914_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or _37356_ (_05916_, _05914_, _05913_);
  or _37357_ (_05917_, _05916_, _05912_);
  and _37358_ (_05918_, _05917_, _05876_);
  and _37359_ (_05919_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _37360_ (_05920_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or _37361_ (_05921_, _05920_, _05919_);
  and _37362_ (_05922_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _37363_ (_05923_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _37364_ (_05924_, _05923_, _05922_);
  or _37365_ (_05925_, _05924_, _05921_);
  and _37366_ (_05926_, _05925_, _00168_);
  or _37367_ (_05927_, _05926_, _05918_);
  and _37368_ (_05928_, _05927_, _05909_);
  and _37369_ (_05929_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _37370_ (_05930_, _05929_, _05876_);
  and _37371_ (_05931_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _37372_ (_05932_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _37373_ (_05933_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _37374_ (_05934_, _05933_, _05932_);
  or _37375_ (_05935_, _05934_, _05931_);
  or _37376_ (_05936_, _05935_, _05930_);
  nor _37377_ (_05937_, _00058_, _00014_);
  and _37378_ (_05938_, _05937_, _05936_);
  and _37379_ (_05939_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _37380_ (_05940_, _05939_, _00168_);
  and _37381_ (_05941_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _37382_ (_05942_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _37383_ (_05943_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _37384_ (_05944_, _05943_, _05942_);
  or _37385_ (_05945_, _05944_, _05941_);
  or _37386_ (_05946_, _05945_, _05940_);
  and _37387_ (_05947_, _05946_, _05901_);
  and _37388_ (_05948_, _05947_, _05938_);
  or _37389_ (_05950_, _05948_, _05928_);
  or _37390_ (_05951_, _05950_, _05906_);
  or _37391_ (_05952_, _05951_, _05889_);
  and _37392_ (_05953_, _05734_, _26817_);
  and _37393_ (_05954_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _37394_ (_05955_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _37395_ (_05957_, _05955_, _05954_);
  and _37396_ (_05958_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _37397_ (_05959_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _37398_ (_05960_, _05959_, _05958_);
  or _37399_ (_05961_, _05960_, _05957_);
  and _37400_ (_05962_, _05961_, _05953_);
  and _37401_ (_05963_, _00014_, _26817_);
  and _37402_ (_05965_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _37403_ (_05966_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _37404_ (_05967_, _05966_, _05965_);
  and _37405_ (_05969_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _37406_ (_05970_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _37407_ (_05972_, _05970_, _05969_);
  or _37408_ (_05973_, _05972_, _05967_);
  and _37409_ (_05975_, _05973_, _05963_);
  or _37410_ (_05976_, _05975_, _05962_);
  and _37411_ (_05977_, _05976_, _00168_);
  and _37412_ (_05978_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _37413_ (_05979_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _37414_ (_05980_, _05979_, _05978_);
  and _37415_ (_05981_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _37416_ (_05982_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _37417_ (_05983_, _05982_, _05981_);
  or _37418_ (_05984_, _05983_, _05980_);
  and _37419_ (_05985_, _05984_, _05963_);
  and _37420_ (_05986_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _37421_ (_05988_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _37422_ (_05989_, _05988_, _05986_);
  and _37423_ (_05990_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _37424_ (_05992_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _37425_ (_05993_, _05992_, _05990_);
  or _37426_ (_05994_, _05993_, _05989_);
  and _37427_ (_05996_, _05994_, _05953_);
  or _37428_ (_05997_, _05996_, _05985_);
  and _37429_ (_05998_, _05997_, _05876_);
  or _37430_ (_05999_, _05998_, _05977_);
  and _37431_ (_06000_, _05999_, _05893_);
  and _37432_ (_06001_, _02397_, _00014_);
  and _37433_ (_06002_, _06001_, _05901_);
  and _37434_ (_06003_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and _37435_ (_06004_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _37436_ (_06005_, _06004_, _06003_);
  and _37437_ (_06006_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _37438_ (_06007_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _37439_ (_06008_, _06007_, _06006_);
  or _37440_ (_06010_, _06008_, _06005_);
  and _37441_ (_06011_, _06010_, _00168_);
  and _37442_ (_06012_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _37443_ (_06013_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _37444_ (_06014_, _06013_, _06012_);
  and _37445_ (_06015_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _37446_ (_06017_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _37447_ (_06018_, _06017_, _06015_);
  or _37448_ (_06019_, _06018_, _06014_);
  and _37449_ (_06020_, _06019_, _05876_);
  or _37450_ (_06021_, _06020_, _06011_);
  and _37451_ (_06022_, _06021_, _06002_);
  and _37452_ (_06024_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _37453_ (_06025_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _37454_ (_06026_, _06025_, _06024_);
  and _37455_ (_06027_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _37456_ (_06028_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _37457_ (_06029_, _06028_, _06027_);
  or _37458_ (_06030_, _06029_, _06026_);
  and _37459_ (_06032_, _06030_, _05876_);
  and _37460_ (_06033_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _37461_ (_06034_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _37462_ (_06035_, _06034_, _06033_);
  and _37463_ (_06036_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _37464_ (_06037_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _37465_ (_06038_, _06037_, _06036_);
  or _37466_ (_06039_, _06038_, _06035_);
  and _37467_ (_06040_, _06039_, _00168_);
  or _37468_ (_06042_, _06040_, _06032_);
  and _37469_ (_06043_, _06042_, _05894_);
  or _37470_ (_06044_, _06043_, _06022_);
  and _37471_ (_06045_, _05908_, _05896_);
  and _37472_ (_06046_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _37473_ (_06047_, _06046_, _05876_);
  and _37474_ (_06048_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _37475_ (_06049_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _37476_ (_06050_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _37477_ (_06052_, _06050_, _06049_);
  or _37478_ (_06053_, _06052_, _06048_);
  or _37479_ (_06054_, _06053_, _06047_);
  and _37480_ (_06055_, _05868_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _37481_ (_06056_, _06055_, _00168_);
  and _37482_ (_06057_, _05881_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _37483_ (_06058_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _37484_ (_06059_, _05874_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _37485_ (_06060_, _06059_, _06058_);
  or _37486_ (_06061_, _06060_, _06057_);
  or _37487_ (_06062_, _06061_, _06056_);
  and _37488_ (_06063_, _06062_, _06054_);
  and _37489_ (_06064_, _06063_, _06045_);
  or _37490_ (_06065_, _06064_, _06044_);
  or _37491_ (_06066_, _06065_, _06000_);
  or _37492_ (_06067_, _06066_, _05952_);
  or _37493_ (_06068_, _04982_, _26662_);
  or _37494_ (_06069_, _02254_, _26663_);
  or _37495_ (_06070_, _06069_, _24591_);
  and _37496_ (_06071_, _26625_, _24588_);
  or _37497_ (_06072_, _06071_, _04978_);
  and _37498_ (_06073_, _26625_, _24616_);
  or _37499_ (_06074_, _06073_, _02262_);
  or _37500_ (_06075_, _06074_, _06072_);
  or _37501_ (_06076_, _06075_, _26615_);
  or _37502_ (_06078_, _06076_, _06070_);
  or _37503_ (_06079_, _26620_, _24617_);
  and _37504_ (_06080_, _24618_, _24613_);
  or _37505_ (_06081_, _05063_, _06080_);
  or _37506_ (_06082_, _06081_, _06079_);
  or _37507_ (_06083_, _06082_, _06078_);
  or _37508_ (_06084_, _06083_, _06068_);
  or _37509_ (_06086_, _06084_, _26659_);
  and _37510_ (_06087_, _06086_, _26572_);
  or _37511_ (_06089_, _06087_, p2_in[1]);
  not _37512_ (_06090_, _06087_);
  or _37513_ (_06091_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _37514_ (_06092_, _06091_, _06089_);
  and _37515_ (_06094_, _06092_, _05881_);
  nor _37516_ (_06095_, _06087_, p2_in[0]);
  and _37517_ (_06096_, _06087_, _25336_);
  nor _37518_ (_06097_, _06096_, _06095_);
  and _37519_ (_06099_, _06097_, _05863_);
  or _37520_ (_06101_, _06099_, _06094_);
  or _37521_ (_06102_, _06087_, p2_in[2]);
  or _37522_ (_06104_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _37523_ (_06105_, _06104_, _06102_);
  and _37524_ (_06106_, _06105_, _05868_);
  or _37525_ (_06107_, _06087_, p2_in[3]);
  or _37526_ (_06108_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _37527_ (_06110_, _06108_, _06107_);
  and _37528_ (_06111_, _06110_, _05874_);
  or _37529_ (_06113_, _06111_, _06106_);
  or _37530_ (_06114_, _06113_, _06101_);
  and _37531_ (_06115_, _06114_, _05896_);
  or _37532_ (_06117_, _06087_, p3_in[3]);
  or _37533_ (_06118_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _37534_ (_06119_, _06118_, _06117_);
  and _37535_ (_06120_, _06119_, _05874_);
  or _37536_ (_06122_, _06087_, p3_in[1]);
  or _37537_ (_06124_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _37538_ (_06125_, _06124_, _06122_);
  and _37539_ (_06126_, _06125_, _05881_);
  or _37540_ (_06127_, _06126_, _06120_);
  or _37541_ (_06128_, _06087_, p3_in[2]);
  or _37542_ (_06129_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _37543_ (_06130_, _06129_, _06128_);
  and _37544_ (_06132_, _06130_, _05868_);
  nor _37545_ (_06133_, _06087_, p3_in[0]);
  and _37546_ (_06135_, _06087_, _25217_);
  nor _37547_ (_06136_, _06135_, _06133_);
  and _37548_ (_06137_, _06136_, _05863_);
  or _37549_ (_06138_, _06137_, _06132_);
  or _37550_ (_06139_, _06138_, _06127_);
  and _37551_ (_06140_, _06139_, _05737_);
  or _37552_ (_06142_, _06140_, _06115_);
  and _37553_ (_06143_, _06142_, _00168_);
  nor _37554_ (_06144_, _06087_, p3_in[6]);
  and _37555_ (_06145_, _06087_, _25234_);
  nor _37556_ (_06146_, _06145_, _06144_);
  and _37557_ (_06147_, _06146_, _05868_);
  nor _37558_ (_06148_, _06087_, p3_in[4]);
  not _37559_ (_06149_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _37560_ (_06150_, _06087_, _06149_);
  nor _37561_ (_06152_, _06150_, _06148_);
  and _37562_ (_06153_, _06152_, _05863_);
  or _37563_ (_06154_, _06153_, _06147_);
  or _37564_ (_06155_, _06087_, p3_in[7]);
  or _37565_ (_06156_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _37566_ (_06157_, _06156_, _06155_);
  and _37567_ (_06158_, _06157_, _05874_);
  or _37568_ (_06159_, _06087_, p3_in[5]);
  or _37569_ (_06161_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _37570_ (_06162_, _06161_, _06159_);
  and _37571_ (_06164_, _06162_, _05881_);
  or _37572_ (_06165_, _06164_, _06158_);
  or _37573_ (_06166_, _06165_, _06154_);
  and _37574_ (_06167_, _06166_, _05737_);
  or _37575_ (_06169_, _06087_, p2_in[5]);
  or _37576_ (_06172_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _37577_ (_06173_, _06172_, _06169_);
  and _37578_ (_06174_, _06173_, _05881_);
  nor _37579_ (_06175_, _06087_, p2_in[4]);
  and _37580_ (_06177_, _06087_, _25300_);
  nor _37581_ (_06179_, _06177_, _06175_);
  and _37582_ (_06181_, _06179_, _05863_);
  or _37583_ (_06182_, _06181_, _06174_);
  nor _37584_ (_06183_, _06087_, p2_in[6]);
  not _37585_ (_06185_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _37586_ (_06186_, _06087_, _06185_);
  nor _37587_ (_06187_, _06186_, _06183_);
  and _37588_ (_06188_, _06187_, _05868_);
  or _37589_ (_06189_, _06087_, p2_in[7]);
  or _37590_ (_06190_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _37591_ (_06191_, _06190_, _06189_);
  and _37592_ (_06192_, _06191_, _05874_);
  or _37593_ (_06193_, _06192_, _06188_);
  or _37594_ (_06194_, _06193_, _06182_);
  and _37595_ (_06195_, _06194_, _05896_);
  or _37596_ (_06196_, _06195_, _06167_);
  and _37597_ (_06197_, _06196_, _05876_);
  or _37598_ (_06198_, _06197_, _06143_);
  and _37599_ (_06199_, _06198_, _05953_);
  or _37600_ (_06200_, _06087_, p0_in[1]);
  or _37601_ (_06201_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _37602_ (_06202_, _06201_, _06200_);
  and _37603_ (_06203_, _06202_, _05881_);
  nor _37604_ (_06204_, _06087_, p0_in[0]);
  and _37605_ (_06206_, _06087_, _25483_);
  nor _37606_ (_06207_, _06206_, _06204_);
  and _37607_ (_06208_, _06207_, _05863_);
  or _37608_ (_06209_, _06208_, _06203_);
  or _37609_ (_06210_, _06087_, p0_in[2]);
  or _37610_ (_06211_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _37611_ (_06212_, _06211_, _06210_);
  and _37612_ (_06213_, _06212_, _05868_);
  or _37613_ (_06214_, _06087_, p0_in[3]);
  or _37614_ (_06215_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _37615_ (_06216_, _06215_, _06214_);
  and _37616_ (_06217_, _06216_, _05874_);
  or _37617_ (_06218_, _06217_, _06213_);
  or _37618_ (_06219_, _06218_, _06209_);
  and _37619_ (_06220_, _06219_, _05896_);
  or _37620_ (_06221_, _06087_, p1_in[2]);
  or _37621_ (_06222_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _37622_ (_06223_, _06222_, _06221_);
  and _37623_ (_06224_, _06223_, _05868_);
  or _37624_ (_06225_, _06087_, p1_in[3]);
  or _37625_ (_06226_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _37626_ (_06227_, _06226_, _06225_);
  and _37627_ (_06228_, _06227_, _05874_);
  or _37628_ (_06229_, _06228_, _06224_);
  or _37629_ (_06230_, _06087_, p1_in[1]);
  or _37630_ (_06231_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _37631_ (_06232_, _06231_, _06230_);
  and _37632_ (_06234_, _06232_, _05881_);
  nor _37633_ (_06235_, _06087_, p1_in[0]);
  and _37634_ (_06236_, _06087_, _25400_);
  nor _37635_ (_06237_, _06236_, _06235_);
  and _37636_ (_06238_, _06237_, _05863_);
  or _37637_ (_06239_, _06238_, _06234_);
  or _37638_ (_06240_, _06239_, _06229_);
  and _37639_ (_06241_, _06240_, _05737_);
  or _37640_ (_06242_, _06241_, _06220_);
  and _37641_ (_06243_, _06242_, _00168_);
  or _37642_ (_06244_, _06087_, p1_in[5]);
  or _37643_ (_06245_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _37644_ (_06246_, _06245_, _06244_);
  and _37645_ (_06247_, _06246_, _05881_);
  nor _37646_ (_06248_, _06087_, p1_in[4]);
  not _37647_ (_06249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _37648_ (_06250_, _06087_, _06249_);
  nor _37649_ (_06251_, _06250_, _06248_);
  and _37650_ (_06252_, _06251_, _05863_);
  or _37651_ (_06253_, _06252_, _06247_);
  nor _37652_ (_06255_, _06087_, p1_in[6]);
  and _37653_ (_06256_, _06087_, _25418_);
  nor _37654_ (_06258_, _06256_, _06255_);
  and _37655_ (_06259_, _06258_, _05868_);
  or _37656_ (_06260_, _06087_, p1_in[7]);
  or _37657_ (_06261_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _37658_ (_06262_, _06261_, _06260_);
  and _37659_ (_06263_, _06262_, _05874_);
  or _37660_ (_06265_, _06263_, _06259_);
  or _37661_ (_06266_, _06265_, _06253_);
  and _37662_ (_06268_, _06266_, _05737_);
  or _37663_ (_06269_, _06087_, p0_in[5]);
  or _37664_ (_06270_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _37665_ (_06272_, _06270_, _06269_);
  and _37666_ (_06274_, _06272_, _05881_);
  nor _37667_ (_06275_, _06087_, p0_in[4]);
  and _37668_ (_06277_, _06087_, _25531_);
  nor _37669_ (_06278_, _06277_, _06275_);
  and _37670_ (_06279_, _06278_, _05863_);
  or _37671_ (_06281_, _06279_, _06274_);
  nor _37672_ (_06282_, _06087_, p0_in[6]);
  and _37673_ (_06283_, _06087_, _25517_);
  nor _37674_ (_06284_, _06283_, _06282_);
  and _37675_ (_06285_, _06284_, _05868_);
  or _37676_ (_06286_, _06087_, p0_in[7]);
  or _37677_ (_06287_, _06090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _37678_ (_06288_, _06287_, _06286_);
  and _37679_ (_06290_, _06288_, _05874_);
  or _37680_ (_06291_, _06290_, _06285_);
  or _37681_ (_06292_, _06291_, _06281_);
  and _37682_ (_06294_, _06292_, _05896_);
  or _37683_ (_06295_, _06294_, _06268_);
  and _37684_ (_06296_, _06295_, _05876_);
  or _37685_ (_06297_, _06296_, _06243_);
  and _37686_ (_06298_, _06297_, _05963_);
  or _37687_ (_06299_, _06298_, _06199_);
  or _37688_ (_06300_, _06299_, _06067_);
  or _37689_ (_06301_, _06300_, _05888_);
  and _37690_ (_06302_, _06045_, _00260_);
  nor _37691_ (_06303_, _06302_, _00184_);
  nand _37692_ (_06304_, _05889_, _23594_);
  and _37693_ (_06305_, _06304_, _06303_);
  and _37694_ (_06306_, _06305_, _06301_);
  and _37695_ (_06307_, _05868_, _23816_);
  or _37696_ (_06308_, _06307_, _05876_);
  and _37697_ (_06309_, _05863_, _24685_);
  and _37698_ (_06310_, _05881_, _23892_);
  and _37699_ (_06311_, _05874_, _23738_);
  or _37700_ (_06312_, _06311_, _06310_);
  or _37701_ (_06313_, _06312_, _06309_);
  or _37702_ (_06314_, _06313_, _06308_);
  and _37703_ (_06315_, _05868_, _24043_);
  or _37704_ (_06316_, _06315_, _00168_);
  and _37705_ (_06317_, _05863_, _23642_);
  and _37706_ (_06318_, _05881_, _23939_);
  and _37707_ (_06319_, _05874_, _26750_);
  or _37708_ (_06320_, _06319_, _06318_);
  or _37709_ (_06321_, _06320_, _06317_);
  or _37710_ (_06322_, _06321_, _06316_);
  nand _37711_ (_06323_, _06322_, _06314_);
  nor _37712_ (_06324_, _06323_, _06303_);
  or _37713_ (_06325_, _06324_, _06306_);
  and _37714_ (_27305_, _06325_, _22762_);
  nor _37715_ (_06327_, _26817_, _02444_);
  and _37716_ (_06328_, _00168_, _00037_);
  and _37717_ (_06329_, _06328_, _05863_);
  nor _37718_ (_06330_, _02397_, _00014_);
  and _37719_ (_06331_, _06330_, _06329_);
  and _37720_ (_06333_, _06331_, _06327_);
  and _37721_ (_06334_, _06333_, _00260_);
  not _37722_ (_06335_, _24646_);
  and _37723_ (_06336_, _05874_, _05876_);
  nor _37724_ (_06337_, _06336_, _06335_);
  and _37725_ (_06339_, _06337_, _00065_);
  nor _37726_ (_06340_, _06339_, _06334_);
  and _37727_ (_06341_, _06340_, _00178_);
  and _37728_ (_06343_, _00259_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _37729_ (_06344_, _05963_, _05892_);
  and _37730_ (_06345_, _06328_, _05874_);
  and _37731_ (_06346_, _06345_, _06344_);
  and _37732_ (_06347_, _06346_, _06343_);
  not _37733_ (_06348_, _06347_);
  and _37734_ (_06349_, _06333_, _00256_);
  and _37735_ (_06350_, _06329_, _06001_);
  and _37736_ (_06351_, _06350_, _06327_);
  and _37737_ (_06352_, _06351_, _00278_);
  nor _37738_ (_06353_, _06352_, _06349_);
  and _37739_ (_06354_, _06353_, _06348_);
  nor _37740_ (_06355_, _06354_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _37741_ (_06356_, _06355_);
  and _37742_ (_06357_, _06356_, _06341_);
  and _37743_ (_06358_, _06344_, _05868_);
  and _37744_ (_06359_, _06358_, _06328_);
  and _37745_ (_06361_, _06359_, _06343_);
  or _37746_ (_06362_, _06361_, rst);
  nor _37747_ (_27306_, _06362_, _06357_);
  and _37748_ (_06363_, _05892_, _05735_);
  and _37749_ (_06365_, _00168_, _05891_);
  and _37750_ (_06366_, _06365_, _05863_);
  and _37751_ (_06367_, _06366_, _06363_);
  nor _37752_ (_06369_, _00168_, _00037_);
  and _37753_ (_06371_, _06369_, _05863_);
  and _37754_ (_06372_, _06371_, _06363_);
  or _37755_ (_06373_, _06372_, _06367_);
  and _37756_ (_06374_, _06365_, _05868_);
  and _37757_ (_06375_, _06374_, _06363_);
  and _37758_ (_06376_, _06369_, _05881_);
  and _37759_ (_06377_, _06376_, _06363_);
  or _37760_ (_06378_, _06377_, _06375_);
  nor _37761_ (_06379_, _06378_, _06373_);
  and _37762_ (_06380_, _06330_, _05900_);
  and _37763_ (_06381_, _06380_, _06366_);
  and _37764_ (_06382_, _06336_, _00037_);
  and _37765_ (_06383_, _05937_, _05900_);
  and _37766_ (_06384_, _06383_, _06382_);
  nor _37767_ (_06385_, _06384_, _06381_);
  and _37768_ (_06387_, _06366_, _06344_);
  and _37769_ (_06388_, _06365_, _05874_);
  and _37770_ (_06389_, _06388_, _06363_);
  nor _37771_ (_06390_, _06389_, _06387_);
  and _37772_ (_06392_, _06390_, _06385_);
  and _37773_ (_06393_, _06392_, _06379_);
  and _37774_ (_06394_, _06388_, _06344_);
  and _37775_ (_06396_, _06365_, _05881_);
  and _37776_ (_06397_, _06396_, _06344_);
  nor _37777_ (_06399_, _06397_, _06394_);
  and _37778_ (_06400_, _06376_, _06344_);
  and _37779_ (_06402_, _06374_, _06344_);
  nor _37780_ (_06404_, _06402_, _06400_);
  and _37781_ (_06405_, _06404_, _06399_);
  and _37782_ (_06406_, _06371_, _06344_);
  and _37783_ (_06407_, _06382_, _06344_);
  nor _37784_ (_06408_, _06407_, _06406_);
  and _37785_ (_06409_, _05963_, _05736_);
  and _37786_ (_06410_, _06409_, _06396_);
  and _37787_ (_06411_, _06409_, _06366_);
  nor _37788_ (_06412_, _06411_, _06410_);
  and _37789_ (_06413_, _06412_, _06408_);
  and _37790_ (_06414_, _06413_, _06405_);
  and _37791_ (_06416_, _06414_, _06393_);
  or _37792_ (_06417_, _06351_, _06333_);
  and _37793_ (_06418_, _06329_, _05900_);
  or _37794_ (_06419_, _06359_, _06346_);
  and _37795_ (_06420_, _06344_, _05881_);
  and _37796_ (_06421_, _06420_, _06328_);
  and _37797_ (_06422_, _05937_, _06327_);
  and _37798_ (_06423_, _06422_, _06329_);
  or _37799_ (_06424_, _06423_, _06421_);
  or _37800_ (_06425_, _06424_, _06419_);
  or _37801_ (_06426_, _06425_, _06418_);
  nor _37802_ (_06427_, _06426_, _06417_);
  and _37803_ (_06428_, _06427_, _06416_);
  not _37804_ (_06429_, _06428_);
  and _37805_ (_06431_, _06429_, _06357_);
  not _37806_ (_06432_, _06431_);
  and _37807_ (_06433_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _37808_ (_06434_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _37809_ (_06435_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _37810_ (_06436_, _06435_, _06434_);
  and _37811_ (_06437_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _37812_ (_06438_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _37813_ (_06439_, _06438_, _06437_);
  or _37814_ (_06441_, _06439_, _06436_);
  and _37815_ (_06442_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _37816_ (_06443_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or _37817_ (_06444_, _06443_, _06442_);
  and _37818_ (_06445_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _37819_ (_06447_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _37820_ (_06448_, _06447_, _06445_);
  or _37821_ (_06449_, _06448_, _06444_);
  or _37822_ (_06451_, _06449_, _06441_);
  and _37823_ (_06452_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _37824_ (_06453_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or _37825_ (_06454_, _06453_, _06452_);
  and _37826_ (_06455_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _37827_ (_06456_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _37828_ (_06458_, _06456_, _06455_);
  or _37829_ (_06459_, _06458_, _06454_);
  and _37830_ (_06460_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and _37831_ (_06462_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _37832_ (_06463_, _06462_, _06460_);
  and _37833_ (_06464_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _37834_ (_06465_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _37835_ (_06466_, _06465_, _06464_);
  or _37836_ (_06467_, _06466_, _06463_);
  or _37837_ (_06469_, _06467_, _06459_);
  or _37838_ (_06471_, _06469_, _06451_);
  and _37839_ (_06472_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _37840_ (_06474_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or _37841_ (_06475_, _06474_, _06472_);
  and _37842_ (_06476_, _06421_, _26727_);
  and _37843_ (_06477_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or _37844_ (_06478_, _06477_, _06476_);
  or _37845_ (_06479_, _06478_, _06475_);
  and _37846_ (_06480_, _06418_, _05937_);
  and _37847_ (_06481_, _06480_, _06157_);
  and _37848_ (_06482_, _06331_, _05900_);
  and _37849_ (_06483_, _06482_, _06191_);
  or _37850_ (_06485_, _06483_, _06481_);
  and _37851_ (_06486_, _06344_, _06329_);
  and _37852_ (_06487_, _06486_, _06288_);
  and _37853_ (_06488_, _06409_, _06329_);
  and _37854_ (_06489_, _06488_, _06262_);
  or _37855_ (_06490_, _06489_, _06487_);
  or _37856_ (_06491_, _06490_, _06485_);
  or _37857_ (_06493_, _06491_, _06479_);
  and _37858_ (_06494_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _37859_ (_06495_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _37860_ (_06496_, _06495_, _06494_);
  or _37861_ (_06497_, _06496_, _06493_);
  or _37862_ (_06498_, _06497_, _06471_);
  and _37863_ (_06499_, _06498_, _06357_);
  or _37864_ (_06500_, _06499_, _06361_);
  or _37865_ (_06501_, _06500_, _06433_);
  not _37866_ (_06502_, _06361_);
  or _37867_ (_06503_, _06502_, _00875_);
  and _37868_ (_06504_, _06503_, _22762_);
  and _37869_ (_27307_[7], _06504_, _06501_);
  and _37870_ (_06505_, _23753_, _22946_);
  and _37871_ (_06506_, _06505_, _23661_);
  and _37872_ (_06507_, _06506_, _24010_);
  not _37873_ (_06508_, _06507_);
  and _37874_ (_06509_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and _37875_ (_06510_, _06507_, _23898_);
  or _37876_ (_25285_, _06510_, _06509_);
  and _37877_ (_06511_, _02325_, _23656_);
  and _37878_ (_06513_, _06511_, _24050_);
  not _37879_ (_06514_, _06511_);
  and _37880_ (_06515_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or _37881_ (_25288_, _06515_, _06513_);
  and _37882_ (_06517_, _02325_, _25078_);
  and _37883_ (_06518_, _06517_, _23824_);
  not _37884_ (_06520_, _06517_);
  and _37885_ (_06522_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or _37886_ (_27151_, _06522_, _06518_);
  and _37887_ (_06524_, _02325_, _24282_);
  and _37888_ (_06525_, _06524_, _23649_);
  not _37889_ (_06527_, _06524_);
  and _37890_ (_06529_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  or _37891_ (_25295_, _06529_, _06525_);
  and _37892_ (_06530_, _02325_, _23911_);
  and _37893_ (_06531_, _06530_, _23898_);
  not _37894_ (_06532_, _06530_);
  and _37895_ (_06533_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  or _37896_ (_25298_, _06533_, _06531_);
  and _37897_ (_06534_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and _37898_ (_06536_, _05705_, _23747_);
  or _37899_ (_25344_, _06536_, _06534_);
  and _37900_ (_06538_, _05429_, _23778_);
  and _37901_ (_06539_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or _37902_ (_25347_, _06539_, _06538_);
  and _37903_ (_06540_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and _37904_ (_06541_, _05705_, _23824_);
  or _37905_ (_25351_, _06541_, _06540_);
  and _37906_ (_06544_, _02325_, _24010_);
  and _37907_ (_06545_, _06544_, _23946_);
  not _37908_ (_06547_, _06544_);
  and _37909_ (_06548_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or _37910_ (_25357_, _06548_, _06545_);
  and _37911_ (_06550_, _06544_, _23778_);
  and _37912_ (_06551_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or _37913_ (_25366_, _06551_, _06550_);
  and _37914_ (_06552_, _02325_, _24085_);
  and _37915_ (_06553_, _06552_, _23898_);
  not _37916_ (_06554_, _06552_);
  and _37917_ (_06555_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or _37918_ (_27143_, _06555_, _06553_);
  and _37919_ (_06557_, _05454_, _23778_);
  and _37920_ (_06558_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _37921_ (_25392_, _06558_, _06557_);
  and _37922_ (_06559_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and _37923_ (_06561_, _05705_, _23707_);
  or _37924_ (_25413_, _06561_, _06559_);
  and _37925_ (_06563_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and _37926_ (_06564_, _05705_, _24050_);
  or _37927_ (_25424_, _06564_, _06563_);
  and _37928_ (_06566_, _24581_, _26650_);
  or _37929_ (_06567_, _02261_, _23950_);
  or _37930_ (_06568_, _06567_, _06566_);
  nor _37931_ (_06569_, _06568_, _24595_);
  nand _37932_ (_06570_, _06569_, _24543_);
  or _37933_ (_06572_, _05087_, _05090_);
  or _37934_ (_06573_, _06572_, _26662_);
  or _37935_ (_06574_, _06573_, _06570_);
  or _37936_ (_06575_, _26654_, _26644_);
  or _37937_ (_06576_, _06575_, _04952_);
  or _37938_ (_06577_, _03276_, _26651_);
  and _37939_ (_06578_, _26645_, _24448_);
  or _37940_ (_06579_, _06578_, _04959_);
  or _37941_ (_06580_, _06579_, _06577_);
  or _37942_ (_06581_, _06580_, _06576_);
  or _37943_ (_06582_, _06581_, _06574_);
  or _37944_ (_06583_, _06582_, _04989_);
  or _37945_ (_06584_, _24559_, _26572_);
  or _37946_ (_06586_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _22766_);
  and _37947_ (_06587_, _06586_, _22762_);
  and _37948_ (_06588_, _06587_, _06584_);
  and _37949_ (_26871_[0], _06588_, _06583_);
  and _37950_ (_06589_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and _37951_ (_06590_, _05705_, _23946_);
  or _37952_ (_25428_, _06590_, _06589_);
  and _37953_ (_06592_, _05454_, _23824_);
  and _37954_ (_06593_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or _37955_ (_25436_, _06593_, _06592_);
  and _37956_ (_06594_, _05042_, _23747_);
  and _37957_ (_06596_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or _37958_ (_25440_, _06596_, _06594_);
  nor _37959_ (_26897_[3], _00566_, rst);
  and _37960_ (_06597_, _05454_, _23898_);
  and _37961_ (_06598_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _37962_ (_25452_, _06598_, _06597_);
  and _37963_ (_06599_, _23778_, _23665_);
  and _37964_ (_06600_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or _37965_ (_25454_, _06600_, _06599_);
  and _37966_ (_06602_, _02325_, _23069_);
  and _37967_ (_06603_, _06602_, _23649_);
  not _37968_ (_06604_, _06602_);
  and _37969_ (_06605_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  or _37970_ (_25457_, _06605_, _06603_);
  and _37971_ (_06606_, _06602_, _23898_);
  and _37972_ (_06607_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  or _37973_ (_25458_, _06607_, _06606_);
  and _37974_ (_06608_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  and _37975_ (_06609_, _05354_, _23747_);
  or _37976_ (_25463_, _06609_, _06608_);
  and _37977_ (_06610_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  and _37978_ (_06612_, _05354_, _23946_);
  or _37979_ (_25465_, _06612_, _06610_);
  and _37980_ (_06613_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  and _37981_ (_06614_, _05354_, _23649_);
  or _37982_ (_25471_, _06614_, _06613_);
  and _37983_ (_06615_, _01758_, _24085_);
  and _37984_ (_06616_, _06615_, _23649_);
  not _37985_ (_06618_, _06615_);
  and _37986_ (_06619_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or _37987_ (_25478_, _06619_, _06616_);
  and _37988_ (_06620_, _06615_, _23747_);
  and _37989_ (_06621_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or _37990_ (_25487_, _06621_, _06620_);
  and _37991_ (_06622_, _02326_, _24050_);
  and _37992_ (_06623_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or _37993_ (_25492_, _06623_, _06622_);
  and _37994_ (_06624_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  and _37995_ (_06625_, _05354_, _23707_);
  or _37996_ (_25513_, _06625_, _06624_);
  nor _37997_ (_26887_[6], _26811_, rst);
  and _37998_ (_06626_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and _37999_ (_06627_, _05705_, _23778_);
  or _38000_ (_25522_, _06627_, _06626_);
  and _38001_ (_06628_, _06615_, _24050_);
  and _38002_ (_06629_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or _38003_ (_27082_, _06629_, _06628_);
  and _38004_ (_06630_, _06615_, _23946_);
  and _38005_ (_06632_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or _38006_ (_25535_, _06632_, _06630_);
  or _38007_ (_06634_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and _38008_ (_26915_, _06634_, _05209_);
  and _38009_ (_06636_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  and _38010_ (_06637_, _05354_, _23898_);
  or _38011_ (_25567_, _06637_, _06636_);
  and _38012_ (_06639_, _02325_, _24275_);
  and _38013_ (_06641_, _06639_, _23747_);
  not _38014_ (_06643_, _06639_);
  and _38015_ (_06644_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or _38016_ (_25569_, _06644_, _06641_);
  and _38017_ (_06646_, _02325_, _24005_);
  and _38018_ (_06647_, _06646_, _23747_);
  not _38019_ (_06649_, _06646_);
  and _38020_ (_06650_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or _38021_ (_25575_, _06650_, _06647_);
  nor _38022_ (_26897_[6], _00814_, rst);
  and _38023_ (_06651_, _02325_, _23752_);
  and _38024_ (_06652_, _06651_, _23946_);
  not _38025_ (_06653_, _06651_);
  and _38026_ (_06654_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  or _38027_ (_25578_, _06654_, _06652_);
  and _38028_ (_06655_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  and _38029_ (_06656_, _04748_, _23824_);
  or _38030_ (_25580_, _06656_, _06655_);
  and _38031_ (_06657_, _24852_, _23747_);
  and _38032_ (_06658_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  or _38033_ (_27205_, _06658_, _06657_);
  and _38034_ (_06659_, _06615_, _23778_);
  and _38035_ (_06661_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or _38036_ (_25585_, _06661_, _06659_);
  and _38037_ (_06662_, _06511_, _23778_);
  and _38038_ (_06663_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or _38039_ (_25589_, _06663_, _06662_);
  and _38040_ (_06665_, _24275_, _23664_);
  and _38041_ (_06666_, _06665_, _23824_);
  not _38042_ (_06667_, _06665_);
  and _38043_ (_06668_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  or _38044_ (_27088_, _06668_, _06666_);
  and _38045_ (_06669_, _06665_, _23898_);
  and _38046_ (_06670_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  or _38047_ (_25600_, _06670_, _06669_);
  and _38048_ (_06671_, _06665_, _23778_);
  and _38049_ (_06672_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or _38050_ (_25606_, _06672_, _06671_);
  or _38051_ (_06673_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and _38052_ (_25614_, _06673_, _05467_);
  or _38053_ (_06674_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and _38054_ (_25617_, _06674_, _05463_);
  and _38055_ (_06675_, _24593_, _24448_);
  or _38056_ (_06676_, _04978_, _24591_);
  or _38057_ (_06677_, _06676_, _05067_);
  or _38058_ (_06678_, _06677_, _06675_);
  or _38059_ (_06680_, _26652_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _38060_ (_06681_, _06680_, _24587_);
  or _38061_ (_06682_, _26665_, _24559_);
  or _38062_ (_06683_, _06682_, _06681_);
  or _38063_ (_06685_, _06683_, _06678_);
  and _38064_ (_06686_, _04973_, _24445_);
  and _38065_ (_06687_, _24606_, _24447_);
  or _38066_ (_06688_, _06687_, _04970_);
  or _38067_ (_06690_, _06688_, _06686_);
  or _38068_ (_06691_, _06690_, _06068_);
  or _38069_ (_06692_, _06691_, _06685_);
  and _38070_ (_06693_, _26614_, _24556_);
  or _38071_ (_06694_, _06693_, _03316_);
  or _38072_ (_06696_, _06694_, _05088_);
  or _38073_ (_06697_, _26599_, _24617_);
  or _38074_ (_06698_, _04969_, _04947_);
  or _38075_ (_06699_, _06698_, _06697_);
  or _38076_ (_06700_, _06699_, _06696_);
  or _38077_ (_06701_, _06700_, _06692_);
  or _38078_ (_06703_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _22766_);
  and _38079_ (_06704_, _06703_, _22762_);
  and _38080_ (_06706_, _06704_, _06584_);
  and _38081_ (_26871_[1], _06706_, _06701_);
  and _38082_ (_06708_, _25733_, _23898_);
  and _38083_ (_06710_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or _38084_ (_25628_, _06710_, _06708_);
  and _38085_ (_06712_, _05042_, _23707_);
  and _38086_ (_06713_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or _38087_ (_25632_, _06713_, _06712_);
  and _38088_ (_06715_, _06665_, _23946_);
  and _38089_ (_06716_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or _38090_ (_25637_, _06716_, _06715_);
  and _38091_ (_06717_, _06665_, _23649_);
  and _38092_ (_06718_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  or _38093_ (_25643_, _06718_, _06717_);
  or _38094_ (_06719_, _03274_, _26665_);
  or _38095_ (_06720_, _05089_, _02381_);
  or _38096_ (_06722_, _06720_, _06719_);
  or _38097_ (_06723_, _04982_, _24617_);
  or _38098_ (_06724_, _06723_, _06676_);
  and _38099_ (_06725_, _24616_, _24448_);
  or _38100_ (_06726_, _26661_, _24585_);
  or _38101_ (_06727_, _06726_, _06725_);
  or _38102_ (_06728_, _06727_, _06724_);
  or _38103_ (_06729_, _06728_, _06690_);
  or _38104_ (_06730_, _06729_, _06694_);
  or _38105_ (_06731_, _06730_, _06722_);
  and _38106_ (_06732_, _06731_, _22768_);
  and _38107_ (_06733_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _38108_ (_06734_, _24558_, _22766_);
  or _38109_ (_06735_, _06734_, _06733_);
  or _38110_ (_06736_, _06735_, _06732_);
  and _38111_ (_26871_[2], _06736_, _22762_);
  or _38112_ (_06737_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and _38113_ (_25648_, _06737_, _05478_);
  and _38114_ (_06738_, _02326_, _23946_);
  and _38115_ (_06739_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or _38116_ (_27153_, _06739_, _06738_);
  and _38117_ (_06740_, _06665_, _23747_);
  and _38118_ (_06741_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  or _38119_ (_25655_, _06741_, _06740_);
  or _38120_ (_06743_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and _38121_ (_25658_, _06743_, _05474_);
  and _38122_ (_06746_, _05701_, _23649_);
  and _38123_ (_06747_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or _38124_ (_25670_, _06747_, _06746_);
  and _38125_ (_06749_, _05714_, _24050_);
  and _38126_ (_06750_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  or _38127_ (_25673_, _06750_, _06749_);
  and _38128_ (_06751_, _23898_, _23665_);
  and _38129_ (_06753_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  or _38130_ (_25732_, _06753_, _06751_);
  and _38131_ (_06755_, _02325_, _23986_);
  and _38132_ (_06756_, _06755_, _23778_);
  not _38133_ (_06757_, _06755_);
  and _38134_ (_06759_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or _38135_ (_25747_, _06759_, _06756_);
  and _38136_ (_06761_, _02359_, _23824_);
  and _38137_ (_06763_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  or _38138_ (_25758_, _06763_, _06761_);
  and _38139_ (_06764_, _05701_, _23707_);
  and _38140_ (_06766_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or _38141_ (_25767_, _06766_, _06764_);
  and _38142_ (_06768_, _05701_, _24050_);
  and _38143_ (_06769_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or _38144_ (_25768_, _06769_, _06768_);
  and _38145_ (_06771_, _06651_, _24050_);
  and _38146_ (_06772_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  or _38147_ (_25771_, _06772_, _06771_);
  not _38148_ (_06773_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _38149_ (_06774_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not _38150_ (_06775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor _38151_ (_06776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _38152_ (_06778_, _06776_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and _38153_ (_06779_, _06778_, _06775_);
  and _38154_ (_06780_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _04488_);
  or _38155_ (_06781_, _06780_, _06779_);
  nor _38156_ (_06783_, _06781_, _06774_);
  nand _38157_ (_06785_, _06783_, _06773_);
  nor _38158_ (_06786_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor _38159_ (_06788_, _06786_, _06783_);
  nand _38160_ (_06789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _38161_ (_06791_, _06789_, _06788_);
  and _38162_ (_06792_, _06791_, _22762_);
  and _38163_ (_25778_, _06792_, _06785_);
  not _38164_ (_06795_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  and _38165_ (_06796_, _04449_, _06795_);
  and _38166_ (_06797_, _04567_, _04454_);
  and _38167_ (_06798_, _06797_, _06796_);
  and _38168_ (_06799_, _06798_, _04563_);
  not _38169_ (_06800_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or _38170_ (_06801_, _04569_, _06800_);
  nor _38171_ (_06803_, _06801_, _06799_);
  or _38172_ (_06804_, _06803_, _04462_);
  and _38173_ (_25781_, _06804_, _22762_);
  nand _38174_ (_06805_, _24504_, _24399_);
  nor _38175_ (_06806_, _06805_, _24461_);
  and _38176_ (_06807_, _22765_, _23839_);
  nand _38177_ (_06808_, _06807_, _25644_);
  nor _38178_ (_06809_, _06808_, _23863_);
  and _38179_ (_06810_, _24526_, _24482_);
  and _38180_ (_06811_, _06810_, _06809_);
  and _38181_ (_06813_, _24431_, _24349_);
  and _38182_ (_06814_, _06813_, _06811_);
  and _38183_ (_26898_, _06814_, _06806_);
  and _38184_ (_25786_, _06788_, _22762_);
  and _38185_ (_06815_, _05410_, _24050_);
  and _38186_ (_06816_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  or _38187_ (_25792_, _06816_, _06815_);
  and _38188_ (_06817_, _04457_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  or _38189_ (_06818_, _06817_, _04462_);
  nor _38190_ (_06819_, _04490_, rst);
  and _38191_ (_25796_, _06819_, _06818_);
  or _38192_ (_06820_, _04780_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand _38193_ (_06821_, _04780_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _38194_ (_06822_, _06821_, _06820_);
  nand _38195_ (_06823_, _06822_, _22762_);
  nor _38196_ (_25800_, _06823_, _04462_);
  not _38197_ (_06825_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _38198_ (_06826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _38199_ (_06827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _38200_ (_06828_, _06778_, _06827_);
  or _38201_ (_06829_, _06828_, _06780_);
  nor _38202_ (_06830_, _06829_, _06826_);
  nand _38203_ (_06832_, _06830_, _06825_);
  nor _38204_ (_06834_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor _38205_ (_06835_, _06834_, _06830_);
  nand _38206_ (_06836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand _38207_ (_06838_, _06836_, _06835_);
  and _38208_ (_06839_, _06838_, _22762_);
  and _38209_ (_25814_, _06839_, _06832_);
  and _38210_ (_25815_, _06835_, _22762_);
  and _38211_ (_06840_, _06665_, _23707_);
  and _38212_ (_06841_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  or _38213_ (_25819_, _06841_, _06840_);
  and _38214_ (_06842_, _04917_, _23898_);
  and _38215_ (_06843_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or _38216_ (_27108_, _06843_, _06842_);
  not _38217_ (_06845_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not _38218_ (_06846_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _38219_ (_06847_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _06846_);
  not _38220_ (_06848_, _06847_);
  nor _38221_ (_06849_, _04376_, _04609_);
  and _38222_ (_06850_, _06849_, _06848_);
  and _38223_ (_06851_, _06850_, _04628_);
  nor _38224_ (_06852_, _06851_, _06845_);
  and _38225_ (_06853_, _06851_, rxd_i);
  or _38226_ (_06854_, _06853_, rst);
  or _38227_ (_25872_, _06854_, _06852_);
  or _38228_ (_06855_, _04605_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _38229_ (_06856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _38230_ (_06857_, _06856_, _04376_);
  or _38231_ (_06858_, _06857_, _04579_);
  nand _38232_ (_06860_, _06858_, _06855_);
  nand _38233_ (_25874_, _06860_, _02066_);
  and _38234_ (_06861_, _25618_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or _38235_ (_06862_, _26599_, _26583_);
  or _38236_ (_06863_, _06862_, _02380_);
  or _38237_ (_06865_, _06863_, _06572_);
  or _38238_ (_06867_, _04958_, _05080_);
  or _38239_ (_06868_, _04979_, _04943_);
  or _38240_ (_06870_, _06868_, _06867_);
  or _38241_ (_06871_, _05070_, _26635_);
  or _38242_ (_06872_, _06871_, _25622_);
  or _38243_ (_06873_, _06872_, _05060_);
  or _38244_ (_06874_, _06873_, _06870_);
  or _38245_ (_06875_, _06874_, _06865_);
  and _38246_ (_06876_, _06875_, _25644_);
  or _38247_ (_26872_[0], _06876_, _06861_);
  and _38248_ (_06877_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and _38249_ (_06878_, _05398_, _23824_);
  or _38250_ (_25944_, _06878_, _06877_);
  and _38251_ (_06879_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and _38252_ (_06880_, _05398_, _23898_);
  or _38253_ (_25951_, _06880_, _06879_);
  and _38254_ (_06881_, _05410_, _23707_);
  and _38255_ (_06882_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  or _38256_ (_25972_, _06882_, _06881_);
  and _38257_ (_06883_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and _38258_ (_06884_, _05398_, _23747_);
  or _38259_ (_25999_, _06884_, _06883_);
  nor _38260_ (_26897_[4], _00640_, rst);
  and _38261_ (_06886_, _23785_, _23753_);
  and _38262_ (_06888_, _06886_, _24005_);
  not _38263_ (_06889_, _06888_);
  and _38264_ (_06890_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  and _38265_ (_06892_, _06888_, _23946_);
  or _38266_ (_27014_, _06892_, _06890_);
  and _38267_ (_06894_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  and _38268_ (_06895_, _06888_, _23649_);
  or _38269_ (_26025_, _06895_, _06894_);
  and _38270_ (_06896_, _24766_, _24010_);
  not _38271_ (_06897_, _06896_);
  and _38272_ (_06898_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and _38273_ (_06899_, _06896_, _23778_);
  or _38274_ (_26050_, _06899_, _06898_);
  and _38275_ (_06900_, _24766_, _24085_);
  not _38276_ (_06902_, _06900_);
  and _38277_ (_06903_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and _38278_ (_06904_, _06900_, _23824_);
  or _38279_ (_26054_, _06904_, _06903_);
  and _38280_ (_06905_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and _38281_ (_06906_, _06900_, _23747_);
  or _38282_ (_26057_, _06906_, _06905_);
  and _38283_ (_06907_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and _38284_ (_06908_, _06900_, _23946_);
  or _38285_ (_26059_, _06908_, _06907_);
  and _38286_ (_06910_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and _38287_ (_06912_, _06900_, _24050_);
  or _38288_ (_26066_, _06912_, _06910_);
  and _38289_ (_06914_, _04811_, _23824_);
  and _38290_ (_06916_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  or _38291_ (_26068_, _06916_, _06914_);
  and _38292_ (_06918_, _06886_, _23903_);
  not _38293_ (_06919_, _06918_);
  and _38294_ (_06920_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and _38295_ (_06921_, _06918_, _24050_);
  or _38296_ (_26071_, _06921_, _06920_);
  and _38297_ (_06922_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and _38298_ (_06924_, _06918_, _23707_);
  or _38299_ (_27017_, _06924_, _06922_);
  and _38300_ (_06927_, _06886_, _23991_);
  not _38301_ (_06928_, _06927_);
  and _38302_ (_06930_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and _38303_ (_06931_, _06927_, _23898_);
  or _38304_ (_26081_, _06931_, _06930_);
  and _38305_ (_06933_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and _38306_ (_06935_, _06927_, _23824_);
  or _38307_ (_26087_, _06935_, _06933_);
  and _38308_ (_06936_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and _38309_ (_06937_, _06927_, _23946_);
  or _38310_ (_26093_, _06937_, _06936_);
  nor _38311_ (_27304_[0], \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or _38312_ (_06940_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor _38313_ (_06941_, _05727_, rst);
  and _38314_ (_27304_[1], _06941_, _06940_);
  nor _38315_ (_06942_, _05727_, _05726_);
  or _38316_ (_06943_, _06942_, _05728_);
  and _38317_ (_06944_, _05731_, _22762_);
  and _38318_ (_27304_[2], _06944_, _06943_);
  nand _38319_ (_06945_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _38320_ (_06946_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _38321_ (_06947_, _06946_, _06945_);
  nand _38322_ (_06948_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _38323_ (_06949_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _38324_ (_06950_, _06949_, _06948_);
  and _38325_ (_06951_, _06950_, _06947_);
  nand _38326_ (_06952_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand _38327_ (_06953_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _38328_ (_06954_, _06953_, _06952_);
  nand _38329_ (_06955_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand _38330_ (_06956_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _38331_ (_06957_, _06956_, _06955_);
  and _38332_ (_06958_, _06957_, _06954_);
  and _38333_ (_06959_, _06958_, _06951_);
  nand _38334_ (_06961_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand _38335_ (_06962_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _38336_ (_06963_, _06962_, _06961_);
  nand _38337_ (_06964_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand _38338_ (_06966_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _38339_ (_06967_, _06966_, _06964_);
  and _38340_ (_06968_, _06967_, _06963_);
  nand _38341_ (_06970_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  nand _38342_ (_06971_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _38343_ (_06973_, _06971_, _06970_);
  nand _38344_ (_06975_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand _38345_ (_06976_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _38346_ (_06978_, _06976_, _06975_);
  and _38347_ (_06979_, _06978_, _06973_);
  and _38348_ (_06980_, _06979_, _06968_);
  and _38349_ (_06981_, _06980_, _06959_);
  nand _38350_ (_06982_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nand _38351_ (_06983_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _38352_ (_06984_, _06983_, _06982_);
  nand _38353_ (_06985_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _38354_ (_06987_, _06421_, _00113_);
  and _38355_ (_06988_, _06987_, _06985_);
  and _38356_ (_06989_, _06988_, _06984_);
  nand _38357_ (_06990_, _06480_, _06136_);
  nand _38358_ (_06991_, _06482_, _06097_);
  and _38359_ (_06992_, _06991_, _06990_);
  nand _38360_ (_06993_, _06486_, _06207_);
  nand _38361_ (_06995_, _06488_, _06237_);
  and _38362_ (_06996_, _06995_, _06993_);
  and _38363_ (_06997_, _06996_, _06992_);
  and _38364_ (_06998_, _06997_, _06989_);
  not _38365_ (_07000_, _06351_);
  or _38366_ (_07001_, _07000_, _05860_);
  nand _38367_ (_07002_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _38368_ (_07003_, _07002_, _07001_);
  and _38369_ (_07004_, _07003_, _06998_);
  nand _38370_ (_07005_, _07004_, _06981_);
  and _38371_ (_07006_, _07005_, _06357_);
  nand _38372_ (_07007_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _38373_ (_07008_, _07007_, _06502_);
  or _38374_ (_07009_, _07008_, _07006_);
  or _38375_ (_07010_, _06502_, _26565_);
  and _38376_ (_07012_, _07010_, _22762_);
  and _38377_ (_27307_[0], _07012_, _07009_);
  and _38378_ (_07014_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _38379_ (_07015_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _38380_ (_07016_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _38381_ (_07017_, _07016_, _07015_);
  and _38382_ (_07019_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _38383_ (_07020_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _38384_ (_07021_, _07020_, _07019_);
  or _38385_ (_07023_, _07021_, _07017_);
  and _38386_ (_07024_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _38387_ (_07025_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _38388_ (_07026_, _07025_, _07024_);
  and _38389_ (_07027_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _38390_ (_07028_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _38391_ (_07029_, _07028_, _07027_);
  or _38392_ (_07030_, _07029_, _07026_);
  or _38393_ (_07031_, _07030_, _07023_);
  and _38394_ (_07032_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _38395_ (_07033_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _38396_ (_07035_, _07033_, _07032_);
  and _38397_ (_07036_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _38398_ (_07037_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _38399_ (_07038_, _07037_, _07036_);
  or _38400_ (_07039_, _07038_, _07035_);
  and _38401_ (_07040_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and _38402_ (_07041_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _38403_ (_07042_, _07041_, _07040_);
  and _38404_ (_07043_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _38405_ (_07044_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or _38406_ (_07045_, _07044_, _07043_);
  or _38407_ (_07046_, _07045_, _07042_);
  or _38408_ (_07047_, _07046_, _07039_);
  or _38409_ (_07048_, _07047_, _07031_);
  and _38410_ (_07049_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _38411_ (_07050_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _38412_ (_07051_, _07050_, _07049_);
  and _38413_ (_07052_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _38414_ (_07054_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or _38415_ (_07056_, _07054_, _07052_);
  and _38416_ (_07057_, _06421_, _00078_);
  and _38417_ (_07058_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _38418_ (_07059_, _07058_, _07057_);
  or _38419_ (_07060_, _07059_, _07056_);
  and _38420_ (_07062_, _06480_, _06125_);
  and _38421_ (_07063_, _06482_, _06092_);
  or _38422_ (_07064_, _07063_, _07062_);
  and _38423_ (_07065_, _06486_, _06202_);
  and _38424_ (_07066_, _06488_, _06232_);
  or _38425_ (_07067_, _07066_, _07065_);
  or _38426_ (_07068_, _07067_, _07064_);
  or _38427_ (_07069_, _07068_, _07060_);
  or _38428_ (_07070_, _07069_, _07051_);
  or _38429_ (_07071_, _07070_, _07048_);
  and _38430_ (_07072_, _07071_, _06357_);
  or _38431_ (_07073_, _07072_, _06361_);
  or _38432_ (_07074_, _07073_, _07014_);
  nand _38433_ (_07075_, _06361_, _00372_);
  and _38434_ (_07076_, _07075_, _22762_);
  and _38435_ (_27307_[1], _07076_, _07074_);
  and _38436_ (_07077_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _38437_ (_07078_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _38438_ (_07079_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _38439_ (_07080_, _07079_, _07078_);
  and _38440_ (_07082_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _38441_ (_07083_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _38442_ (_07084_, _07083_, _07082_);
  or _38443_ (_07085_, _07084_, _07080_);
  and _38444_ (_07087_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _38445_ (_07088_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _38446_ (_07090_, _07088_, _07087_);
  and _38447_ (_07091_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _38448_ (_07093_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _38449_ (_07094_, _07093_, _07091_);
  or _38450_ (_07095_, _07094_, _07090_);
  or _38451_ (_07096_, _07095_, _07085_);
  and _38452_ (_07097_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _38453_ (_07099_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or _38454_ (_07100_, _07099_, _07097_);
  and _38455_ (_07101_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _38456_ (_07102_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _38457_ (_07103_, _07102_, _07101_);
  or _38458_ (_07104_, _07103_, _07100_);
  and _38459_ (_07105_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and _38460_ (_07107_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _38461_ (_07108_, _07107_, _07105_);
  and _38462_ (_07109_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _38463_ (_07111_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or _38464_ (_07112_, _07111_, _07109_);
  or _38465_ (_07113_, _07112_, _07108_);
  or _38466_ (_07114_, _07113_, _07104_);
  or _38467_ (_07115_, _07114_, _07096_);
  and _38468_ (_07116_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _38469_ (_07117_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _38470_ (_07118_, _07117_, _07116_);
  and _38471_ (_07119_, _06421_, _00148_);
  and _38472_ (_07120_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _38473_ (_07121_, _07120_, _07119_);
  or _38474_ (_07122_, _07121_, _07118_);
  and _38475_ (_07123_, _06480_, _06130_);
  and _38476_ (_07124_, _06482_, _06105_);
  or _38477_ (_07125_, _07124_, _07123_);
  and _38478_ (_07126_, _06486_, _06212_);
  and _38479_ (_07127_, _06488_, _06223_);
  or _38480_ (_07128_, _07127_, _07126_);
  or _38481_ (_07129_, _07128_, _07125_);
  or _38482_ (_07130_, _07129_, _07122_);
  and _38483_ (_07131_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _38484_ (_07132_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _38485_ (_07133_, _07132_, _07131_);
  or _38486_ (_07134_, _07133_, _07130_);
  or _38487_ (_07135_, _07134_, _07115_);
  and _38488_ (_07136_, _07135_, _06357_);
  or _38489_ (_07137_, _07136_, _06361_);
  or _38490_ (_07138_, _07137_, _07077_);
  or _38491_ (_07139_, _06502_, _00451_);
  and _38492_ (_07140_, _07139_, _22762_);
  and _38493_ (_27307_[2], _07140_, _07138_);
  and _38494_ (_07141_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _38495_ (_07142_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _38496_ (_07143_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _38497_ (_07144_, _07143_, _07142_);
  and _38498_ (_07145_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _38499_ (_07146_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _38500_ (_07147_, _07146_, _07145_);
  or _38501_ (_07148_, _07147_, _07144_);
  and _38502_ (_07149_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _38503_ (_07151_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or _38504_ (_07152_, _07151_, _07149_);
  and _38505_ (_07153_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _38506_ (_07154_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _38507_ (_07155_, _07154_, _07153_);
  or _38508_ (_07156_, _07155_, _07152_);
  or _38509_ (_07157_, _07156_, _07148_);
  and _38510_ (_07158_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _38511_ (_07159_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or _38512_ (_07160_, _07159_, _07158_);
  and _38513_ (_07161_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _38514_ (_07162_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _38515_ (_07163_, _07162_, _07161_);
  or _38516_ (_07164_, _07163_, _07160_);
  and _38517_ (_07165_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and _38518_ (_07166_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _38519_ (_07167_, _07166_, _07165_);
  and _38520_ (_07168_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _38521_ (_07169_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _38522_ (_07170_, _07169_, _07168_);
  or _38523_ (_07171_, _07170_, _07167_);
  or _38524_ (_07172_, _07171_, _07164_);
  or _38525_ (_07174_, _07172_, _07157_);
  and _38526_ (_07175_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _38527_ (_07176_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or _38528_ (_07177_, _07176_, _07175_);
  and _38529_ (_07178_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _38530_ (_07179_, _06421_, _00030_);
  or _38531_ (_07180_, _07179_, _07178_);
  or _38532_ (_07181_, _07180_, _07177_);
  and _38533_ (_07182_, _06480_, _06119_);
  and _38534_ (_07183_, _06482_, _06110_);
  or _38535_ (_07184_, _07183_, _07182_);
  and _38536_ (_07186_, _06486_, _06216_);
  and _38537_ (_07187_, _06488_, _06227_);
  or _38538_ (_07188_, _07187_, _07186_);
  or _38539_ (_07189_, _07188_, _07184_);
  or _38540_ (_07190_, _07189_, _07181_);
  and _38541_ (_07192_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _38542_ (_07193_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _38543_ (_07194_, _07193_, _07192_);
  or _38544_ (_07196_, _07194_, _07190_);
  or _38545_ (_07197_, _07196_, _07174_);
  and _38546_ (_07198_, _07197_, _06357_);
  or _38547_ (_07199_, _07198_, _06361_);
  or _38548_ (_07200_, _07199_, _07141_);
  or _38549_ (_07201_, _06502_, _00545_);
  and _38550_ (_07202_, _07201_, _22762_);
  and _38551_ (_27307_[3], _07202_, _07200_);
  and _38552_ (_07204_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _38553_ (_07205_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand _38554_ (_07206_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _38555_ (_07207_, _07206_, _07205_);
  nand _38556_ (_07209_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand _38557_ (_07210_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _38558_ (_07211_, _07210_, _07209_);
  and _38559_ (_07212_, _07211_, _07207_);
  nand _38560_ (_07213_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nand _38561_ (_07214_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _38562_ (_07215_, _07214_, _07213_);
  nand _38563_ (_07216_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand _38564_ (_07217_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _38565_ (_07219_, _07217_, _07216_);
  and _38566_ (_07220_, _07219_, _07215_);
  and _38567_ (_07221_, _07220_, _07212_);
  nand _38568_ (_07223_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand _38569_ (_07224_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _38570_ (_07225_, _07224_, _07223_);
  nand _38571_ (_07227_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _38572_ (_07229_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _38573_ (_07230_, _07229_, _07227_);
  and _38574_ (_07232_, _07230_, _07225_);
  nand _38575_ (_07233_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  nand _38576_ (_07235_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _38577_ (_07236_, _07235_, _07233_);
  nand _38578_ (_07238_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  nand _38579_ (_07239_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _38580_ (_07240_, _07239_, _07238_);
  and _38581_ (_07242_, _07240_, _07236_);
  and _38582_ (_07243_, _07242_, _07232_);
  and _38583_ (_07245_, _07243_, _07221_);
  nand _38584_ (_07247_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand _38585_ (_07248_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _38586_ (_07249_, _07248_, _07247_);
  nand _38587_ (_07251_, _06421_, _00047_);
  nand _38588_ (_07252_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _38589_ (_07254_, _07252_, _07251_);
  and _38590_ (_07255_, _07254_, _07249_);
  nand _38591_ (_07256_, _06480_, _06152_);
  nand _38592_ (_07257_, _06482_, _06179_);
  and _38593_ (_07258_, _07257_, _07256_);
  nand _38594_ (_07259_, _06486_, _06278_);
  nand _38595_ (_07260_, _06488_, _06251_);
  and _38596_ (_07261_, _07260_, _07259_);
  and _38597_ (_07262_, _07261_, _07258_);
  and _38598_ (_07263_, _07262_, _07255_);
  nand _38599_ (_07264_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nand _38600_ (_07265_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _38601_ (_07266_, _07265_, _07264_);
  and _38602_ (_07267_, _07266_, _07263_);
  and _38603_ (_07268_, _07267_, _07245_);
  nor _38604_ (_07269_, _06341_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or _38605_ (_07270_, _07269_, _06355_);
  nor _38606_ (_07271_, _07270_, _07268_);
  or _38607_ (_07272_, _07271_, _06361_);
  or _38608_ (_07273_, _07272_, _07204_);
  or _38609_ (_07274_, _06502_, _00620_);
  and _38610_ (_07275_, _07274_, _22762_);
  and _38611_ (_27307_[4], _07275_, _07273_);
  and _38612_ (_07276_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _38613_ (_07277_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _38614_ (_07279_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _38615_ (_07280_, _07279_, _07277_);
  and _38616_ (_07283_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _38617_ (_07284_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _38618_ (_07285_, _07284_, _07283_);
  or _38619_ (_07286_, _07285_, _07280_);
  and _38620_ (_07288_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _38621_ (_07289_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _38622_ (_07291_, _07289_, _07288_);
  and _38623_ (_07292_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _38624_ (_07293_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _38625_ (_07294_, _07293_, _07292_);
  or _38626_ (_07295_, _07294_, _07291_);
  or _38627_ (_07296_, _07295_, _07286_);
  and _38628_ (_07297_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _38629_ (_07298_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _38630_ (_07299_, _07298_, _07297_);
  and _38631_ (_07301_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _38632_ (_07302_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _38633_ (_07303_, _07302_, _07301_);
  or _38634_ (_07304_, _07303_, _07299_);
  and _38635_ (_07306_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and _38636_ (_07307_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _38637_ (_07308_, _07307_, _07306_);
  and _38638_ (_07309_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _38639_ (_07311_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or _38640_ (_07312_, _07311_, _07309_);
  or _38641_ (_07313_, _07312_, _07308_);
  or _38642_ (_07314_, _07313_, _07304_);
  or _38643_ (_07315_, _07314_, _07296_);
  and _38644_ (_07316_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _38645_ (_07317_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or _38646_ (_07318_, _07317_, _07316_);
  and _38647_ (_07319_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _38648_ (_07320_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or _38649_ (_07321_, _07320_, _07319_);
  not _38650_ (_07322_, _26826_);
  and _38651_ (_07323_, _06421_, _07322_);
  and _38652_ (_07324_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or _38653_ (_07325_, _07324_, _07323_);
  or _38654_ (_07326_, _07325_, _07321_);
  and _38655_ (_07327_, _06480_, _06162_);
  and _38656_ (_07328_, _06482_, _06173_);
  or _38657_ (_07329_, _07328_, _07327_);
  and _38658_ (_07330_, _06486_, _06272_);
  and _38659_ (_07331_, _06488_, _06246_);
  or _38660_ (_07332_, _07331_, _07330_);
  or _38661_ (_07333_, _07332_, _07329_);
  or _38662_ (_07334_, _07333_, _07326_);
  or _38663_ (_07335_, _07334_, _07318_);
  or _38664_ (_07336_, _07335_, _07315_);
  and _38665_ (_07337_, _07336_, _06357_);
  or _38666_ (_07339_, _07337_, _06361_);
  or _38667_ (_07340_, _07339_, _07276_);
  or _38668_ (_07341_, _06502_, _00708_);
  and _38669_ (_07343_, _07341_, _22762_);
  and _38670_ (_27307_[5], _07343_, _07340_);
  and _38671_ (_07344_, _06432_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _38672_ (_07345_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand _38673_ (_07346_, _06367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _38674_ (_07347_, _07346_, _07345_);
  nand _38675_ (_07348_, _06375_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nand _38676_ (_07349_, _06377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _38677_ (_07350_, _07349_, _07348_);
  and _38678_ (_07351_, _07350_, _07347_);
  nand _38679_ (_07352_, _06389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nand _38680_ (_07353_, _06387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _38681_ (_07354_, _07353_, _07352_);
  and _38682_ (_07355_, _06381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _38683_ (_07356_, _06384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nor _38684_ (_07357_, _07356_, _07355_);
  and _38685_ (_07358_, _07357_, _07354_);
  and _38686_ (_07360_, _07358_, _07351_);
  nand _38687_ (_07361_, _06410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  nand _38688_ (_07362_, _06411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _38689_ (_07364_, _07362_, _07361_);
  nand _38690_ (_07365_, _06407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  nand _38691_ (_07366_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _38692_ (_07367_, _07366_, _07365_);
  and _38693_ (_07368_, _07367_, _07364_);
  nand _38694_ (_07369_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand _38695_ (_07370_, _06397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _38696_ (_07371_, _07370_, _07369_);
  nand _38697_ (_07372_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _38698_ (_07373_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _38699_ (_07374_, _07373_, _07372_);
  and _38700_ (_07375_, _07374_, _07371_);
  and _38701_ (_07376_, _07375_, _07368_);
  and _38702_ (_07377_, _07376_, _07360_);
  nand _38703_ (_07378_, _06346_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nand _38704_ (_07379_, _06359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _38705_ (_07380_, _07379_, _07378_);
  not _38706_ (_07381_, _26788_);
  nand _38707_ (_07382_, _06421_, _07381_);
  nand _38708_ (_07383_, _06423_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _38709_ (_07384_, _07383_, _07382_);
  and _38710_ (_07385_, _07384_, _07380_);
  nand _38711_ (_07386_, _06480_, _06146_);
  nand _38712_ (_07387_, _06482_, _06187_);
  and _38713_ (_07388_, _07387_, _07386_);
  nand _38714_ (_07389_, _06486_, _06284_);
  nand _38715_ (_07391_, _06488_, _06258_);
  and _38716_ (_07392_, _07391_, _07389_);
  and _38717_ (_07393_, _07392_, _07388_);
  and _38718_ (_07394_, _07393_, _07385_);
  nand _38719_ (_07395_, _06333_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand _38720_ (_07397_, _06351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _38721_ (_07398_, _07397_, _07395_);
  and _38722_ (_07399_, _07398_, _07394_);
  and _38723_ (_07400_, _07399_, _07377_);
  nor _38724_ (_07401_, _06341_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or _38725_ (_07403_, _07401_, _06355_);
  nor _38726_ (_07404_, _07403_, _07400_);
  or _38727_ (_07405_, _07404_, _06361_);
  or _38728_ (_07406_, _07405_, _07344_);
  nand _38729_ (_07407_, _06361_, _00793_);
  and _38730_ (_07409_, _07407_, _22762_);
  and _38731_ (_27307_[6], _07409_, _07406_);
  and _38732_ (_07410_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and _38733_ (_07411_, _06927_, _24050_);
  or _38734_ (_26132_, _07411_, _07410_);
  or _38735_ (_07412_, _04891_, _23642_);
  nand _38736_ (_07413_, _04882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _38737_ (_07414_, _04882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _38738_ (_07415_, _07414_, _26097_);
  and _38739_ (_07417_, _07415_, _07413_);
  and _38740_ (_07418_, _04864_, _24309_);
  or _38741_ (_07419_, _07418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _38742_ (_07420_, _05158_, _04864_);
  not _38743_ (_07421_, _07420_);
  and _38744_ (_07422_, _07421_, _04860_);
  and _38745_ (_07423_, _07422_, _07419_);
  and _38746_ (_07424_, _04876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _38747_ (_07426_, _07424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _38748_ (_07427_, _07424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _38749_ (_07429_, _07427_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _38750_ (_07430_, _07429_, _07426_);
  or _38751_ (_07431_, _07430_, _07423_);
  or _38752_ (_07432_, _07431_, _07417_);
  or _38753_ (_07433_, _07432_, _24299_);
  and _38754_ (_07434_, _07433_, _24294_);
  and _38755_ (_07436_, _07434_, _07412_);
  and _38756_ (_07437_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _38757_ (_07438_, _07437_, _07436_);
  and _38758_ (_26617_, _07438_, _22762_);
  and _38759_ (_07439_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  and _38760_ (_07440_, _02298_, _23747_);
  or _38761_ (_26642_, _07440_, _07439_);
  and _38762_ (_07442_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  and _38763_ (_07443_, _02298_, _23649_);
  or _38764_ (_26649_, _07443_, _07442_);
  and _38765_ (_07444_, _04917_, _23778_);
  and _38766_ (_07446_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or _38767_ (_26664_, _07446_, _07444_);
  and _38768_ (_07447_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  and _38769_ (_07448_, _02298_, _23946_);
  or _38770_ (_26667_, _07448_, _07447_);
  or _38771_ (_07449_, _04891_, _23939_);
  not _38772_ (_07450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _38773_ (_07451_, _07420_, _26099_);
  nor _38774_ (_07452_, _07451_, _07450_);
  and _38775_ (_07454_, _07451_, _07450_);
  or _38776_ (_07455_, _07454_, _07452_);
  and _38777_ (_07456_, _07455_, _04861_);
  and _38778_ (_07457_, _05158_, _24300_);
  or _38779_ (_07458_, _07457_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _38780_ (_07459_, _07458_, _24302_);
  nor _38781_ (_07460_, _07459_, _05151_);
  or _38782_ (_07461_, _05164_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _38783_ (_07462_, _05165_, _26098_);
  and _38784_ (_07463_, _07462_, _07461_);
  or _38785_ (_07464_, _07463_, _07460_);
  or _38786_ (_07465_, _07464_, _07456_);
  or _38787_ (_07466_, _07465_, _24299_);
  and _38788_ (_07467_, _07466_, _24294_);
  and _38789_ (_07468_, _07467_, _07449_);
  and _38790_ (_07469_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _38791_ (_07470_, _07469_, _07468_);
  and _38792_ (_26690_, _07470_, _22762_);
  and _38793_ (_07471_, _01809_, _24010_);
  and _38794_ (_07472_, _07471_, _23946_);
  not _38795_ (_07473_, _07471_);
  and _38796_ (_07474_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  or _38797_ (_27107_, _07474_, _07472_);
  and _38798_ (_07475_, _04811_, _23707_);
  and _38799_ (_07476_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or _38800_ (_26706_, _07476_, _07475_);
  and _38801_ (_07477_, _07471_, _23649_);
  and _38802_ (_07478_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  or _38803_ (_26720_, _07478_, _07477_);
  and _38804_ (_07479_, _07471_, _23824_);
  and _38805_ (_07480_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  or _38806_ (_26726_, _07480_, _07479_);
  and _38807_ (_07482_, _07471_, _23778_);
  and _38808_ (_07483_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  or _38809_ (_26731_, _07483_, _07482_);
  and _38810_ (_07484_, _05445_, _24050_);
  and _38811_ (_07486_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  or _38812_ (_26748_, _07486_, _07484_);
  and _38813_ (_07488_, _05445_, _23946_);
  and _38814_ (_07489_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  or _38815_ (_26764_, _07489_, _07488_);
  and _38816_ (_07492_, _24329_, _24201_);
  not _38817_ (_07493_, _07492_);
  and _38818_ (_07494_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and _38819_ (_07496_, _07492_, _24050_);
  or _38820_ (_26769_, _07496_, _07494_);
  and _38821_ (_07497_, _25142_, _23649_);
  and _38822_ (_07499_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  or _38823_ (_26771_, _07499_, _07497_);
  and _38824_ (_07500_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _38825_ (_07501_, _24128_, _24043_);
  not _38826_ (_07502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _38827_ (_07503_, _25684_, _07502_);
  and _38828_ (_07504_, _25684_, _07502_);
  or _38829_ (_07505_, _07504_, _07503_);
  or _38830_ (_07506_, _07505_, _24127_);
  and _38831_ (_07508_, _07506_, _24166_);
  and _38832_ (_07509_, _07508_, _07501_);
  or _38833_ (_26774_, _07509_, _07500_);
  and _38834_ (_07510_, _25733_, _23824_);
  and _38835_ (_07511_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or _38836_ (_26780_, _07511_, _07510_);
  and _38837_ (_26860_[1], _23866_, _22762_);
  and _38838_ (_07513_, _04760_, _23069_);
  not _38839_ (_07514_, _07513_);
  and _38840_ (_07515_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and _38841_ (_07516_, _07513_, _23898_);
  or _38842_ (_26963_, _07516_, _07515_);
  and _38843_ (_26860_[2], _24436_, _22762_);
  and _38844_ (_07517_, _05445_, _23747_);
  and _38845_ (_07518_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  or _38846_ (_26805_, _07518_, _07517_);
  and _38847_ (_07519_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  and _38848_ (_07521_, _07492_, _23946_);
  or _38849_ (_26828_, _07521_, _07519_);
  and _38850_ (_07522_, _05445_, _23898_);
  and _38851_ (_07524_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  or _38852_ (_26834_, _07524_, _07522_);
  and _38853_ (_07525_, _06886_, _24275_);
  not _38854_ (_07526_, _07525_);
  and _38855_ (_07527_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  and _38856_ (_07530_, _07525_, _23778_);
  or _38857_ (_00090_, _07530_, _07527_);
  and _38858_ (_26910_, _02443_, _22762_);
  and _38859_ (_26911_[7], _23706_, _22762_);
  nor _38860_ (_26913_[2], _00168_, rst);
  and _38861_ (_07533_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  and _38862_ (_07534_, _07525_, _23898_);
  or _38863_ (_00200_, _07534_, _07533_);
  and _38864_ (_07536_, _01809_, _25078_);
  and _38865_ (_07537_, _07536_, _23778_);
  not _38866_ (_07539_, _07536_);
  and _38867_ (_07541_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  or _38868_ (_00203_, _07541_, _07537_);
  and _38869_ (_07542_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  and _38870_ (_07543_, _07525_, _23649_);
  or _38871_ (_00206_, _07543_, _07542_);
  and _38872_ (_07544_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  and _38873_ (_07545_, _07525_, _23946_);
  or _38874_ (_00269_, _07545_, _07544_);
  and _38875_ (_07547_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  and _38876_ (_07550_, _07525_, _23707_);
  or _38877_ (_00275_, _07550_, _07547_);
  and _38878_ (_07551_, _24766_, _23784_);
  not _38879_ (_07552_, _07551_);
  and _38880_ (_07553_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  and _38881_ (_07554_, _07551_, _23778_);
  or _38882_ (_00279_, _07554_, _07553_);
  nor _38883_ (_26887_[2], _00163_, rst);
  and _38884_ (_07555_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  and _38885_ (_07556_, _07551_, _23824_);
  or _38886_ (_00296_, _07556_, _07555_);
  and _38887_ (_07557_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  and _38888_ (_07558_, _07551_, _23649_);
  or _38889_ (_00299_, _07558_, _07557_);
  and _38890_ (_07559_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  and _38891_ (_07560_, _07551_, _24050_);
  or _38892_ (_00309_, _07560_, _07559_);
  and _38893_ (_26911_[0], _23777_, _22762_);
  and _38894_ (_26911_[1], _23897_, _22762_);
  and _38895_ (_26911_[2], _23823_, _22762_);
  and _38896_ (_26911_[3], _23746_, _22762_);
  and _38897_ (_26911_[4], _23648_, _22762_);
  and _38898_ (_26911_[5], _23945_, _22762_);
  and _38899_ (_26911_[6], _24049_, _22762_);
  and _38900_ (_07562_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  and _38901_ (_07563_, _07551_, _23707_);
  or _38902_ (_00385_, _07563_, _07562_);
  nor _38903_ (_26913_[0], _00134_, rst);
  nor _38904_ (_26913_[1], _00099_, rst);
  nor _38905_ (_07566_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _38906_ (_07568_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _23978_);
  nor _38907_ (_07570_, _07568_, _07566_);
  not _38908_ (_07572_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _38909_ (_07574_, _00587_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _38910_ (_07576_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _23978_);
  nor _38911_ (_07577_, _07576_, _07574_);
  and _38912_ (_07578_, _07577_, _07572_);
  nor _38913_ (_07580_, _07577_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _38914_ (_07581_, _07580_, _07578_);
  not _38915_ (_07582_, _07581_);
  nor _38916_ (_07583_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _38917_ (_07584_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _23978_);
  nor _38918_ (_07585_, _07584_, _07583_);
  not _38919_ (_07586_, _07585_);
  nor _38920_ (_07588_, _00495_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _38921_ (_07589_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _23978_);
  nor _38922_ (_07590_, _07589_, _07588_);
  and _38923_ (_07591_, _07590_, _07586_);
  nand _38924_ (_07592_, _07591_, _07582_);
  and _38925_ (_07594_, _07592_, _07570_);
  nor _38926_ (_07597_, _07590_, _07586_);
  not _38927_ (_07599_, _07597_);
  not _38928_ (_07600_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _38929_ (_07601_, _07577_, _07600_);
  and _38930_ (_07603_, _07577_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _38931_ (_07605_, _07603_, _07601_);
  nor _38932_ (_07606_, _07605_, _07599_);
  and _38933_ (_07608_, _07590_, _07585_);
  not _38934_ (_07610_, _07608_);
  not _38935_ (_07612_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _38936_ (_07613_, _07577_, _07612_);
  nor _38937_ (_07615_, _07577_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _38938_ (_07616_, _07615_, _07613_);
  nor _38939_ (_07618_, _07616_, _07610_);
  nor _38940_ (_07619_, _07618_, _07606_);
  not _38941_ (_07621_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _38942_ (_07623_, _07577_, _07621_);
  nor _38943_ (_07624_, _07590_, _07585_);
  not _38944_ (_07626_, _07624_);
  nor _38945_ (_07628_, _07577_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _38946_ (_07631_, _07628_, _07626_);
  or _38947_ (_07632_, _07631_, _07623_);
  and _38948_ (_07634_, _07632_, _07619_);
  and _38949_ (_07636_, _07634_, _07594_);
  not _38950_ (_07637_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _38951_ (_07639_, _07577_, _07637_);
  nor _38952_ (_07641_, _07577_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _38953_ (_07642_, _07641_, _07639_);
  nor _38954_ (_07643_, _07642_, _07610_);
  nor _38955_ (_07645_, _07643_, _07570_);
  and _38956_ (_07647_, _07577_, \oc8051_symbolic_cxrom1.regvalid [12]);
  not _38957_ (_07648_, _07577_);
  and _38958_ (_07649_, _07648_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _38959_ (_07650_, _07649_, _07647_);
  not _38960_ (_07652_, _07650_);
  nand _38961_ (_07653_, _07652_, _07591_);
  and _38962_ (_07655_, _07577_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not _38963_ (_07657_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _38964_ (_07659_, _07577_, _07657_);
  nor _38965_ (_07660_, _07659_, _07655_);
  nor _38966_ (_07662_, _07660_, _07599_);
  nor _38967_ (_07663_, _07577_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not _38968_ (_07664_, _07663_);
  not _38969_ (_07665_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _38970_ (_07666_, _07577_, _07665_);
  nor _38971_ (_07667_, _07666_, _07626_);
  and _38972_ (_07668_, _07667_, _07664_);
  nor _38973_ (_07669_, _07668_, _07662_);
  and _38974_ (_07670_, _07669_, _07653_);
  and _38975_ (_07671_, _07670_, _07645_);
  nor _38976_ (_07672_, _07671_, _07636_);
  not _38977_ (_07673_, _07672_);
  and _38978_ (_07674_, _07673_, word_in[7]);
  not _38979_ (_07675_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand _38980_ (_07676_, _07570_, _07675_);
  or _38981_ (_07677_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _38982_ (_07678_, _07677_, _07676_);
  and _38983_ (_07679_, _07678_, _07624_);
  or _38984_ (_07681_, _07679_, _07577_);
  not _38985_ (_07682_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _38986_ (_07684_, _07570_, _07682_);
  or _38987_ (_07685_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _38988_ (_07686_, _07685_, _07684_);
  and _38989_ (_07687_, _07686_, _07608_);
  not _38990_ (_07689_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand _38991_ (_07691_, _07570_, _07689_);
  or _38992_ (_07692_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _38993_ (_07693_, _07692_, _07691_);
  and _38994_ (_07695_, _07693_, _07591_);
  not _38995_ (_07696_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _38996_ (_07698_, _07570_, _07696_);
  or _38997_ (_07700_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _38998_ (_07701_, _07700_, _07698_);
  and _38999_ (_07703_, _07701_, _07597_);
  or _39000_ (_07704_, _07703_, _07695_);
  or _39001_ (_07706_, _07704_, _07687_);
  or _39002_ (_07707_, _07706_, _07681_);
  not _39003_ (_07709_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _39004_ (_07710_, _07570_, _07709_);
  or _39005_ (_07711_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _39006_ (_07713_, _07711_, _07710_);
  and _39007_ (_07714_, _07713_, _07624_);
  or _39008_ (_07715_, _07714_, _07648_);
  not _39009_ (_07717_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _39010_ (_07718_, _07570_, _07717_);
  or _39011_ (_07720_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _39012_ (_07721_, _07720_, _07718_);
  and _39013_ (_07722_, _07721_, _07591_);
  not _39014_ (_07723_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _39015_ (_07725_, _07570_, _07723_);
  or _39016_ (_07726_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _39017_ (_07727_, _07726_, _07725_);
  and _39018_ (_07728_, _07727_, _07608_);
  or _39019_ (_07730_, _07728_, _07722_);
  not _39020_ (_07731_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _39021_ (_07732_, _07570_, _07731_);
  or _39022_ (_07733_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _39023_ (_07734_, _07733_, _07732_);
  and _39024_ (_07735_, _07734_, _07597_);
  or _39025_ (_07736_, _07735_, _07730_);
  or _39026_ (_07738_, _07736_, _07715_);
  and _39027_ (_07740_, _07738_, _07707_);
  and _39028_ (_07742_, _07740_, _07672_);
  or _39029_ (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _07742_, _07674_);
  and _39030_ (_07743_, _24085_, _23664_);
  and _39031_ (_07745_, _07743_, _23898_);
  not _39032_ (_07747_, _07743_);
  and _39033_ (_07748_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  or _39034_ (_27072_, _07748_, _07745_);
  not _39035_ (_07749_, _07570_);
  and _39036_ (_07751_, _07585_, _07749_);
  not _39037_ (_07753_, _07751_);
  and _39038_ (_07754_, _07585_, _07570_);
  and _39039_ (_07755_, _07754_, _07590_);
  nor _39040_ (_07756_, _07754_, _07590_);
  nor _39041_ (_07757_, _07756_, _07755_);
  not _39042_ (_07758_, _07757_);
  nor _39043_ (_07759_, _07758_, _07616_);
  nor _39044_ (_07760_, _07755_, _07648_);
  not _39045_ (_07761_, _07590_);
  nor _39046_ (_07762_, _07761_, _07577_);
  and _39047_ (_07763_, _07754_, _07762_);
  nor _39048_ (_07764_, _07763_, _07760_);
  and _39049_ (_07766_, _07764_, _07758_);
  and _39050_ (_07768_, _07766_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _39051_ (_07770_, _07764_, _07757_);
  and _39052_ (_07772_, _07770_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _39053_ (_07774_, _07772_, _07768_);
  nor _39054_ (_07776_, _07774_, _07759_);
  nor _39055_ (_07778_, _07776_, _07753_);
  nor _39056_ (_07780_, _07585_, _07570_);
  not _39057_ (_07782_, _07780_);
  nor _39058_ (_07783_, _07758_, _07581_);
  and _39059_ (_07784_, _07766_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _39060_ (_07785_, _07770_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _39061_ (_07786_, _07785_, _07784_);
  nor _39062_ (_07787_, _07786_, _07783_);
  nor _39063_ (_07788_, _07787_, _07782_);
  nor _39064_ (_07789_, _07788_, _07778_);
  and _39065_ (_07790_, _07586_, _07570_);
  not _39066_ (_07791_, _07790_);
  nor _39067_ (_07792_, _07758_, _07642_);
  and _39068_ (_07793_, _07766_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _39069_ (_07794_, _07770_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _39070_ (_07795_, _07794_, _07793_);
  nor _39071_ (_07796_, _07795_, _07792_);
  nor _39072_ (_07798_, _07796_, _07791_);
  not _39073_ (_07799_, _07754_);
  nor _39074_ (_07801_, _07758_, _07650_);
  and _39075_ (_07803_, _07766_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _39076_ (_07804_, _07770_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _39077_ (_07806_, _07804_, _07803_);
  nor _39078_ (_07807_, _07806_, _07801_);
  nor _39079_ (_07808_, _07807_, _07799_);
  nor _39080_ (_07809_, _07808_, _07798_);
  and _39081_ (_07810_, _07809_, _07789_);
  or _39082_ (_07811_, _07780_, _07754_);
  not _39083_ (_07812_, _07811_);
  not _39084_ (_07813_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _39085_ (_07814_, _07570_, _07813_);
  or _39086_ (_07815_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _39087_ (_07816_, _07815_, _07814_);
  and _39088_ (_07817_, _07816_, _07812_);
  not _39089_ (_07819_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _39090_ (_07821_, _07570_, _07819_);
  or _39091_ (_07822_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _39092_ (_07824_, _07822_, _07821_);
  and _39093_ (_07825_, _07824_, _07811_);
  or _39094_ (_07826_, _07825_, _07817_);
  and _39095_ (_07827_, _07826_, _07770_);
  not _39096_ (_07829_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand _39097_ (_07831_, _07570_, _07829_);
  or _39098_ (_07833_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _39099_ (_07835_, _07833_, _07831_);
  and _39100_ (_07836_, _07835_, _07812_);
  not _39101_ (_07837_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand _39102_ (_07839_, _07570_, _07837_);
  or _39103_ (_07840_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _39104_ (_07841_, _07840_, _07839_);
  and _39105_ (_07842_, _07841_, _07811_);
  or _39106_ (_07843_, _07842_, _07836_);
  and _39107_ (_07844_, _07843_, _07766_);
  and _39108_ (_07845_, _07757_, _07648_);
  not _39109_ (_07846_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand _39110_ (_07847_, _07570_, _07846_);
  or _39111_ (_07848_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _39112_ (_07849_, _07848_, _07847_);
  and _39113_ (_07850_, _07849_, _07812_);
  not _39114_ (_07852_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand _39115_ (_07853_, _07570_, _07852_);
  or _39116_ (_07855_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _39117_ (_07856_, _07855_, _07853_);
  and _39118_ (_07857_, _07856_, _07811_);
  or _39119_ (_07858_, _07857_, _07850_);
  and _39120_ (_07859_, _07858_, _07845_);
  and _39121_ (_07860_, _07757_, _07577_);
  not _39122_ (_07861_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _39123_ (_07862_, _07570_, _07861_);
  or _39124_ (_07863_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _39125_ (_07864_, _07863_, _07862_);
  and _39126_ (_07865_, _07864_, _07812_);
  not _39127_ (_07866_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _39128_ (_07867_, _07570_, _07866_);
  or _39129_ (_07868_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _39130_ (_07869_, _07868_, _07867_);
  and _39131_ (_07870_, _07869_, _07811_);
  or _39132_ (_07871_, _07870_, _07865_);
  and _39133_ (_07872_, _07871_, _07860_);
  or _39134_ (_07873_, _07872_, _07859_);
  or _39135_ (_07874_, _07873_, _07844_);
  nor _39136_ (_07875_, _07874_, _07827_);
  nor _39137_ (_07876_, _07875_, _07810_);
  and _39138_ (_07877_, _07810_, word_in[15]);
  or _39139_ (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _07877_, _07876_);
  nor _39140_ (_07878_, _07608_, _07624_);
  and _39141_ (_07879_, _07608_, _07577_);
  nor _39142_ (_07880_, _07608_, _07577_);
  nor _39143_ (_07881_, _07880_, _07879_);
  nor _39144_ (_07882_, _07881_, _07878_);
  and _39145_ (_07883_, _07882_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not _39146_ (_07884_, _07883_);
  not _39147_ (_07885_, _07878_);
  nor _39148_ (_07886_, _07885_, _07581_);
  and _39149_ (_07887_, _07881_, _07885_);
  and _39150_ (_07888_, _07887_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _39151_ (_07889_, _07888_, _07886_);
  and _39152_ (_07890_, _07889_, _07884_);
  nor _39153_ (_07891_, _07890_, _07799_);
  nor _39154_ (_07892_, _07885_, _07616_);
  and _39155_ (_07893_, _07887_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _39156_ (_07895_, _07882_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or _39157_ (_07896_, _07895_, _07893_);
  nor _39158_ (_07897_, _07896_, _07892_);
  nor _39159_ (_07898_, _07897_, _07791_);
  nor _39160_ (_07899_, _07898_, _07891_);
  nor _39161_ (_07900_, _07885_, _07642_);
  and _39162_ (_07901_, _07882_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _39163_ (_07902_, _07887_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _39164_ (_07903_, _07902_, _07901_);
  nor _39165_ (_07904_, _07903_, _07900_);
  nor _39166_ (_07905_, _07904_, _07782_);
  and _39167_ (_07906_, _07882_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not _39168_ (_07907_, _07906_);
  nor _39169_ (_07908_, _07885_, _07650_);
  and _39170_ (_07909_, _07887_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _39171_ (_07910_, _07909_, _07908_);
  and _39172_ (_07911_, _07910_, _07907_);
  nor _39173_ (_07912_, _07911_, _07753_);
  nor _39174_ (_07913_, _07912_, _07905_);
  and _39175_ (_07914_, _07913_, _07899_);
  not _39176_ (_07915_, _07881_);
  and _39177_ (_07916_, _07686_, _07591_);
  and _39178_ (_07917_, _07678_, _07577_);
  or _39179_ (_07918_, _07917_, _07916_);
  and _39180_ (_07919_, _07693_, _07597_);
  and _39181_ (_07920_, _07701_, _07624_);
  or _39182_ (_07921_, _07920_, _07919_);
  or _39183_ (_07922_, _07921_, _07918_);
  and _39184_ (_07923_, _07922_, _07915_);
  and _39185_ (_07924_, _07721_, _07597_);
  and _39186_ (_07926_, _07734_, _07624_);
  or _39187_ (_07927_, _07926_, _07924_);
  and _39188_ (_07928_, _07727_, _07591_);
  and _39189_ (_07929_, _07713_, _07608_);
  or _39190_ (_07930_, _07929_, _07928_);
  or _39191_ (_07931_, _07930_, _07927_);
  and _39192_ (_07932_, _07931_, _07881_);
  nor _39193_ (_07933_, _07932_, _07923_);
  nor _39194_ (_07934_, _07933_, _07914_);
  and _39195_ (_07935_, _07914_, word_in[23]);
  or _39196_ (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _07935_, _07934_);
  and _39197_ (_07936_, _05281_, _23824_);
  and _39198_ (_07937_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or _39199_ (_00562_, _07937_, _07936_);
  nor _39200_ (_07938_, _07782_, _07590_);
  and _39201_ (_07939_, _07938_, _07601_);
  not _39202_ (_07940_, _07938_);
  nand _39203_ (_07941_, _07782_, _07590_);
  and _39204_ (_07942_, _07941_, _07940_);
  not _39205_ (_07943_, _07942_);
  nor _39206_ (_07945_, _07943_, _07581_);
  nor _39207_ (_07946_, _07941_, _07577_);
  and _39208_ (_07947_, _07941_, _07577_);
  nor _39209_ (_07948_, _07947_, _07946_);
  and _39210_ (_07949_, _07948_, _07943_);
  and _39211_ (_07950_, _07949_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _39212_ (_07951_, _07948_, _07942_);
  and _39213_ (_07952_, _07951_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _39214_ (_07953_, _07952_, _07950_);
  nor _39215_ (_07954_, _07953_, _07945_);
  nor _39216_ (_07955_, _07954_, _07753_);
  nor _39217_ (_07956_, _07955_, _07939_);
  nor _39218_ (_07957_, _07943_, _07616_);
  and _39219_ (_07958_, _07951_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _39220_ (_07959_, _07958_, _07957_);
  nor _39221_ (_07960_, _07959_, _07782_);
  nor _39222_ (_07961_, _07943_, _07642_);
  and _39223_ (_07962_, _07949_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _39224_ (_07963_, _07951_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _39225_ (_07964_, _07963_, _07962_);
  nor _39226_ (_07965_, _07964_, _07961_);
  nor _39227_ (_07966_, _07965_, _07799_);
  nor _39228_ (_07967_, _07943_, _07650_);
  and _39229_ (_07968_, _07949_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _39230_ (_07969_, _07951_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _39231_ (_07970_, _07969_, _07968_);
  nor _39232_ (_07971_, _07970_, _07967_);
  nor _39233_ (_07972_, _07971_, _07791_);
  or _39234_ (_07973_, _07972_, _07966_);
  nor _39235_ (_07974_, _07973_, _07960_);
  and _39236_ (_07975_, _07974_, _07956_);
  and _39237_ (_07976_, _07824_, _07812_);
  and _39238_ (_07977_, _07816_, _07811_);
  or _39239_ (_07978_, _07977_, _07976_);
  and _39240_ (_07979_, _07978_, _07951_);
  and _39241_ (_07980_, _07841_, _07812_);
  and _39242_ (_07981_, _07835_, _07811_);
  or _39243_ (_07982_, _07981_, _07980_);
  and _39244_ (_07983_, _07982_, _07949_);
  and _39245_ (_07984_, _07942_, _07648_);
  and _39246_ (_07985_, _07856_, _07812_);
  and _39247_ (_07986_, _07849_, _07811_);
  or _39248_ (_07987_, _07986_, _07985_);
  and _39249_ (_07988_, _07987_, _07984_);
  and _39250_ (_07989_, _07869_, _07812_);
  and _39251_ (_07990_, _07864_, _07811_);
  or _39252_ (_07991_, _07990_, _07989_);
  and _39253_ (_07992_, _07947_, _07940_);
  and _39254_ (_07993_, _07992_, _07991_);
  or _39255_ (_07994_, _07993_, _07988_);
  or _39256_ (_07996_, _07994_, _07983_);
  nor _39257_ (_07997_, _07996_, _07979_);
  nor _39258_ (_07998_, _07997_, _07975_);
  and _39259_ (_07999_, _07975_, word_in[31]);
  or _39260_ (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _07999_, _07998_);
  and _39261_ (_08000_, _07590_, _07577_);
  or _39262_ (_08001_, _08000_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _39263_ (_26842_[15], _08001_, _22762_);
  and _39264_ (_08002_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and _39265_ (_08003_, _06896_, _23824_);
  or _39266_ (_00617_, _08003_, _08002_);
  and _39267_ (_08004_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and _39268_ (_08005_, _06896_, _23649_);
  or _39269_ (_00626_, _08005_, _08004_);
  and _39270_ (_08006_, _07914_, _22762_);
  and _39271_ (_08007_, _08006_, _07878_);
  and _39272_ (_08008_, _08007_, _07881_);
  and _39273_ (_08009_, _08008_, _07790_);
  and _39274_ (_08010_, _07810_, _22762_);
  and _39275_ (_08011_, _08010_, _07751_);
  and _39276_ (_08012_, _08011_, _07860_);
  and _39277_ (_08013_, _07636_, _22762_);
  and _39278_ (_08014_, _08013_, _07585_);
  nor _39279_ (_08015_, _07672_, rst);
  and _39280_ (_08016_, _08015_, _08000_);
  and _39281_ (_08017_, _08016_, _08014_);
  nor _39282_ (_08018_, _08017_, _07723_);
  and _39283_ (_08019_, _08015_, word_in[7]);
  and _39284_ (_08020_, _08019_, _08017_);
  or _39285_ (_08021_, _08020_, _08018_);
  or _39286_ (_08022_, _08021_, _08012_);
  not _39287_ (_08023_, _08012_);
  or _39288_ (_08024_, _08023_, word_in[15]);
  and _39289_ (_08025_, _08024_, _08022_);
  or _39290_ (_08026_, _08025_, _08009_);
  and _39291_ (_08027_, _08000_, _07780_);
  and _39292_ (_08028_, _07975_, _22762_);
  and _39293_ (_08029_, _08028_, _08027_);
  not _39294_ (_08030_, _08029_);
  not _39295_ (_08031_, _08009_);
  and _39296_ (_08033_, _08006_, word_in[23]);
  or _39297_ (_08034_, _08033_, _08031_);
  and _39298_ (_08035_, _08034_, _08030_);
  and _39299_ (_08036_, _08035_, _08026_);
  and _39300_ (_08037_, _08029_, word_in[31]);
  or _39301_ (_26849_[7], _08037_, _08036_);
  or _39302_ (_08038_, _07949_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _39303_ (_26859_, _08038_, _22762_);
  not _39304_ (_08039_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _39305_ (_08040_, _07626_, _07577_);
  nand _39306_ (_08041_, _08040_, _08039_);
  or _39307_ (_08042_, _08041_, _07879_);
  and _39308_ (_26842_[1], _08042_, _22762_);
  and _39309_ (_08043_, _24329_, _23076_);
  and _39310_ (_08044_, _08043_, _24050_);
  not _39311_ (_08045_, _08043_);
  and _39312_ (_08046_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or _39313_ (_27212_, _08046_, _08044_);
  and _39314_ (_08047_, _05410_, _23778_);
  and _39315_ (_08048_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  or _39316_ (_27213_, _08048_, _08047_);
  and _39317_ (_08050_, _07755_, _07577_);
  not _39318_ (_08051_, _08040_);
  nor _39319_ (_08052_, _08051_, _08050_);
  and _39320_ (_08053_, _07984_, _07751_);
  nor _39321_ (_08054_, _08053_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand _39322_ (_08055_, _08054_, _08052_);
  and _39323_ (_26842_[2], _08055_, _22762_);
  not _39324_ (_08056_, _07766_);
  and _39325_ (_08057_, _07984_, _07754_);
  or _39326_ (_08058_, _07590_, _07577_);
  or _39327_ (_08059_, _08058_, _07751_);
  and _39328_ (_08060_, _08059_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or _39329_ (_08061_, _08060_, _08057_);
  and _39330_ (_08062_, _08061_, _08056_);
  and _39331_ (_08063_, _07601_, _07624_);
  or _39332_ (_08064_, _08063_, _08053_);
  or _39333_ (_08065_, _08064_, _08062_);
  and _39334_ (_08066_, _08065_, _08052_);
  or _39335_ (_08067_, _08063_, _08061_);
  and _39336_ (_08068_, _08067_, _08050_);
  or _39337_ (_08069_, _08068_, _08051_);
  or _39338_ (_08070_, _08069_, _08066_);
  and _39339_ (_26842_[3], _08070_, _22762_);
  and _39340_ (_08071_, _08043_, _23707_);
  and _39341_ (_08072_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or _39342_ (_00764_, _08072_, _08071_);
  and _39343_ (_08073_, _07780_, _07762_);
  or _39344_ (_08074_, _08073_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _39345_ (_08075_, _08074_, _08058_);
  or _39346_ (_08076_, _08075_, _08057_);
  and _39347_ (_08077_, _08076_, _08056_);
  and _39348_ (_08078_, _08074_, _08050_);
  and _39349_ (_08079_, _07790_, _07984_);
  and _39350_ (_08080_, _07938_, _07648_);
  and _39351_ (_08081_, _08080_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _39352_ (_08082_, _08081_, _08079_);
  or _39353_ (_08083_, _08082_, _08078_);
  or _39354_ (_08084_, _08083_, _08053_);
  or _39355_ (_08085_, _08084_, _08077_);
  and _39356_ (_26842_[4], _08085_, _22762_);
  and _39357_ (_08087_, _02200_, _23824_);
  and _39358_ (_08088_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or _39359_ (_00828_, _08088_, _08087_);
  and _39360_ (_08091_, _02321_, _23898_);
  and _39361_ (_08093_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  or _39362_ (_27138_, _08093_, _08091_);
  or _39363_ (_08095_, _07760_, _07946_);
  or _39364_ (_08096_, _08095_, _08050_);
  not _39365_ (_08097_, _07880_);
  or _39366_ (_08098_, _08073_, _08057_);
  or _39367_ (_08099_, _08098_, _08097_);
  and _39368_ (_08101_, _08099_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _39369_ (_08102_, _08053_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _39370_ (_08104_, _07790_, _07762_);
  and _39371_ (_08105_, _08051_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _39372_ (_08106_, _08105_, _08104_);
  or _39373_ (_08108_, _08106_, _08102_);
  or _39374_ (_08109_, _08108_, _08101_);
  and _39375_ (_08111_, _08109_, _08096_);
  or _39376_ (_08112_, _08105_, _08053_);
  or _39377_ (_08113_, _08112_, _08098_);
  or _39378_ (_08114_, _08113_, _08111_);
  and _39379_ (_26842_[5], _08114_, _22762_);
  and _39380_ (_08116_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  and _39381_ (_08117_, _05199_, _23824_);
  or _39382_ (_00874_, _08117_, _08116_);
  and _39383_ (_08119_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  and _39384_ (_08120_, _05199_, _23649_);
  or _39385_ (_00921_, _08120_, _08119_);
  nor _39386_ (_08121_, _07880_, _08050_);
  and _39387_ (_08122_, _07751_, _07762_);
  or _39388_ (_08123_, _08122_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _39389_ (_08124_, _08123_, _08121_);
  and _39390_ (_08125_, _08098_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _39391_ (_08126_, _08125_, _08104_);
  or _39392_ (_08127_, _08126_, _08124_);
  and _39393_ (_08128_, _08127_, _08095_);
  and _39394_ (_08129_, _08123_, _08050_);
  and _39395_ (_08130_, _08053_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _39396_ (_08132_, _08051_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _39397_ (_08133_, _08132_, _08057_);
  or _39398_ (_08134_, _08133_, _08073_);
  or _39399_ (_08135_, _08134_, _08130_);
  or _39400_ (_08136_, _08135_, _08129_);
  or _39401_ (_08137_, _08136_, _08128_);
  and _39402_ (_26842_[6], _08137_, _22762_);
  not _39403_ (_08138_, _07764_);
  and _39404_ (_08139_, _08080_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _39405_ (_08140_, _07984_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _39406_ (_08141_, _08140_, _07782_);
  or _39407_ (_08142_, _08141_, _08139_);
  or _39408_ (_08143_, _08122_, _07577_);
  and _39409_ (_08144_, _08143_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not _39410_ (_08145_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _39411_ (_08146_, _07585_, _08145_);
  and _39412_ (_08147_, _08146_, _07762_);
  or _39413_ (_08148_, _08147_, _07763_);
  or _39414_ (_08149_, _08148_, _08144_);
  or _39415_ (_08150_, _08149_, _08142_);
  and _39416_ (_08151_, _08150_, _08138_);
  and _39417_ (_08152_, _08140_, _07570_);
  and _39418_ (_08153_, _08053_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _39419_ (_08154_, _08147_, _08122_);
  or _39420_ (_08155_, _08154_, _08153_);
  or _39421_ (_08156_, _08155_, _08152_);
  or _39422_ (_08157_, _08156_, _08151_);
  and _39423_ (_08158_, _08157_, _08121_);
  and _39424_ (_08159_, _08150_, _08050_);
  or _39425_ (_08160_, _08139_, _08073_);
  or _39426_ (_08163_, _08160_, _08104_);
  or _39427_ (_08164_, _08163_, _08140_);
  or _39428_ (_08165_, _08164_, _08159_);
  or _39429_ (_08166_, _08165_, _08158_);
  and _39430_ (_26842_[7], _08166_, _22762_);
  and _39431_ (_08167_, _01809_, _24005_);
  and _39432_ (_08168_, _08167_, _23946_);
  not _39433_ (_08169_, _08167_);
  and _39434_ (_08171_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or _39435_ (_00995_, _08171_, _08168_);
  and _39436_ (_08173_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  and _39437_ (_08174_, _05199_, _23747_);
  or _39438_ (_01020_, _08174_, _08173_);
  not _39439_ (_08176_, _08058_);
  nor _39440_ (_08177_, _07984_, _07951_);
  and _39441_ (_08178_, _08177_, _07577_);
  or _39442_ (_08180_, _08178_, _08176_);
  and _39443_ (_08182_, _08180_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _39444_ (_08184_, _07938_, _07577_);
  and _39445_ (_08185_, _07762_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nand _39446_ (_08186_, _07764_, _07782_);
  and _39447_ (_08187_, _08186_, _08185_);
  or _39448_ (_08189_, _08104_, _07763_);
  or _39449_ (_08191_, _08189_, _08187_);
  or _39450_ (_08192_, _08191_, _08184_);
  or _39451_ (_08193_, _08192_, _08122_);
  or _39452_ (_08194_, _08193_, _08182_);
  and _39453_ (_26842_[8], _08194_, _22762_);
  and _39454_ (_08196_, _06602_, _23778_);
  and _39455_ (_08197_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  or _39456_ (_01104_, _08197_, _08196_);
  and _39457_ (_08198_, _23903_, _23664_);
  and _39458_ (_08199_, _08198_, _23898_);
  not _39459_ (_08200_, _08198_);
  and _39460_ (_08201_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or _39461_ (_01130_, _08201_, _08199_);
  and _39462_ (_08204_, _07880_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _39463_ (_08206_, _07760_, _07940_);
  and _39464_ (_08207_, _07992_, _07790_);
  nor _39465_ (_08209_, _07880_, _07621_);
  or _39466_ (_08211_, _08209_, _08207_);
  and _39467_ (_08212_, _08211_, _08206_);
  or _39468_ (_08213_, _08212_, _08184_);
  and _39469_ (_08214_, _07608_, _07648_);
  and _39470_ (_08216_, _08211_, _08050_);
  or _39471_ (_08217_, _08216_, _08214_);
  or _39472_ (_08218_, _08217_, _08213_);
  or _39473_ (_08219_, _08218_, _08204_);
  and _39474_ (_26842_[9], _08219_, _22762_);
  and _39475_ (_08220_, _07947_, _07751_);
  not _39476_ (_08222_, _07756_);
  and _39477_ (_08223_, _08222_, _07655_);
  or _39478_ (_08224_, _08223_, _08220_);
  not _39479_ (_08225_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _39480_ (_08226_, _08040_, _08225_);
  and _39481_ (_08227_, _07878_, _07648_);
  and _39482_ (_08228_, _08227_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _39483_ (_08229_, _08122_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _39484_ (_08230_, _08229_, _07763_);
  or _39485_ (_08231_, _08230_, _08228_);
  or _39486_ (_08232_, _08231_, _08226_);
  or _39487_ (_08233_, _08232_, _08207_);
  or _39488_ (_08234_, _08233_, _08224_);
  or _39489_ (_08235_, _08234_, _08184_);
  and _39490_ (_26842_[10], _08235_, _22762_);
  and _39491_ (_08236_, _08198_, _23778_);
  and _39492_ (_08237_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or _39493_ (_01277_, _08237_, _08236_);
  and _39494_ (_08238_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  and _39495_ (_08239_, _05193_, _23898_);
  or _39496_ (_01285_, _08239_, _08238_);
  and _39497_ (_08241_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  and _39498_ (_08242_, _05193_, _23778_);
  or _39499_ (_01296_, _08242_, _08241_);
  nor _39500_ (_08243_, _24628_, rst);
  and _39501_ (_26888_, _08243_, _00289_);
  and _39502_ (_08244_, _07947_, _07754_);
  and _39503_ (_08245_, _08000_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _39504_ (_08246_, _08245_, _08244_);
  and _39505_ (_08247_, _07845_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _39506_ (_08248_, _08080_, _07763_);
  and _39507_ (_08249_, _08248_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _39508_ (_08250_, _07812_, _07984_);
  and _39509_ (_08251_, _08250_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _39510_ (_08252_, _08251_, _08184_);
  or _39511_ (_08253_, _08252_, _08249_);
  or _39512_ (_08254_, _08253_, _08220_);
  or _39513_ (_08255_, _08254_, _08247_);
  or _39514_ (_08256_, _08255_, _08207_);
  or _39515_ (_08257_, _08256_, _08246_);
  and _39516_ (_26842_[11], _08257_, _22762_);
  and _39517_ (_08259_, _02359_, _23707_);
  and _39518_ (_08260_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  or _39519_ (_01344_, _08260_, _08259_);
  and _39520_ (_08261_, _08198_, _23649_);
  and _39521_ (_08262_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or _39522_ (_01348_, _08262_, _08261_);
  and _39523_ (_08263_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  and _39524_ (_08264_, _05193_, _23649_);
  or _39525_ (_27228_, _08264_, _08263_);
  and _39526_ (_08265_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and _39527_ (_08266_, _04761_, _23898_);
  or _39528_ (_01372_, _08266_, _08265_);
  and _39529_ (_08267_, _08000_, _07782_);
  and _39530_ (_08268_, _08267_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _39531_ (_08269_, _07597_, _07648_);
  and _39532_ (_08270_, _08269_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nand _39533_ (_08271_, _08040_, _07940_);
  and _39534_ (_08272_, _08271_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _39535_ (_08273_, _07762_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _39536_ (_08274_, _08273_, _07992_);
  or _39537_ (_08275_, _08274_, _08272_);
  or _39538_ (_08276_, _08275_, _08270_);
  or _39539_ (_08277_, _08276_, _08268_);
  and _39540_ (_26842_[12], _08277_, _22762_);
  and _39541_ (_08278_, _04333_, _24654_);
  nand _39542_ (_08279_, _08278_, _23594_);
  or _39543_ (_08280_, _08278_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _39544_ (_08281_, _08280_, _04339_);
  and _39545_ (_08282_, _08281_, _08279_);
  nor _39546_ (_08283_, _04339_, _23702_);
  or _39547_ (_08284_, _08283_, _08282_);
  and _39548_ (_01382_, _08284_, _22762_);
  or _39549_ (_08285_, _04805_, _04725_);
  and _39550_ (_08286_, _08285_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _39551_ (_08287_, _08286_, _04768_);
  and _39552_ (_01384_, _08287_, _22762_);
  nor _39553_ (_01386_, _06776_, rst);
  and _39554_ (_08288_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  and _39555_ (_08289_, _05193_, _23747_);
  or _39556_ (_01393_, _08289_, _08288_);
  and _39557_ (_08290_, _08198_, _23747_);
  and _39558_ (_08291_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or _39559_ (_01396_, _08291_, _08290_);
  and _39560_ (_08292_, _02064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _39561_ (_08293_, _02066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or _39562_ (_01407_, _08293_, _08292_);
  or _39563_ (_08294_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _39564_ (_08295_, _08294_, _22762_);
  and _39565_ (_08296_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or _39566_ (_08297_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _39567_ (_08298_, _08297_, rxd_i);
  or _39568_ (_08299_, _08298_, _08296_);
  and _39569_ (_08300_, _08299_, _04589_);
  and _39570_ (_08301_, _04612_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _39571_ (_08302_, _08301_, _08300_);
  and _39572_ (_08303_, _04602_, rxd_i);
  or _39573_ (_08304_, _08303_, _04609_);
  or _39574_ (_08305_, _08304_, _08302_);
  and _39575_ (_01419_, _08305_, _08295_);
  or _39576_ (_08306_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _39577_ (_08307_, _00273_, _24729_);
  or _39578_ (_08308_, _08307_, _08306_);
  nand _39579_ (_08309_, _05838_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _39580_ (_08310_, _08309_, _08307_);
  or _39581_ (_08311_, _08310_, _05839_);
  and _39582_ (_08312_, _08311_, _08308_);
  and _39583_ (_08313_, _01975_, _24735_);
  or _39584_ (_08314_, _08313_, _08312_);
  nand _39585_ (_08315_, _08313_, _23702_);
  and _39586_ (_08316_, _08315_, _22762_);
  and _39587_ (_01438_, _08316_, _08314_);
  or _39588_ (_08317_, _08053_, _07763_);
  or _39589_ (_08318_, _08057_, _08122_);
  or _39590_ (_08319_, _08318_, _08317_);
  or _39591_ (_08320_, _08319_, _07879_);
  and _39592_ (_08321_, _08320_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _39593_ (_08322_, _07597_, _07577_);
  or _39594_ (_08323_, _08027_, _08322_);
  nor _39595_ (_08324_, _08000_, _07572_);
  or _39596_ (_08325_, _08324_, _08267_);
  and _39597_ (_08326_, _08325_, _07586_);
  or _39598_ (_08327_, _08326_, _08323_);
  or _39599_ (_08328_, _08327_, _08321_);
  and _39600_ (_26842_[13], _08328_, _22762_);
  and _39601_ (_08329_, _04743_, _04582_);
  and _39602_ (_08330_, _04727_, _08329_);
  nand _39603_ (_08331_, _08330_, _04770_);
  or _39604_ (_08332_, _08330_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _39605_ (_08333_, _08332_, _22762_);
  and _39606_ (_01452_, _08333_, _08331_);
  or _39607_ (_08334_, _06845_, rxd_i);
  nand _39608_ (_08335_, _08334_, _04595_);
  or _39609_ (_08336_, _04596_, _04578_);
  and _39610_ (_08337_, _08336_, _08335_);
  or _39611_ (_08338_, _04601_, _04579_);
  or _39612_ (_08339_, _08338_, _04594_);
  or _39613_ (_08340_, _08339_, _08337_);
  and _39614_ (_01455_, _08340_, _02066_);
  or _39615_ (_08341_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _39616_ (_08342_, _08341_, _22762_);
  nand _39617_ (_08343_, _02034_, _23702_);
  and _39618_ (_01457_, _08343_, _08342_);
  nand _39619_ (_08344_, _04454_, _04449_);
  and _39620_ (_08345_, _08344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _39621_ (_08346_, _08345_, _06799_);
  nor _39622_ (_08347_, _04448_, _06800_);
  and _39623_ (_08348_, _08347_, _08346_);
  or _39624_ (_08349_, _08348_, _04569_);
  nand _39625_ (_08350_, _08349_, _22762_);
  nor _39626_ (_01466_, _08350_, _04462_);
  and _39627_ (_08351_, _24201_, _24010_);
  not _39628_ (_08352_, _08351_);
  and _39629_ (_08353_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and _39630_ (_08354_, _08351_, _23747_);
  or _39631_ (_01495_, _08354_, _08353_);
  or _39632_ (_08355_, _07860_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _39633_ (_26842_[14], _08355_, _22762_);
  and _39634_ (_08356_, _23665_, _23649_);
  and _39635_ (_08357_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  or _39636_ (_01521_, _08357_, _08356_);
  and _39637_ (_08358_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and _39638_ (_08359_, _08351_, _23824_);
  or _39639_ (_01524_, _08359_, _08358_);
  and _39640_ (_08360_, _24005_, _23664_);
  and _39641_ (_08361_, _08360_, _23747_);
  not _39642_ (_08362_, _08360_);
  and _39643_ (_08363_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  or _39644_ (_01538_, _08363_, _08361_);
  and _39645_ (_08364_, _08360_, _23824_);
  and _39646_ (_08366_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  or _39647_ (_01542_, _08366_, _08364_);
  and _39648_ (_08367_, _23747_, _23665_);
  and _39649_ (_08368_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  or _39650_ (_27078_, _08368_, _08367_);
  and _39651_ (_08369_, _05410_, _23824_);
  and _39652_ (_08370_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  or _39653_ (_01566_, _08370_, _08369_);
  and _39654_ (_08371_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and _39655_ (_08372_, _06896_, _24050_);
  or _39656_ (_27022_, _08372_, _08371_);
  and _39657_ (_08373_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and _39658_ (_08374_, _06896_, _23707_);
  or _39659_ (_01690_, _08374_, _08373_);
  and _39660_ (_08375_, _24766_, _23911_);
  not _39661_ (_08376_, _08375_);
  and _39662_ (_08377_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  and _39663_ (_08378_, _08375_, _23898_);
  or _39664_ (_01694_, _08378_, _08377_);
  and _39665_ (_08379_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  and _39666_ (_08381_, _08375_, _23747_);
  or _39667_ (_01696_, _08381_, _08379_);
  and _39668_ (_08382_, _02359_, _23898_);
  and _39669_ (_08383_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  or _39670_ (_01750_, _08383_, _08382_);
  and _39671_ (_08384_, _02326_, _23898_);
  and _39672_ (_08385_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or _39673_ (_01761_, _08385_, _08384_);
  and _39674_ (_08386_, _02326_, _23649_);
  and _39675_ (_08387_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or _39676_ (_01780_, _08387_, _08386_);
  and _39677_ (_08388_, _02345_, _23946_);
  and _39678_ (_08389_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or _39679_ (_01784_, _08389_, _08388_);
  and _39680_ (_08390_, _02359_, _23946_);
  and _39681_ (_08391_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  or _39682_ (_01789_, _08391_, _08390_);
  and _39683_ (_08392_, _08010_, _08050_);
  not _39684_ (_08393_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _39685_ (_08394_, _08015_, _07585_);
  nor _39686_ (_08396_, _08394_, _08013_);
  and _39687_ (_08397_, _08015_, _08058_);
  not _39688_ (_08398_, _08397_);
  and _39689_ (_08399_, _08398_, _08396_);
  and _39690_ (_08400_, _08399_, _08015_);
  nor _39691_ (_08401_, _08400_, _08393_);
  and _39692_ (_08402_, _08015_, word_in[0]);
  and _39693_ (_08403_, _08402_, _08399_);
  or _39694_ (_08404_, _08403_, _08401_);
  or _39695_ (_08405_, _08404_, _08392_);
  and _39696_ (_08406_, _08000_, _07751_);
  and _39697_ (_08407_, _08006_, _08406_);
  not _39698_ (_08408_, _08407_);
  not _39699_ (_08409_, _08392_);
  or _39700_ (_08410_, _08409_, word_in[8]);
  and _39701_ (_08411_, _08410_, _08408_);
  and _39702_ (_08412_, _08411_, _08405_);
  and _39703_ (_08413_, _07790_, _08000_);
  and _39704_ (_08414_, _08028_, _08413_);
  and _39705_ (_08415_, _08407_, word_in[16]);
  or _39706_ (_08417_, _08415_, _08414_);
  or _39707_ (_08418_, _08417_, _08412_);
  not _39708_ (_08419_, _08414_);
  or _39709_ (_08420_, _08419_, word_in[24]);
  and _39710_ (_26843_[0], _08420_, _08418_);
  and _39711_ (_08422_, _08006_, word_in[17]);
  and _39712_ (_08423_, _08422_, _08406_);
  not _39713_ (_08425_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _39714_ (_08426_, _08400_, _08425_);
  and _39715_ (_08428_, _08015_, word_in[1]);
  and _39716_ (_08430_, _08428_, _08399_);
  or _39717_ (_08431_, _08430_, _08426_);
  and _39718_ (_08433_, _08431_, _08409_);
  and _39719_ (_08434_, _08392_, word_in[9]);
  or _39720_ (_08436_, _08434_, _08433_);
  and _39721_ (_08437_, _08436_, _08408_);
  or _39722_ (_08438_, _08437_, _08423_);
  and _39723_ (_08440_, _08438_, _08419_);
  and _39724_ (_08441_, _08414_, word_in[25]);
  or _39725_ (_26843_[1], _08441_, _08440_);
  and _39726_ (_08443_, _02359_, _23747_);
  and _39727_ (_08444_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  or _39728_ (_01806_, _08444_, _08443_);
  and _39729_ (_08445_, _08407_, word_in[18]);
  or _39730_ (_08446_, _08409_, word_in[10]);
  and _39731_ (_08447_, _08446_, _08408_);
  and _39732_ (_08448_, _08400_, word_in[2]);
  not _39733_ (_08450_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _39734_ (_08452_, _08400_, _08450_);
  or _39735_ (_08453_, _08452_, _08448_);
  or _39736_ (_08455_, _08453_, _08392_);
  and _39737_ (_08456_, _08455_, _08447_);
  or _39738_ (_08457_, _08456_, _08445_);
  and _39739_ (_08459_, _08457_, _08419_);
  and _39740_ (_08460_, _08414_, word_in[26]);
  or _39741_ (_26843_[2], _08460_, _08459_);
  and _39742_ (_08461_, _08028_, word_in[27]);
  and _39743_ (_08462_, _08461_, _08413_);
  or _39744_ (_08464_, _08409_, word_in[11]);
  and _39745_ (_08465_, _08464_, _08408_);
  not _39746_ (_08467_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _39747_ (_08468_, _08400_, _08467_);
  and _39748_ (_08469_, _08400_, word_in[3]);
  or _39749_ (_08470_, _08469_, _08468_);
  or _39750_ (_08471_, _08470_, _08392_);
  and _39751_ (_08472_, _08471_, _08465_);
  and _39752_ (_08473_, _08407_, word_in[19]);
  or _39753_ (_08474_, _08473_, _08472_);
  and _39754_ (_08475_, _08474_, _08419_);
  or _39755_ (_26843_[3], _08475_, _08462_);
  and _39756_ (_08477_, _06506_, _23911_);
  not _39757_ (_08478_, _08477_);
  and _39758_ (_08479_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  and _39759_ (_08480_, _08477_, _23707_);
  or _39760_ (_26980_, _08480_, _08479_);
  and _39761_ (_08481_, _08028_, word_in[28]);
  and _39762_ (_08482_, _08481_, _08413_);
  or _39763_ (_08483_, _08409_, word_in[12]);
  and _39764_ (_08484_, _08483_, _08408_);
  not _39765_ (_08485_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _39766_ (_08486_, _08400_, _08485_);
  and _39767_ (_08488_, _08400_, word_in[4]);
  or _39768_ (_08489_, _08488_, _08486_);
  or _39769_ (_08490_, _08489_, _08392_);
  and _39770_ (_08491_, _08490_, _08484_);
  and _39771_ (_08492_, _08407_, word_in[20]);
  or _39772_ (_08493_, _08492_, _08491_);
  and _39773_ (_08494_, _08493_, _08419_);
  or _39774_ (_26843_[4], _08494_, _08482_);
  and _39775_ (_08495_, _08028_, word_in[29]);
  and _39776_ (_08497_, _08495_, _08413_);
  and _39777_ (_08498_, _08407_, word_in[21]);
  not _39778_ (_08499_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _39779_ (_08500_, _08400_, _08499_);
  and _39780_ (_08501_, _08015_, word_in[5]);
  and _39781_ (_08502_, _08501_, _08400_);
  or _39782_ (_08503_, _08502_, _08500_);
  or _39783_ (_08504_, _08503_, _08392_);
  or _39784_ (_08505_, _08409_, word_in[13]);
  and _39785_ (_08506_, _08505_, _08408_);
  and _39786_ (_08507_, _08506_, _08504_);
  or _39787_ (_08508_, _08507_, _08498_);
  and _39788_ (_08509_, _08508_, _08419_);
  or _39789_ (_26843_[5], _08509_, _08497_);
  and _39790_ (_08510_, _08028_, word_in[30]);
  and _39791_ (_08511_, _08510_, _08413_);
  and _39792_ (_08512_, _08407_, word_in[22]);
  or _39793_ (_08513_, _08409_, word_in[14]);
  and _39794_ (_08514_, _08513_, _08408_);
  not _39795_ (_08515_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _39796_ (_08516_, _08400_, _08515_);
  and _39797_ (_08517_, _08400_, word_in[6]);
  or _39798_ (_08518_, _08517_, _08516_);
  or _39799_ (_08519_, _08518_, _08392_);
  and _39800_ (_08520_, _08519_, _08514_);
  or _39801_ (_08521_, _08520_, _08512_);
  and _39802_ (_08523_, _08521_, _08419_);
  or _39803_ (_26843_[6], _08523_, _08511_);
  and _39804_ (_08524_, _05410_, _23898_);
  and _39805_ (_08525_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  or _39806_ (_01820_, _08525_, _08524_);
  or _39807_ (_08527_, _08409_, word_in[15]);
  and _39808_ (_08528_, _08527_, _08408_);
  nor _39809_ (_08529_, _08400_, _07837_);
  and _39810_ (_08530_, _08400_, word_in[7]);
  or _39811_ (_08531_, _08530_, _08529_);
  or _39812_ (_08532_, _08531_, _08392_);
  and _39813_ (_08533_, _08532_, _08528_);
  and _39814_ (_08534_, _08407_, word_in[23]);
  or _39815_ (_08535_, _08534_, _08533_);
  and _39816_ (_08536_, _08535_, _08419_);
  and _39817_ (_08537_, _08414_, word_in[31]);
  or _39818_ (_26843_[7], _08537_, _08536_);
  and _39819_ (_08539_, _06602_, _23747_);
  and _39820_ (_08540_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  or _39821_ (_01833_, _08540_, _08539_);
  and _39822_ (_08541_, _06602_, _23707_);
  and _39823_ (_08542_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  or _39824_ (_01837_, _08542_, _08541_);
  and _39825_ (_08543_, _06602_, _24050_);
  and _39826_ (_08545_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  or _39827_ (_27157_, _08545_, _08543_);
  and _39828_ (_08546_, _05042_, _24050_);
  and _39829_ (_08547_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or _39830_ (_01860_, _08547_, _08546_);
  and _39831_ (_08548_, _01809_, _24275_);
  and _39832_ (_08549_, _08548_, _23747_);
  not _39833_ (_08550_, _08548_);
  and _39834_ (_08551_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  or _39835_ (_01866_, _08551_, _08549_);
  and _39836_ (_08552_, _08028_, _08406_);
  and _39837_ (_08553_, _08010_, _07780_);
  and _39838_ (_08554_, _08553_, _07766_);
  not _39839_ (_08555_, _08554_);
  not _39840_ (_08556_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _39841_ (_08557_, _08013_, _07586_);
  and _39842_ (_08558_, _08557_, _08398_);
  nor _39843_ (_08559_, _08558_, _08556_);
  and _39844_ (_08560_, _08558_, _08402_);
  or _39845_ (_08561_, _08560_, _08559_);
  and _39846_ (_08562_, _08561_, _08555_);
  and _39847_ (_08563_, _08006_, _07754_);
  and _39848_ (_08564_, _08563_, _07882_);
  and _39849_ (_08565_, _08554_, word_in[8]);
  or _39850_ (_08566_, _08565_, _08564_);
  or _39851_ (_08567_, _08566_, _08562_);
  not _39852_ (_08568_, _08564_);
  or _39853_ (_08569_, _08568_, word_in[16]);
  and _39854_ (_08570_, _08569_, _08567_);
  or _39855_ (_08571_, _08570_, _08552_);
  not _39856_ (_08573_, _08552_);
  or _39857_ (_08574_, _08573_, word_in[24]);
  and _39858_ (_26850_[0], _08574_, _08571_);
  not _39859_ (_08575_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _39860_ (_08576_, _08558_, _08575_);
  and _39861_ (_08577_, _08558_, _08428_);
  or _39862_ (_08578_, _08577_, _08576_);
  and _39863_ (_08579_, _08578_, _08555_);
  and _39864_ (_08580_, _08554_, word_in[9]);
  or _39865_ (_08581_, _08580_, _08564_);
  or _39866_ (_08582_, _08581_, _08579_);
  or _39867_ (_08583_, _08568_, word_in[17]);
  and _39868_ (_08584_, _08583_, _08582_);
  or _39869_ (_08585_, _08584_, _08552_);
  or _39870_ (_08586_, _08573_, word_in[25]);
  and _39871_ (_26850_[1], _08586_, _08585_);
  and _39872_ (_08587_, _08548_, _23707_);
  and _39873_ (_08588_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  or _39874_ (_01878_, _08588_, _08587_);
  not _39875_ (_08589_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _39876_ (_08590_, _08558_, _08589_);
  and _39877_ (_08591_, _08015_, word_in[2]);
  and _39878_ (_08592_, _08558_, _08591_);
  or _39879_ (_08593_, _08592_, _08590_);
  and _39880_ (_08594_, _08593_, _08555_);
  and _39881_ (_08595_, _08554_, word_in[10]);
  or _39882_ (_08596_, _08595_, _08564_);
  or _39883_ (_08597_, _08596_, _08594_);
  or _39884_ (_08598_, _08568_, word_in[18]);
  and _39885_ (_08599_, _08598_, _08597_);
  or _39886_ (_08600_, _08599_, _08552_);
  or _39887_ (_08601_, _08573_, word_in[26]);
  and _39888_ (_26850_[2], _08601_, _08600_);
  not _39889_ (_08602_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _39890_ (_08603_, _08558_, _08602_);
  and _39891_ (_08604_, _08015_, word_in[3]);
  and _39892_ (_08605_, _08558_, _08604_);
  or _39893_ (_08606_, _08605_, _08603_);
  and _39894_ (_08607_, _08606_, _08555_);
  and _39895_ (_08608_, _08554_, word_in[11]);
  or _39896_ (_08609_, _08608_, _08564_);
  or _39897_ (_08610_, _08609_, _08607_);
  or _39898_ (_08611_, _08568_, word_in[19]);
  and _39899_ (_08612_, _08611_, _08610_);
  or _39900_ (_08613_, _08612_, _08552_);
  or _39901_ (_08614_, _08573_, word_in[27]);
  and _39902_ (_26850_[3], _08614_, _08613_);
  and _39903_ (_08615_, _08548_, _23946_);
  and _39904_ (_08616_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or _39905_ (_01881_, _08616_, _08615_);
  not _39906_ (_08617_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _39907_ (_08618_, _08558_, _08617_);
  and _39908_ (_08619_, _08015_, word_in[4]);
  and _39909_ (_08620_, _08558_, _08619_);
  or _39910_ (_08621_, _08620_, _08618_);
  and _39911_ (_08622_, _08621_, _08555_);
  and _39912_ (_08623_, _08554_, word_in[12]);
  or _39913_ (_08624_, _08623_, _08564_);
  or _39914_ (_08625_, _08624_, _08622_);
  or _39915_ (_08626_, _08568_, word_in[20]);
  and _39916_ (_08627_, _08626_, _08625_);
  or _39917_ (_08628_, _08627_, _08552_);
  or _39918_ (_08629_, _08573_, word_in[28]);
  and _39919_ (_26850_[4], _08629_, _08628_);
  not _39920_ (_08630_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _39921_ (_08631_, _08558_, _08630_);
  and _39922_ (_08632_, _08558_, _08501_);
  or _39923_ (_08633_, _08632_, _08631_);
  and _39924_ (_08634_, _08633_, _08555_);
  and _39925_ (_08635_, _08554_, word_in[13]);
  or _39926_ (_08636_, _08635_, _08564_);
  or _39927_ (_08637_, _08636_, _08634_);
  or _39928_ (_08638_, _08568_, word_in[21]);
  and _39929_ (_08639_, _08638_, _08637_);
  or _39930_ (_08640_, _08639_, _08552_);
  or _39931_ (_08641_, _08573_, word_in[29]);
  and _39932_ (_26850_[5], _08641_, _08640_);
  and _39933_ (_08642_, _02325_, _23784_);
  and _39934_ (_08643_, _08642_, _23946_);
  not _39935_ (_08644_, _08642_);
  and _39936_ (_08645_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  or _39937_ (_01885_, _08645_, _08643_);
  not _39938_ (_08646_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _39939_ (_08647_, _08558_, _08646_);
  and _39940_ (_08648_, _08015_, word_in[6]);
  and _39941_ (_08649_, _08558_, _08648_);
  or _39942_ (_08650_, _08649_, _08647_);
  and _39943_ (_08651_, _08650_, _08555_);
  and _39944_ (_08652_, _08554_, word_in[14]);
  or _39945_ (_08653_, _08652_, _08564_);
  or _39946_ (_08654_, _08653_, _08651_);
  or _39947_ (_08655_, _08568_, word_in[22]);
  and _39948_ (_08656_, _08655_, _08654_);
  or _39949_ (_08657_, _08656_, _08552_);
  or _39950_ (_08658_, _08573_, word_in[30]);
  and _39951_ (_26850_[6], _08658_, _08657_);
  nor _39952_ (_08659_, _08558_, _07675_);
  and _39953_ (_08660_, _08558_, _08019_);
  or _39954_ (_08661_, _08660_, _08659_);
  and _39955_ (_08662_, _08661_, _08555_);
  and _39956_ (_08663_, _08554_, word_in[15]);
  or _39957_ (_08664_, _08663_, _08564_);
  or _39958_ (_08665_, _08664_, _08662_);
  or _39959_ (_08666_, _08568_, word_in[23]);
  and _39960_ (_08667_, _08666_, _08665_);
  or _39961_ (_08668_, _08667_, _08552_);
  or _39962_ (_08669_, _08573_, word_in[31]);
  and _39963_ (_26850_[7], _08669_, _08668_);
  and _39964_ (_08670_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  and _39965_ (_08671_, _08477_, _24050_);
  or _39966_ (_01901_, _08671_, _08670_);
  and _39967_ (_08673_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and _39968_ (_08674_, _07513_, _23707_);
  or _39969_ (_01928_, _08674_, _08673_);
  and _39970_ (_08675_, _06544_, _23747_);
  and _39971_ (_08676_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or _39972_ (_01933_, _08676_, _08675_);
  and _39973_ (_08677_, _08028_, _08050_);
  and _39974_ (_08678_, _08006_, word_in[16]);
  and _39975_ (_08679_, _08006_, _07780_);
  and _39976_ (_08680_, _08679_, _07882_);
  not _39977_ (_08681_, _08680_);
  or _39978_ (_08682_, _08681_, _08678_);
  and _39979_ (_08683_, _08010_, _07790_);
  and _39980_ (_08684_, _08683_, _07766_);
  not _39981_ (_08685_, _08684_);
  not _39982_ (_08686_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  not _39983_ (_08687_, _08013_);
  and _39984_ (_08688_, _08394_, _08687_);
  and _39985_ (_08689_, _08688_, _08176_);
  nor _39986_ (_08690_, _08689_, _08686_);
  and _39987_ (_08691_, _08689_, _08402_);
  or _39988_ (_08692_, _08691_, _08690_);
  and _39989_ (_08693_, _08692_, _08685_);
  and _39990_ (_08694_, _08684_, word_in[8]);
  or _39991_ (_08695_, _08694_, _08680_);
  or _39992_ (_08696_, _08695_, _08693_);
  and _39993_ (_08697_, _08696_, _08682_);
  or _39994_ (_08698_, _08697_, _08677_);
  not _39995_ (_08699_, _08677_);
  or _39996_ (_08700_, _08699_, word_in[24]);
  and _39997_ (_26851_[0], _08700_, _08698_);
  or _39998_ (_08701_, _08681_, _08422_);
  not _39999_ (_08702_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _40000_ (_08703_, _08689_, _08702_);
  and _40001_ (_08704_, _08689_, _08428_);
  or _40002_ (_08705_, _08704_, _08703_);
  and _40003_ (_08706_, _08705_, _08685_);
  and _40004_ (_08707_, _08684_, word_in[9]);
  or _40005_ (_08708_, _08707_, _08680_);
  or _40006_ (_08709_, _08708_, _08706_);
  and _40007_ (_08710_, _08709_, _08701_);
  or _40008_ (_08711_, _08710_, _08677_);
  or _40009_ (_08712_, _08699_, word_in[25]);
  and _40010_ (_26851_[1], _08712_, _08711_);
  and _40011_ (_08713_, _06544_, _23707_);
  and _40012_ (_08714_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or _40013_ (_01943_, _08714_, _08713_);
  and _40014_ (_08715_, _08006_, word_in[18]);
  or _40015_ (_08716_, _08681_, _08715_);
  not _40016_ (_08717_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _40017_ (_08718_, _08689_, _08717_);
  and _40018_ (_08719_, _08689_, _08591_);
  or _40019_ (_08720_, _08719_, _08718_);
  and _40020_ (_08721_, _08720_, _08685_);
  and _40021_ (_08722_, _08684_, word_in[10]);
  or _40022_ (_08723_, _08722_, _08680_);
  or _40023_ (_08724_, _08723_, _08721_);
  and _40024_ (_08725_, _08724_, _08716_);
  or _40025_ (_08726_, _08725_, _08677_);
  or _40026_ (_08727_, _08699_, word_in[26]);
  and _40027_ (_26851_[2], _08727_, _08726_);
  and _40028_ (_08728_, _08006_, word_in[19]);
  or _40029_ (_08729_, _08681_, _08728_);
  not _40030_ (_08730_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor _40031_ (_08731_, _08689_, _08730_);
  and _40032_ (_08732_, _08689_, _08604_);
  or _40033_ (_08733_, _08732_, _08731_);
  and _40034_ (_08734_, _08733_, _08685_);
  and _40035_ (_08735_, _08684_, word_in[11]);
  or _40036_ (_08736_, _08735_, _08680_);
  or _40037_ (_08737_, _08736_, _08734_);
  and _40038_ (_08738_, _08737_, _08729_);
  or _40039_ (_08739_, _08738_, _08677_);
  or _40040_ (_08741_, _08699_, word_in[27]);
  and _40041_ (_26851_[3], _08741_, _08739_);
  and _40042_ (_08742_, _06530_, _23946_);
  and _40043_ (_08743_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  or _40044_ (_01946_, _08743_, _08742_);
  and _40045_ (_08744_, _08006_, word_in[20]);
  or _40046_ (_08745_, _08681_, _08744_);
  not _40047_ (_08746_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _40048_ (_08747_, _08689_, _08746_);
  and _40049_ (_08748_, _08689_, _08619_);
  or _40050_ (_08750_, _08748_, _08747_);
  and _40051_ (_08751_, _08750_, _08685_);
  and _40052_ (_08752_, _08684_, word_in[12]);
  or _40053_ (_08753_, _08752_, _08680_);
  or _40054_ (_08754_, _08753_, _08751_);
  and _40055_ (_08755_, _08754_, _08745_);
  or _40056_ (_08756_, _08755_, _08677_);
  or _40057_ (_08757_, _08699_, word_in[28]);
  and _40058_ (_26851_[4], _08757_, _08756_);
  and _40059_ (_08758_, _08006_, word_in[21]);
  or _40060_ (_08759_, _08681_, _08758_);
  not _40061_ (_08760_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _40062_ (_08761_, _08689_, _08760_);
  and _40063_ (_08762_, _08689_, _08501_);
  or _40064_ (_08763_, _08762_, _08761_);
  and _40065_ (_08764_, _08763_, _08685_);
  and _40066_ (_08766_, _08684_, word_in[13]);
  or _40067_ (_08767_, _08766_, _08680_);
  or _40068_ (_08768_, _08767_, _08764_);
  and _40069_ (_08769_, _08768_, _08759_);
  or _40070_ (_08770_, _08769_, _08677_);
  or _40071_ (_08772_, _08699_, word_in[29]);
  and _40072_ (_26851_[5], _08772_, _08770_);
  and _40073_ (_08774_, _08006_, word_in[22]);
  or _40074_ (_08775_, _08681_, _08774_);
  not _40075_ (_08776_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _40076_ (_08778_, _08689_, _08776_);
  and _40077_ (_08779_, _08689_, _08648_);
  or _40078_ (_08780_, _08779_, _08778_);
  and _40079_ (_08781_, _08780_, _08685_);
  and _40080_ (_08782_, _08684_, word_in[14]);
  or _40081_ (_08783_, _08782_, _08680_);
  or _40082_ (_08784_, _08783_, _08781_);
  and _40083_ (_08785_, _08784_, _08775_);
  or _40084_ (_08786_, _08785_, _08677_);
  or _40085_ (_08787_, _08699_, word_in[30]);
  and _40086_ (_26851_[6], _08787_, _08786_);
  or _40087_ (_08788_, _08681_, _08033_);
  nor _40088_ (_08789_, _08689_, _07829_);
  and _40089_ (_08790_, _08689_, _08019_);
  or _40090_ (_08791_, _08790_, _08789_);
  and _40091_ (_08792_, _08791_, _08685_);
  and _40092_ (_08793_, _08684_, word_in[15]);
  or _40093_ (_08794_, _08793_, _08680_);
  or _40094_ (_08795_, _08794_, _08792_);
  and _40095_ (_08796_, _08795_, _08788_);
  or _40096_ (_08797_, _08796_, _08677_);
  or _40097_ (_08798_, _08699_, word_in[31]);
  and _40098_ (_26851_[7], _08798_, _08797_);
  and _40099_ (_08799_, _25078_, _23664_);
  and _40100_ (_08800_, _08799_, _23898_);
  not _40101_ (_08801_, _08799_);
  and _40102_ (_08802_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  or _40103_ (_27077_, _08802_, _08800_);
  and _40104_ (_08803_, _06517_, _23946_);
  and _40105_ (_08804_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or _40106_ (_01976_, _08804_, _08803_);
  and _40107_ (_08805_, _06651_, _23649_);
  and _40108_ (_08806_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  or _40109_ (_01991_, _08806_, _08805_);
  and _40110_ (_08807_, _08011_, _07766_);
  not _40111_ (_08808_, _08807_);
  not _40112_ (_08809_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _40113_ (_08810_, _08398_, _08014_);
  nor _40114_ (_08811_, _08810_, _08809_);
  and _40115_ (_08812_, _08810_, _08402_);
  or _40116_ (_08813_, _08812_, _08811_);
  and _40117_ (_08814_, _08813_, _08808_);
  and _40118_ (_08815_, _08006_, _07790_);
  and _40119_ (_08816_, _08815_, _07882_);
  and _40120_ (_08817_, _08807_, word_in[8]);
  or _40121_ (_08818_, _08817_, _08816_);
  or _40122_ (_08819_, _08818_, _08814_);
  and _40123_ (_08820_, _08028_, _08080_);
  not _40124_ (_08821_, _08820_);
  not _40125_ (_08822_, _08816_);
  or _40126_ (_08823_, _08822_, _08678_);
  and _40127_ (_08824_, _08823_, _08821_);
  and _40128_ (_08825_, _08824_, _08819_);
  and _40129_ (_08827_, _08820_, word_in[24]);
  or _40130_ (_26852_[0], _08827_, _08825_);
  and _40131_ (_08829_, _08820_, word_in[25]);
  not _40132_ (_08830_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _40133_ (_08831_, _08810_, _08830_);
  and _40134_ (_08832_, _08810_, _08428_);
  or _40135_ (_08833_, _08832_, _08831_);
  and _40136_ (_08834_, _08833_, _08808_);
  and _40137_ (_08835_, _08807_, word_in[9]);
  or _40138_ (_08836_, _08835_, _08816_);
  or _40139_ (_08837_, _08836_, _08834_);
  or _40140_ (_08838_, _08822_, word_in[17]);
  and _40141_ (_08839_, _08838_, _08821_);
  and _40142_ (_08840_, _08839_, _08837_);
  or _40143_ (_26852_[1], _08840_, _08829_);
  and _40144_ (_08841_, _06755_, _23946_);
  and _40145_ (_08842_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or _40146_ (_02003_, _08842_, _08841_);
  and _40147_ (_08843_, _08820_, word_in[26]);
  not _40148_ (_08844_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor _40149_ (_08845_, _08810_, _08844_);
  and _40150_ (_08846_, _08810_, _08591_);
  or _40151_ (_08847_, _08846_, _08845_);
  and _40152_ (_08848_, _08847_, _08808_);
  and _40153_ (_08849_, _08807_, word_in[10]);
  or _40154_ (_08850_, _08849_, _08816_);
  or _40155_ (_08851_, _08850_, _08848_);
  or _40156_ (_08853_, _08822_, word_in[18]);
  and _40157_ (_08854_, _08853_, _08821_);
  and _40158_ (_08855_, _08854_, _08851_);
  or _40159_ (_26852_[2], _08855_, _08843_);
  and _40160_ (_08856_, _08820_, word_in[27]);
  not _40161_ (_08857_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _40162_ (_08858_, _08810_, _08857_);
  and _40163_ (_08859_, _08810_, _08604_);
  or _40164_ (_08860_, _08859_, _08858_);
  and _40165_ (_08861_, _08860_, _08808_);
  and _40166_ (_08862_, _08807_, word_in[11]);
  or _40167_ (_08863_, _08862_, _08816_);
  or _40168_ (_08864_, _08863_, _08861_);
  or _40169_ (_08865_, _08822_, word_in[19]);
  and _40170_ (_08866_, _08865_, _08821_);
  and _40171_ (_08867_, _08866_, _08864_);
  or _40172_ (_26852_[3], _08867_, _08856_);
  and _40173_ (_08868_, _06755_, _23747_);
  and _40174_ (_08869_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or _40175_ (_02008_, _08869_, _08868_);
  not _40176_ (_08870_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _40177_ (_08871_, _08810_, _08870_);
  and _40178_ (_08872_, _08810_, _08619_);
  or _40179_ (_08873_, _08872_, _08871_);
  and _40180_ (_08874_, _08873_, _08808_);
  and _40181_ (_08875_, _08807_, word_in[12]);
  or _40182_ (_08876_, _08875_, _08816_);
  or _40183_ (_08877_, _08876_, _08874_);
  or _40184_ (_08878_, _08822_, word_in[20]);
  and _40185_ (_08879_, _08878_, _08821_);
  and _40186_ (_08880_, _08879_, _08877_);
  and _40187_ (_08881_, _08820_, word_in[28]);
  or _40188_ (_26852_[4], _08881_, _08880_);
  not _40189_ (_08883_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _40190_ (_08884_, _08810_, _08883_);
  and _40191_ (_08885_, _08810_, _08501_);
  or _40192_ (_08886_, _08885_, _08884_);
  and _40193_ (_08887_, _08886_, _08808_);
  and _40194_ (_08888_, _08807_, word_in[13]);
  or _40195_ (_08889_, _08888_, _08816_);
  or _40196_ (_08890_, _08889_, _08887_);
  or _40197_ (_08891_, _08822_, _08758_);
  and _40198_ (_08892_, _08891_, _08821_);
  and _40199_ (_08893_, _08892_, _08890_);
  and _40200_ (_08894_, _08820_, word_in[29]);
  or _40201_ (_26852_[5], _08894_, _08893_);
  and _40202_ (_08895_, _06646_, _23824_);
  and _40203_ (_08896_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or _40204_ (_02013_, _08896_, _08895_);
  and _40205_ (_08897_, _08820_, word_in[30]);
  not _40206_ (_08898_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _40207_ (_08899_, _08810_, _08898_);
  and _40208_ (_08900_, _08810_, _08648_);
  or _40209_ (_08901_, _08900_, _08899_);
  and _40210_ (_08902_, _08901_, _08808_);
  and _40211_ (_08903_, _08807_, word_in[14]);
  or _40212_ (_08904_, _08903_, _08816_);
  or _40213_ (_08905_, _08904_, _08902_);
  or _40214_ (_08906_, _08822_, word_in[22]);
  and _40215_ (_08907_, _08906_, _08821_);
  and _40216_ (_08910_, _08907_, _08905_);
  or _40217_ (_26852_[6], _08910_, _08897_);
  nor _40218_ (_08911_, _08810_, _07696_);
  and _40219_ (_08912_, _08810_, _08019_);
  or _40220_ (_08913_, _08912_, _08911_);
  and _40221_ (_08914_, _08913_, _08808_);
  and _40222_ (_08915_, _08807_, word_in[15]);
  or _40223_ (_08916_, _08915_, _08816_);
  or _40224_ (_08917_, _08916_, _08914_);
  or _40225_ (_08918_, _08822_, word_in[23]);
  and _40226_ (_08919_, _08918_, _08821_);
  and _40227_ (_08920_, _08919_, _08917_);
  and _40228_ (_08921_, _08820_, word_in[31]);
  or _40229_ (_26852_[7], _08921_, _08920_);
  and _40230_ (_08922_, _06646_, _23946_);
  and _40231_ (_08923_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or _40232_ (_02033_, _08923_, _08922_);
  and _40233_ (_08924_, _05710_, _23898_);
  and _40234_ (_08925_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  or _40235_ (_02062_, _08925_, _08924_);
  and _40236_ (_08927_, _06639_, _23824_);
  and _40237_ (_08928_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or _40238_ (_02068_, _08928_, _08927_);
  and _40239_ (_08929_, _08028_, _07942_);
  and _40240_ (_08930_, _08929_, _07948_);
  and _40241_ (_08932_, _08930_, _07790_);
  and _40242_ (_08933_, _08006_, _08053_);
  not _40243_ (_08934_, _08933_);
  or _40244_ (_08935_, _08934_, word_in[16]);
  and _40245_ (_08936_, _08010_, _08057_);
  not _40246_ (_08937_, _08936_);
  not _40247_ (_08938_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _40248_ (_08940_, _08015_, _07762_);
  and _40249_ (_08941_, _08940_, _08396_);
  nor _40250_ (_08942_, _08941_, _08938_);
  and _40251_ (_08944_, _08941_, _08402_);
  or _40252_ (_08945_, _08944_, _08942_);
  and _40253_ (_08946_, _08945_, _08937_);
  and _40254_ (_08948_, _08936_, word_in[8]);
  or _40255_ (_08949_, _08948_, _08933_);
  or _40256_ (_08950_, _08949_, _08946_);
  and _40257_ (_08952_, _08950_, _08935_);
  or _40258_ (_08953_, _08952_, _08932_);
  and _40259_ (_08954_, _08028_, word_in[24]);
  not _40260_ (_08955_, _08932_);
  or _40261_ (_08956_, _08955_, _08954_);
  and _40262_ (_26853_[0], _08956_, _08953_);
  not _40263_ (_08957_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _40264_ (_08958_, _08941_, _08957_);
  and _40265_ (_08960_, _08941_, word_in[1]);
  or _40266_ (_08961_, _08960_, _08958_);
  and _40267_ (_08962_, _08961_, _08937_);
  and _40268_ (_08964_, _08936_, word_in[9]);
  or _40269_ (_08966_, _08964_, _08962_);
  or _40270_ (_08967_, _08966_, _08933_);
  nor _40271_ (_08968_, _08934_, _08422_);
  nor _40272_ (_08970_, _08968_, _08932_);
  and _40273_ (_08972_, _08970_, _08967_);
  and _40274_ (_08973_, _08028_, word_in[25]);
  and _40275_ (_08974_, _08932_, _08973_);
  or _40276_ (_26853_[1], _08974_, _08972_);
  and _40277_ (_08976_, _06639_, _23707_);
  and _40278_ (_08978_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or _40279_ (_02085_, _08978_, _08976_);
  not _40280_ (_08979_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _40281_ (_08980_, _08941_, _08979_);
  and _40282_ (_08982_, _08941_, word_in[2]);
  or _40283_ (_08984_, _08982_, _08980_);
  and _40284_ (_08985_, _08984_, _08937_);
  and _40285_ (_08986_, _08936_, word_in[10]);
  or _40286_ (_08987_, _08986_, _08985_);
  and _40287_ (_08989_, _08987_, _08934_);
  and _40288_ (_08990_, _08933_, word_in[18]);
  or _40289_ (_08991_, _08990_, _08989_);
  and _40290_ (_08992_, _08991_, _08955_);
  and _40291_ (_08993_, _08028_, word_in[26]);
  and _40292_ (_08994_, _08932_, _08993_);
  or _40293_ (_26853_[2], _08994_, _08992_);
  not _40294_ (_08996_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _40295_ (_08997_, _08941_, _08996_);
  and _40296_ (_08998_, _08941_, word_in[3]);
  or _40297_ (_08999_, _08998_, _08997_);
  and _40298_ (_09000_, _08999_, _08937_);
  and _40299_ (_09001_, _08936_, word_in[11]);
  or _40300_ (_09003_, _09001_, _09000_);
  or _40301_ (_09004_, _09003_, _08933_);
  nor _40302_ (_09005_, _08934_, _08728_);
  nor _40303_ (_09006_, _09005_, _08932_);
  and _40304_ (_09007_, _09006_, _09004_);
  and _40305_ (_09008_, _08932_, _08461_);
  or _40306_ (_26853_[3], _09008_, _09007_);
  or _40307_ (_09012_, _08934_, word_in[20]);
  not _40308_ (_09013_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _40309_ (_09015_, _08941_, _09013_);
  and _40310_ (_09016_, _08941_, _08619_);
  or _40311_ (_09017_, _09016_, _09015_);
  or _40312_ (_09019_, _09017_, _08936_);
  or _40313_ (_09020_, _08937_, word_in[12]);
  and _40314_ (_09021_, _09020_, _09019_);
  or _40315_ (_09023_, _09021_, _08933_);
  and _40316_ (_09024_, _09023_, _09012_);
  or _40317_ (_09026_, _09024_, _08932_);
  or _40318_ (_09027_, _08955_, _08481_);
  and _40319_ (_26853_[4], _09027_, _09026_);
  or _40320_ (_09028_, _08934_, word_in[21]);
  not _40321_ (_09029_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _40322_ (_09030_, _08941_, _09029_);
  and _40323_ (_09031_, _08941_, _08501_);
  or _40324_ (_09032_, _09031_, _09030_);
  or _40325_ (_09033_, _09032_, _08936_);
  or _40326_ (_09034_, _08937_, word_in[13]);
  and _40327_ (_09036_, _09034_, _09033_);
  or _40328_ (_09037_, _09036_, _08933_);
  and _40329_ (_09039_, _09037_, _09028_);
  or _40330_ (_09040_, _09039_, _08932_);
  or _40331_ (_09041_, _08955_, _08495_);
  and _40332_ (_26853_[5], _09041_, _09040_);
  or _40333_ (_09042_, _08934_, word_in[22]);
  not _40334_ (_09043_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _40335_ (_09044_, _08941_, _09043_);
  and _40336_ (_09045_, _08941_, _08648_);
  or _40337_ (_09046_, _09045_, _09044_);
  or _40338_ (_09048_, _09046_, _08936_);
  or _40339_ (_09050_, _08937_, word_in[14]);
  and _40340_ (_09051_, _09050_, _09048_);
  or _40341_ (_09052_, _09051_, _08933_);
  and _40342_ (_09053_, _09052_, _09042_);
  or _40343_ (_09054_, _09053_, _08932_);
  or _40344_ (_09055_, _08955_, _08510_);
  and _40345_ (_26853_[6], _09055_, _09054_);
  and _40346_ (_09057_, _25748_, _23649_);
  and _40347_ (_09058_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or _40348_ (_02098_, _09058_, _09057_);
  nor _40349_ (_09060_, _08941_, _07852_);
  and _40350_ (_09062_, _08941_, word_in[7]);
  or _40351_ (_09063_, _09062_, _09060_);
  and _40352_ (_09064_, _09063_, _08937_);
  and _40353_ (_09065_, _08936_, word_in[15]);
  or _40354_ (_09066_, _09065_, _09064_);
  and _40355_ (_09067_, _09066_, _08934_);
  and _40356_ (_09068_, _08933_, word_in[23]);
  or _40357_ (_09069_, _09068_, _09067_);
  and _40358_ (_09070_, _09069_, _08955_);
  and _40359_ (_09072_, _08028_, word_in[31]);
  and _40360_ (_09073_, _08932_, _09072_);
  or _40361_ (_26853_[7], _09073_, _09070_);
  and _40362_ (_09076_, _08563_, _08227_);
  not _40363_ (_09077_, _09076_);
  and _40364_ (_09078_, _08553_, _07845_);
  not _40365_ (_09080_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _40366_ (_09082_, _08940_, _08557_);
  nor _40367_ (_09083_, _09082_, _09080_);
  and _40368_ (_09084_, _09082_, word_in[0]);
  nor _40369_ (_09085_, _09084_, _09083_);
  nor _40370_ (_09087_, _09085_, _09078_);
  and _40371_ (_09088_, _09078_, word_in[8]);
  or _40372_ (_09089_, _09088_, _09087_);
  and _40373_ (_09090_, _09089_, _09077_);
  and _40374_ (_09091_, _08930_, _07751_);
  and _40375_ (_09092_, _09076_, _08678_);
  or _40376_ (_09093_, _09092_, _09091_);
  or _40377_ (_09095_, _09093_, _09090_);
  not _40378_ (_09096_, _09091_);
  or _40379_ (_09097_, _09096_, word_in[24]);
  and _40380_ (_26854_[0], _09097_, _09095_);
  not _40381_ (_09098_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _40382_ (_09099_, _09082_, _09098_);
  and _40383_ (_09100_, _09082_, word_in[1]);
  nor _40384_ (_09102_, _09100_, _09099_);
  nor _40385_ (_09103_, _09102_, _09078_);
  and _40386_ (_09104_, _09078_, word_in[9]);
  or _40387_ (_09105_, _09104_, _09103_);
  and _40388_ (_09106_, _09105_, _09077_);
  and _40389_ (_09107_, _09076_, _08422_);
  or _40390_ (_09108_, _09107_, _09091_);
  or _40391_ (_09109_, _09108_, _09106_);
  or _40392_ (_09111_, _09096_, word_in[25]);
  and _40393_ (_26854_[1], _09111_, _09109_);
  not _40394_ (_09113_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _40395_ (_09115_, _09082_, _09113_);
  and _40396_ (_09116_, _09082_, word_in[2]);
  nor _40397_ (_09117_, _09116_, _09115_);
  nor _40398_ (_09119_, _09117_, _09078_);
  and _40399_ (_09120_, _09078_, word_in[10]);
  or _40400_ (_09121_, _09120_, _09119_);
  and _40401_ (_09122_, _09121_, _09077_);
  and _40402_ (_09123_, _09076_, _08715_);
  or _40403_ (_09124_, _09123_, _09091_);
  or _40404_ (_09125_, _09124_, _09122_);
  or _40405_ (_09126_, _09096_, word_in[26]);
  and _40406_ (_26854_[2], _09126_, _09125_);
  not _40407_ (_09128_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _40408_ (_09129_, _09082_, _09128_);
  and _40409_ (_09130_, _09082_, word_in[3]);
  nor _40410_ (_09131_, _09130_, _09129_);
  nor _40411_ (_09132_, _09131_, _09078_);
  and _40412_ (_09133_, _09078_, word_in[11]);
  or _40413_ (_09134_, _09133_, _09132_);
  and _40414_ (_09135_, _09134_, _09077_);
  and _40415_ (_09136_, _09076_, _08728_);
  or _40416_ (_09137_, _09136_, _09091_);
  or _40417_ (_09138_, _09137_, _09135_);
  or _40418_ (_09139_, _09096_, word_in[27]);
  and _40419_ (_26854_[3], _09139_, _09138_);
  not _40420_ (_09141_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _40421_ (_09142_, _09082_, _09141_);
  and _40422_ (_09143_, _09082_, word_in[4]);
  nor _40423_ (_09144_, _09143_, _09142_);
  nor _40424_ (_09145_, _09144_, _09078_);
  and _40425_ (_09146_, _09078_, word_in[12]);
  or _40426_ (_09147_, _09146_, _09145_);
  and _40427_ (_09148_, _09147_, _09077_);
  and _40428_ (_09149_, _09076_, _08744_);
  or _40429_ (_09150_, _09149_, _09091_);
  or _40430_ (_09151_, _09150_, _09148_);
  or _40431_ (_09152_, _09096_, word_in[28]);
  and _40432_ (_26854_[4], _09152_, _09151_);
  not _40433_ (_09153_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _40434_ (_09154_, _09082_, _09153_);
  and _40435_ (_09155_, _09082_, word_in[5]);
  nor _40436_ (_09157_, _09155_, _09154_);
  nor _40437_ (_09158_, _09157_, _09078_);
  and _40438_ (_09159_, _09078_, word_in[13]);
  or _40439_ (_09160_, _09159_, _09158_);
  and _40440_ (_09161_, _09160_, _09077_);
  and _40441_ (_09162_, _09076_, _08758_);
  or _40442_ (_09163_, _09162_, _09091_);
  or _40443_ (_09164_, _09163_, _09161_);
  or _40444_ (_09165_, _09096_, word_in[29]);
  and _40445_ (_26854_[5], _09165_, _09164_);
  not _40446_ (_09166_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _40447_ (_09168_, _09082_, _09166_);
  and _40448_ (_09169_, _09082_, word_in[6]);
  nor _40449_ (_09170_, _09169_, _09168_);
  nor _40450_ (_09171_, _09170_, _09078_);
  and _40451_ (_09173_, _09078_, word_in[14]);
  or _40452_ (_09175_, _09173_, _09171_);
  and _40453_ (_09176_, _09175_, _09077_);
  and _40454_ (_09177_, _09076_, _08774_);
  or _40455_ (_09178_, _09177_, _09091_);
  or _40456_ (_09180_, _09178_, _09176_);
  or _40457_ (_09181_, _09096_, word_in[30]);
  and _40458_ (_26854_[6], _09181_, _09180_);
  or _40459_ (_09182_, _09077_, _08033_);
  nor _40460_ (_09183_, _09082_, _07689_);
  and _40461_ (_09185_, _09082_, word_in[7]);
  or _40462_ (_09186_, _09185_, _09183_);
  or _40463_ (_09187_, _09186_, _09078_);
  not _40464_ (_09188_, word_in[15]);
  nand _40465_ (_09189_, _09078_, _09188_);
  and _40466_ (_09192_, _09189_, _09187_);
  or _40467_ (_09193_, _09192_, _09076_);
  and _40468_ (_09195_, _09193_, _09182_);
  or _40469_ (_09196_, _09195_, _09091_);
  or _40470_ (_09197_, _09096_, word_in[31]);
  and _40471_ (_26854_[7], _09197_, _09196_);
  and _40472_ (_09198_, _08930_, _07754_);
  and _40473_ (_09199_, _08683_, _07845_);
  not _40474_ (_09200_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _40475_ (_09201_, _08940_, _08688_);
  nor _40476_ (_09203_, _09201_, _09200_);
  and _40477_ (_09204_, _09201_, _08402_);
  or _40478_ (_09205_, _09204_, _09203_);
  or _40479_ (_09207_, _09205_, _09199_);
  not _40480_ (_09208_, _09199_);
  or _40481_ (_09209_, _09208_, word_in[8]);
  and _40482_ (_09210_, _09209_, _09207_);
  and _40483_ (_09211_, _08007_, _07915_);
  and _40484_ (_09212_, _09211_, _07780_);
  or _40485_ (_09213_, _09212_, _09210_);
  not _40486_ (_09214_, _09212_);
  or _40487_ (_09216_, _09214_, _08678_);
  and _40488_ (_09217_, _09216_, _09213_);
  or _40489_ (_09218_, _09217_, _09198_);
  not _40490_ (_09220_, _09198_);
  or _40491_ (_09221_, _09220_, word_in[24]);
  and _40492_ (_26855_[0], _09221_, _09218_);
  not _40493_ (_09222_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _40494_ (_09223_, _09201_, _09222_);
  and _40495_ (_09224_, _09201_, _08428_);
  or _40496_ (_09226_, _09224_, _09223_);
  and _40497_ (_09227_, _09226_, _09208_);
  and _40498_ (_09229_, _09199_, word_in[9]);
  or _40499_ (_09230_, _09229_, _09227_);
  or _40500_ (_09231_, _09230_, _09212_);
  or _40501_ (_09232_, _09214_, _08422_);
  and _40502_ (_09233_, _09232_, _09231_);
  or _40503_ (_09234_, _09233_, _09198_);
  or _40504_ (_09235_, _09220_, word_in[25]);
  and _40505_ (_26855_[1], _09235_, _09234_);
  not _40506_ (_09236_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor _40507_ (_09237_, _09201_, _09236_);
  and _40508_ (_09238_, _09201_, _08591_);
  or _40509_ (_09239_, _09238_, _09237_);
  or _40510_ (_09240_, _09239_, _09199_);
  or _40511_ (_09241_, _09208_, word_in[10]);
  and _40512_ (_09242_, _09241_, _09240_);
  or _40513_ (_09243_, _09242_, _09212_);
  or _40514_ (_09244_, _09214_, _08715_);
  and _40515_ (_09245_, _09244_, _09243_);
  or _40516_ (_09246_, _09245_, _09198_);
  or _40517_ (_09247_, _09220_, word_in[26]);
  and _40518_ (_26855_[2], _09247_, _09246_);
  not _40519_ (_09248_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _40520_ (_09249_, _09201_, _09248_);
  and _40521_ (_09250_, _09201_, _08604_);
  or _40522_ (_09251_, _09250_, _09249_);
  and _40523_ (_09252_, _09251_, _09208_);
  and _40524_ (_09253_, _09199_, word_in[11]);
  or _40525_ (_09255_, _09253_, _09252_);
  or _40526_ (_09256_, _09255_, _09212_);
  or _40527_ (_09257_, _09214_, _08728_);
  and _40528_ (_09259_, _09257_, _09256_);
  or _40529_ (_09260_, _09259_, _09198_);
  or _40530_ (_09261_, _09220_, word_in[27]);
  and _40531_ (_26855_[3], _09261_, _09260_);
  not _40532_ (_09262_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor _40533_ (_09263_, _09201_, _09262_);
  and _40534_ (_09264_, _09201_, _08619_);
  or _40535_ (_09265_, _09264_, _09263_);
  or _40536_ (_09266_, _09265_, _09199_);
  or _40537_ (_09267_, _09208_, word_in[12]);
  and _40538_ (_09268_, _09267_, _09266_);
  or _40539_ (_09269_, _09268_, _09212_);
  or _40540_ (_09271_, _09214_, _08744_);
  and _40541_ (_09272_, _09271_, _09269_);
  or _40542_ (_09273_, _09272_, _09198_);
  or _40543_ (_09275_, _09220_, word_in[28]);
  and _40544_ (_26855_[4], _09275_, _09273_);
  and _40545_ (_09276_, _02345_, _23707_);
  and _40546_ (_09278_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or _40547_ (_02210_, _09278_, _09276_);
  not _40548_ (_09279_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _40549_ (_09280_, _09201_, _09279_);
  and _40550_ (_09281_, _09201_, _08501_);
  or _40551_ (_09283_, _09281_, _09280_);
  or _40552_ (_09284_, _09283_, _09199_);
  or _40553_ (_09285_, _09208_, word_in[13]);
  and _40554_ (_09286_, _09285_, _09284_);
  or _40555_ (_09287_, _09286_, _09212_);
  nor _40556_ (_09288_, _09214_, _08758_);
  nor _40557_ (_09289_, _09288_, _09198_);
  and _40558_ (_09290_, _09289_, _09287_);
  and _40559_ (_09292_, _09198_, word_in[29]);
  or _40560_ (_26855_[5], _09292_, _09290_);
  not _40561_ (_09293_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _40562_ (_09294_, _09201_, _09293_);
  and _40563_ (_09295_, _09201_, _08648_);
  or _40564_ (_09297_, _09295_, _09294_);
  and _40565_ (_09298_, _09297_, _09208_);
  and _40566_ (_09300_, _09199_, word_in[14]);
  or _40567_ (_09301_, _09300_, _09298_);
  or _40568_ (_09303_, _09301_, _09212_);
  nor _40569_ (_09304_, _09214_, _08774_);
  nor _40570_ (_09306_, _09304_, _09198_);
  and _40571_ (_09307_, _09306_, _09303_);
  and _40572_ (_09308_, _09198_, word_in[30]);
  or _40573_ (_26855_[6], _09308_, _09307_);
  nor _40574_ (_09310_, _09201_, _07846_);
  and _40575_ (_09311_, _09201_, _08019_);
  or _40576_ (_09313_, _09311_, _09310_);
  or _40577_ (_09314_, _09313_, _09199_);
  nand _40578_ (_09316_, _09199_, _09188_);
  and _40579_ (_09318_, _09316_, _09314_);
  or _40580_ (_09319_, _09318_, _09212_);
  nor _40581_ (_09320_, _09214_, _08033_);
  nor _40582_ (_09322_, _09320_, _09198_);
  and _40583_ (_09323_, _09322_, _09319_);
  and _40584_ (_09324_, _09198_, word_in[31]);
  or _40585_ (_26855_[7], _09324_, _09323_);
  and _40586_ (_09325_, _08028_, _08073_);
  not _40587_ (_09326_, _09325_);
  and _40588_ (_09328_, _08227_, _08815_);
  and _40589_ (_09329_, _09328_, _08678_);
  not _40590_ (_09330_, _09328_);
  and _40591_ (_09332_, _08011_, _07845_);
  not _40592_ (_09333_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _40593_ (_09335_, _08940_, _08014_);
  nor _40594_ (_09336_, _09335_, _09333_);
  and _40595_ (_09337_, _09335_, word_in[0]);
  nor _40596_ (_09339_, _09337_, _09336_);
  nor _40597_ (_09341_, _09339_, _09332_);
  and _40598_ (_09342_, _09332_, word_in[8]);
  or _40599_ (_09344_, _09342_, _09341_);
  and _40600_ (_09345_, _09344_, _09330_);
  or _40601_ (_09346_, _09345_, _09329_);
  and _40602_ (_09348_, _09346_, _09326_);
  and _40603_ (_09349_, _09325_, word_in[24]);
  or _40604_ (_26856_[0], _09349_, _09348_);
  and _40605_ (_09351_, _09325_, _08973_);
  not _40606_ (_09352_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor _40607_ (_09353_, _09335_, _09352_);
  and _40608_ (_09355_, _09335_, word_in[1]);
  nor _40609_ (_09356_, _09355_, _09353_);
  nor _40610_ (_09358_, _09356_, _09332_);
  and _40611_ (_09360_, _09332_, word_in[9]);
  or _40612_ (_09361_, _09360_, _09358_);
  and _40613_ (_09362_, _09361_, _09330_);
  and _40614_ (_09363_, _09328_, _08422_);
  or _40615_ (_09364_, _09363_, _09362_);
  and _40616_ (_09367_, _09364_, _09326_);
  or _40617_ (_26856_[1], _09367_, _09351_);
  and _40618_ (_09369_, _09328_, _08715_);
  not _40619_ (_09371_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _40620_ (_09372_, _09335_, _09371_);
  and _40621_ (_09374_, _09335_, word_in[2]);
  nor _40622_ (_09376_, _09374_, _09372_);
  nor _40623_ (_09377_, _09376_, _09332_);
  and _40624_ (_09378_, _09332_, word_in[10]);
  or _40625_ (_09380_, _09378_, _09377_);
  and _40626_ (_09381_, _09380_, _09330_);
  or _40627_ (_09383_, _09381_, _09369_);
  and _40628_ (_09385_, _09383_, _09326_);
  and _40629_ (_09386_, _09325_, word_in[26]);
  or _40630_ (_26856_[2], _09386_, _09385_);
  and _40631_ (_09388_, _09328_, _08728_);
  not _40632_ (_09389_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _40633_ (_09390_, _09335_, _09389_);
  and _40634_ (_09391_, _09335_, word_in[3]);
  nor _40635_ (_09392_, _09391_, _09390_);
  nor _40636_ (_09394_, _09392_, _09332_);
  and _40637_ (_09395_, _09332_, word_in[11]);
  or _40638_ (_09396_, _09395_, _09394_);
  and _40639_ (_09397_, _09396_, _09330_);
  or _40640_ (_09398_, _09397_, _09388_);
  and _40641_ (_09399_, _09398_, _09326_);
  and _40642_ (_09400_, _09325_, word_in[27]);
  or _40643_ (_26856_[3], _09400_, _09399_);
  and _40644_ (_09401_, _09328_, _08744_);
  not _40645_ (_09402_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor _40646_ (_09403_, _09335_, _09402_);
  and _40647_ (_09404_, _09335_, word_in[4]);
  nor _40648_ (_09405_, _09404_, _09403_);
  nor _40649_ (_09406_, _09405_, _09332_);
  and _40650_ (_09407_, _09332_, word_in[12]);
  or _40651_ (_09408_, _09407_, _09406_);
  and _40652_ (_09409_, _09408_, _09330_);
  or _40653_ (_09410_, _09409_, _09401_);
  and _40654_ (_09411_, _09410_, _09326_);
  and _40655_ (_09412_, _09325_, word_in[28]);
  or _40656_ (_26856_[4], _09412_, _09411_);
  and _40657_ (_09414_, _09325_, _08495_);
  not _40658_ (_09415_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor _40659_ (_09416_, _09335_, _09415_);
  and _40660_ (_09417_, _09335_, word_in[5]);
  nor _40661_ (_09418_, _09417_, _09416_);
  nor _40662_ (_09419_, _09418_, _09332_);
  and _40663_ (_09420_, _09332_, word_in[13]);
  or _40664_ (_09422_, _09420_, _09419_);
  and _40665_ (_09423_, _09422_, _09330_);
  and _40666_ (_09424_, _09328_, _08758_);
  or _40667_ (_09425_, _09424_, _09423_);
  and _40668_ (_09426_, _09425_, _09326_);
  or _40669_ (_26856_[5], _09426_, _09414_);
  and _40670_ (_09427_, _09328_, _08774_);
  not _40671_ (_09428_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor _40672_ (_09429_, _09335_, _09428_);
  and _40673_ (_09430_, _09335_, word_in[6]);
  nor _40674_ (_09431_, _09430_, _09429_);
  nor _40675_ (_09432_, _09431_, _09332_);
  and _40676_ (_09434_, _09332_, word_in[14]);
  or _40677_ (_09435_, _09434_, _09432_);
  and _40678_ (_09436_, _09435_, _09330_);
  or _40679_ (_09437_, _09436_, _09427_);
  and _40680_ (_09438_, _09437_, _09326_);
  and _40681_ (_09439_, _09325_, word_in[30]);
  or _40682_ (_26856_[6], _09439_, _09438_);
  and _40683_ (_09440_, _09328_, _08033_);
  nor _40684_ (_09441_, _09335_, _07682_);
  and _40685_ (_09442_, _09335_, word_in[7]);
  nor _40686_ (_09443_, _09442_, _09441_);
  nor _40687_ (_09444_, _09443_, _09332_);
  and _40688_ (_09445_, _09332_, word_in[15]);
  or _40689_ (_09446_, _09445_, _09444_);
  and _40690_ (_09447_, _09446_, _09330_);
  or _40691_ (_09448_, _09447_, _09440_);
  and _40692_ (_09449_, _09448_, _09326_);
  and _40693_ (_09450_, _09325_, word_in[31]);
  or _40694_ (_26856_[7], _09450_, _09449_);
  and _40695_ (_09451_, _08006_, _08122_);
  and _40696_ (_09452_, _08010_, _07763_);
  not _40697_ (_09453_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nand _40698_ (_09454_, _07761_, _07577_);
  not _40699_ (_09455_, _09454_);
  and _40700_ (_09456_, _08015_, _09455_);
  and _40701_ (_09457_, _09456_, _08396_);
  nor _40702_ (_09458_, _09457_, _09453_);
  and _40703_ (_09459_, _09457_, _08402_);
  or _40704_ (_09460_, _09459_, _09458_);
  or _40705_ (_09461_, _09460_, _09452_);
  not _40706_ (_09462_, _09452_);
  or _40707_ (_09463_, _09462_, word_in[8]);
  and _40708_ (_09464_, _09463_, _09461_);
  or _40709_ (_09465_, _09464_, _09451_);
  and _40710_ (_09466_, _08028_, _07951_);
  and _40711_ (_09467_, _09466_, _07790_);
  not _40712_ (_09468_, _09451_);
  nor _40713_ (_09469_, _09468_, word_in[16]);
  nor _40714_ (_09470_, _09469_, _09467_);
  and _40715_ (_09471_, _09470_, _09465_);
  and _40716_ (_09472_, _09467_, word_in[24]);
  or _40717_ (_26857_[0], _09472_, _09471_);
  or _40718_ (_09473_, _09468_, word_in[17]);
  not _40719_ (_09474_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _40720_ (_09475_, _09457_, _09474_);
  and _40721_ (_09476_, _09457_, _08428_);
  or _40722_ (_09477_, _09476_, _09475_);
  or _40723_ (_09478_, _09477_, _09452_);
  or _40724_ (_09479_, _09462_, word_in[9]);
  and _40725_ (_09480_, _09479_, _09478_);
  or _40726_ (_09481_, _09480_, _09451_);
  and _40727_ (_09482_, _09481_, _09473_);
  or _40728_ (_09483_, _09482_, _09467_);
  not _40729_ (_09484_, _09467_);
  or _40730_ (_09485_, _09484_, word_in[25]);
  and _40731_ (_26857_[1], _09485_, _09483_);
  not _40732_ (_09486_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _40733_ (_09487_, _09457_, _09486_);
  and _40734_ (_09488_, _09457_, word_in[2]);
  or _40735_ (_09489_, _09488_, _09487_);
  and _40736_ (_09491_, _09489_, _09462_);
  and _40737_ (_09492_, _09452_, word_in[10]);
  or _40738_ (_09493_, _09492_, _09491_);
  and _40739_ (_09494_, _09493_, _09468_);
  and _40740_ (_09495_, _09451_, word_in[18]);
  or _40741_ (_09496_, _09495_, _09494_);
  and _40742_ (_09497_, _09496_, _09484_);
  and _40743_ (_09498_, _09467_, word_in[26]);
  or _40744_ (_26857_[2], _09498_, _09497_);
  not _40745_ (_09499_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _40746_ (_09500_, _09457_, _09499_);
  and _40747_ (_09501_, _09457_, _08604_);
  or _40748_ (_09502_, _09501_, _09500_);
  or _40749_ (_09503_, _09502_, _09452_);
  or _40750_ (_09504_, _09462_, word_in[11]);
  and _40751_ (_09505_, _09504_, _09468_);
  and _40752_ (_09506_, _09505_, _09503_);
  and _40753_ (_09507_, _09451_, word_in[19]);
  or _40754_ (_09508_, _09507_, _09506_);
  or _40755_ (_09509_, _09508_, _09467_);
  or _40756_ (_09510_, _09484_, word_in[27]);
  and _40757_ (_26857_[3], _09510_, _09509_);
  or _40758_ (_09511_, _09468_, word_in[20]);
  not _40759_ (_09512_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _40760_ (_09513_, _09457_, _09512_);
  and _40761_ (_09514_, _09457_, _08619_);
  or _40762_ (_09515_, _09514_, _09513_);
  or _40763_ (_09516_, _09515_, _09452_);
  or _40764_ (_09517_, _09462_, word_in[12]);
  and _40765_ (_09518_, _09517_, _09516_);
  or _40766_ (_09520_, _09518_, _09451_);
  and _40767_ (_09521_, _09520_, _09511_);
  or _40768_ (_09522_, _09521_, _09467_);
  or _40769_ (_09524_, _09484_, word_in[28]);
  and _40770_ (_26857_[4], _09524_, _09522_);
  not _40771_ (_09525_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _40772_ (_09526_, _09457_, _09525_);
  and _40773_ (_09527_, _09457_, _08501_);
  or _40774_ (_09528_, _09527_, _09526_);
  or _40775_ (_09529_, _09528_, _09452_);
  or _40776_ (_09530_, _09462_, word_in[13]);
  and _40777_ (_09531_, _09530_, _09529_);
  or _40778_ (_09532_, _09531_, _09451_);
  or _40779_ (_09533_, _09468_, word_in[21]);
  and _40780_ (_09534_, _09533_, _09532_);
  or _40781_ (_09535_, _09534_, _09467_);
  or _40782_ (_09536_, _09484_, word_in[29]);
  and _40783_ (_26857_[5], _09536_, _09535_);
  not _40784_ (_09537_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _40785_ (_09538_, _09457_, _09537_);
  and _40786_ (_09539_, _09457_, _08648_);
  or _40787_ (_09540_, _09539_, _09538_);
  or _40788_ (_09541_, _09540_, _09452_);
  or _40789_ (_09542_, _09462_, word_in[14]);
  and _40790_ (_09543_, _09542_, _09541_);
  or _40791_ (_09544_, _09543_, _09451_);
  nor _40792_ (_09545_, _09468_, word_in[22]);
  nor _40793_ (_09546_, _09545_, _09467_);
  and _40794_ (_09547_, _09546_, _09544_);
  and _40795_ (_09548_, _09467_, word_in[30]);
  or _40796_ (_26857_[6], _09548_, _09547_);
  nor _40797_ (_09549_, _09457_, _07819_);
  and _40798_ (_09550_, _09457_, word_in[7]);
  or _40799_ (_09551_, _09550_, _09549_);
  and _40800_ (_09552_, _09551_, _09462_);
  and _40801_ (_09553_, _09452_, word_in[15]);
  or _40802_ (_09554_, _09553_, _09552_);
  or _40803_ (_09555_, _09554_, _09451_);
  nor _40804_ (_09556_, _09468_, word_in[23]);
  nor _40805_ (_09557_, _09556_, _09467_);
  and _40806_ (_09558_, _09557_, _09555_);
  and _40807_ (_09559_, _09467_, word_in[31]);
  or _40808_ (_26857_[7], _09559_, _09558_);
  nor _40809_ (_26860_[7], _24508_, rst);
  and _40810_ (_09560_, _08799_, _23747_);
  and _40811_ (_09561_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  or _40812_ (_02338_, _09561_, _09560_);
  and _40813_ (_09562_, _24371_, _23898_);
  and _40814_ (_09563_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or _40815_ (_27197_, _09563_, _09562_);
  nor _40816_ (_26887_[7], _26770_, rst);
  and _40817_ (_09564_, _08799_, _23824_);
  and _40818_ (_09565_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  or _40819_ (_02348_, _09565_, _09564_);
  nor _40820_ (_26860_[5], _24530_, rst);
  and _40821_ (_09566_, _08043_, _23898_);
  and _40822_ (_09567_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or _40823_ (_02362_, _09567_, _09566_);
  and _40824_ (_09568_, _08563_, _07887_);
  and _40825_ (_09569_, _08553_, _07770_);
  not _40826_ (_09570_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _40827_ (_09571_, _09456_, _08557_);
  nor _40828_ (_09572_, _09571_, _09570_);
  and _40829_ (_09573_, _09571_, _08402_);
  or _40830_ (_09574_, _09573_, _09572_);
  or _40831_ (_09575_, _09574_, _09569_);
  not _40832_ (_09576_, _09569_);
  or _40833_ (_09577_, _09576_, word_in[8]);
  and _40834_ (_09578_, _09577_, _09575_);
  or _40835_ (_09579_, _09578_, _09568_);
  and _40836_ (_09580_, _09466_, _07751_);
  not _40837_ (_09581_, _09568_);
  nor _40838_ (_09582_, _09581_, _08678_);
  nor _40839_ (_09583_, _09582_, _09580_);
  and _40840_ (_09584_, _09583_, _09579_);
  and _40841_ (_09585_, _09580_, word_in[24]);
  or _40842_ (_26858_[0], _09585_, _09584_);
  not _40843_ (_09586_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _40844_ (_09587_, _09571_, _09586_);
  and _40845_ (_09588_, _09571_, _08428_);
  or _40846_ (_09589_, _09588_, _09587_);
  or _40847_ (_09590_, _09589_, _09569_);
  or _40848_ (_09591_, _09576_, word_in[9]);
  and _40849_ (_09592_, _09591_, _09590_);
  or _40850_ (_09593_, _09592_, _09568_);
  nor _40851_ (_09594_, _09581_, _08422_);
  nor _40852_ (_09595_, _09594_, _09580_);
  and _40853_ (_09596_, _09595_, _09593_);
  and _40854_ (_09597_, _09580_, word_in[25]);
  or _40855_ (_26858_[1], _09597_, _09596_);
  not _40856_ (_09598_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _40857_ (_09599_, _09571_, _09598_);
  and _40858_ (_09601_, _09571_, _08591_);
  or _40859_ (_09602_, _09601_, _09599_);
  or _40860_ (_09603_, _09602_, _09569_);
  or _40861_ (_09604_, _09576_, word_in[10]);
  and _40862_ (_09605_, _09604_, _09603_);
  or _40863_ (_09606_, _09605_, _09568_);
  nor _40864_ (_09607_, _09581_, _08715_);
  nor _40865_ (_09608_, _09607_, _09580_);
  and _40866_ (_09610_, _09608_, _09606_);
  and _40867_ (_09611_, _09580_, word_in[26]);
  or _40868_ (_26858_[2], _09611_, _09610_);
  not _40869_ (_09613_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _40870_ (_09614_, _09571_, _09613_);
  and _40871_ (_09615_, _09571_, _08604_);
  or _40872_ (_09616_, _09615_, _09614_);
  or _40873_ (_09617_, _09616_, _09569_);
  or _40874_ (_09618_, _09576_, word_in[11]);
  and _40875_ (_09619_, _09618_, _09617_);
  or _40876_ (_09620_, _09619_, _09568_);
  nor _40877_ (_09621_, _09581_, _08728_);
  nor _40878_ (_09622_, _09621_, _09580_);
  and _40879_ (_09623_, _09622_, _09620_);
  and _40880_ (_09624_, _09580_, word_in[27]);
  or _40881_ (_26858_[3], _09624_, _09623_);
  not _40882_ (_09625_, _09580_);
  not _40883_ (_09627_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _40884_ (_09628_, _09571_, _09627_);
  and _40885_ (_09629_, _09571_, _08619_);
  nor _40886_ (_09630_, _09629_, _09628_);
  nor _40887_ (_09631_, _09630_, _09569_);
  and _40888_ (_09632_, _09569_, word_in[12]);
  or _40889_ (_09633_, _09632_, _09568_);
  or _40890_ (_09634_, _09633_, _09631_);
  or _40891_ (_09635_, _09581_, _08744_);
  and _40892_ (_09636_, _09635_, _09634_);
  and _40893_ (_09637_, _09636_, _09625_);
  and _40894_ (_09639_, _09580_, word_in[28]);
  or _40895_ (_26858_[4], _09639_, _09637_);
  or _40896_ (_09640_, _09581_, _08758_);
  not _40897_ (_09641_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _40898_ (_09642_, _09571_, _09641_);
  and _40899_ (_09643_, _09571_, _08501_);
  nor _40900_ (_09644_, _09643_, _09642_);
  nor _40901_ (_09645_, _09644_, _09569_);
  and _40902_ (_09646_, _09569_, word_in[13]);
  or _40903_ (_09647_, _09646_, _09568_);
  or _40904_ (_09648_, _09647_, _09645_);
  and _40905_ (_09649_, _09648_, _09640_);
  and _40906_ (_09651_, _09649_, _09625_);
  and _40907_ (_09653_, _09580_, word_in[29]);
  or _40908_ (_26858_[5], _09653_, _09651_);
  not _40909_ (_09654_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _40910_ (_09655_, _09571_, _09654_);
  and _40911_ (_09656_, _09571_, _08648_);
  or _40912_ (_09657_, _09656_, _09655_);
  or _40913_ (_09658_, _09657_, _09569_);
  or _40914_ (_09659_, _09576_, word_in[14]);
  and _40915_ (_09660_, _09659_, _09658_);
  or _40916_ (_09661_, _09660_, _09568_);
  nor _40917_ (_09662_, _09581_, _08774_);
  nor _40918_ (_09663_, _09662_, _09580_);
  and _40919_ (_09664_, _09663_, _09661_);
  and _40920_ (_09665_, _09580_, word_in[30]);
  or _40921_ (_26858_[6], _09665_, _09664_);
  nor _40922_ (_09666_, _09571_, _07709_);
  and _40923_ (_09667_, _09571_, _08019_);
  or _40924_ (_09669_, _09667_, _09666_);
  or _40925_ (_09670_, _09669_, _09569_);
  nand _40926_ (_09671_, _09569_, _09188_);
  and _40927_ (_09672_, _09671_, _09670_);
  or _40928_ (_09673_, _09672_, _09568_);
  nor _40929_ (_09674_, _09581_, _08033_);
  nor _40930_ (_09675_, _09674_, _09580_);
  and _40931_ (_09676_, _09675_, _09673_);
  and _40932_ (_09677_, _09580_, word_in[31]);
  or _40933_ (_26858_[7], _09677_, _09676_);
  and _40934_ (_09678_, _24371_, _23778_);
  and _40935_ (_09679_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or _40936_ (_27196_, _09679_, _09678_);
  and _40937_ (_09682_, _09466_, _07754_);
  and _40938_ (_09683_, _08679_, _07887_);
  not _40939_ (_09684_, _09683_);
  or _40940_ (_09685_, _09684_, _08678_);
  not _40941_ (_09686_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _40942_ (_09687_, _08688_, _09455_);
  nor _40943_ (_09688_, _09687_, _09686_);
  and _40944_ (_09689_, _09687_, _08402_);
  or _40945_ (_09690_, _09689_, _09688_);
  and _40946_ (_09691_, _08010_, _07770_);
  and _40947_ (_09692_, _09691_, _08683_);
  not _40948_ (_09693_, _09692_);
  and _40949_ (_09694_, _09693_, _09690_);
  and _40950_ (_09695_, _08683_, _07770_);
  and _40951_ (_09696_, _09695_, word_in[8]);
  or _40952_ (_09697_, _09696_, _09683_);
  or _40953_ (_09698_, _09697_, _09694_);
  and _40954_ (_09699_, _09698_, _09685_);
  or _40955_ (_09700_, _09699_, _09682_);
  not _40956_ (_09701_, _09682_);
  or _40957_ (_09702_, _09701_, word_in[24]);
  and _40958_ (_26844_[0], _09702_, _09700_);
  not _40959_ (_09703_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _40960_ (_09704_, _09687_, _09703_);
  and _40961_ (_09705_, _09687_, _08428_);
  or _40962_ (_09706_, _09705_, _09704_);
  or _40963_ (_09707_, _09706_, _09695_);
  not _40964_ (_09708_, _09695_);
  or _40965_ (_09709_, _09708_, word_in[9]);
  and _40966_ (_09710_, _09709_, _09707_);
  or _40967_ (_09711_, _09710_, _09683_);
  nor _40968_ (_09712_, _09684_, _08422_);
  nor _40969_ (_09713_, _09712_, _09682_);
  and _40970_ (_09714_, _09713_, _09711_);
  and _40971_ (_09715_, _09682_, word_in[25]);
  or _40972_ (_26844_[1], _09715_, _09714_);
  not _40973_ (_09716_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _40974_ (_09717_, _09687_, _09716_);
  and _40975_ (_09718_, _09687_, _08591_);
  or _40976_ (_09719_, _09718_, _09717_);
  or _40977_ (_09720_, _09719_, _09695_);
  or _40978_ (_09721_, _09708_, word_in[10]);
  and _40979_ (_09722_, _09721_, _09720_);
  or _40980_ (_09723_, _09722_, _09683_);
  nor _40981_ (_09724_, _09684_, _08715_);
  nor _40982_ (_09725_, _09724_, _09682_);
  and _40983_ (_09726_, _09725_, _09723_);
  and _40984_ (_09727_, _09682_, word_in[26]);
  or _40985_ (_26844_[2], _09727_, _09726_);
  and _40986_ (_09729_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and _40987_ (_09730_, _08351_, _24050_);
  or _40988_ (_02446_, _09730_, _09729_);
  not _40989_ (_09732_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _40990_ (_09734_, _09687_, _09732_);
  and _40991_ (_09735_, _09687_, _08604_);
  or _40992_ (_09736_, _09735_, _09734_);
  or _40993_ (_09738_, _09736_, _09695_);
  or _40994_ (_09739_, _09708_, word_in[11]);
  and _40995_ (_09740_, _09739_, _09738_);
  or _40996_ (_09741_, _09740_, _09683_);
  nor _40997_ (_09742_, _09684_, _08728_);
  nor _40998_ (_09743_, _09742_, _09682_);
  and _40999_ (_09744_, _09743_, _09741_);
  and _41000_ (_09745_, _09682_, word_in[27]);
  or _41001_ (_26844_[3], _09745_, _09744_);
  not _41002_ (_09746_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor _41003_ (_09747_, _09687_, _09746_);
  and _41004_ (_09748_, _09687_, _08619_);
  or _41005_ (_09749_, _09748_, _09747_);
  or _41006_ (_09751_, _09749_, _09695_);
  or _41007_ (_09752_, _09708_, word_in[12]);
  and _41008_ (_09754_, _09752_, _09751_);
  or _41009_ (_09755_, _09754_, _09683_);
  nor _41010_ (_09756_, _09684_, _08744_);
  nor _41011_ (_09757_, _09756_, _09682_);
  and _41012_ (_09758_, _09757_, _09755_);
  and _41013_ (_09759_, _09682_, word_in[28]);
  or _41014_ (_26844_[4], _09759_, _09758_);
  not _41015_ (_09760_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _41016_ (_09761_, _09687_, _09760_);
  and _41017_ (_09762_, _09687_, _08501_);
  or _41018_ (_09763_, _09762_, _09761_);
  or _41019_ (_09764_, _09763_, _09695_);
  or _41020_ (_09765_, _09708_, word_in[13]);
  and _41021_ (_09766_, _09765_, _09764_);
  or _41022_ (_09767_, _09766_, _09683_);
  nor _41023_ (_09768_, _09684_, _08758_);
  nor _41024_ (_09770_, _09768_, _09682_);
  and _41025_ (_09771_, _09770_, _09767_);
  and _41026_ (_09773_, _09682_, word_in[29]);
  or _41027_ (_26844_[5], _09773_, _09771_);
  not _41028_ (_09774_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _41029_ (_09775_, _09687_, _09774_);
  and _41030_ (_09776_, _09687_, _08648_);
  or _41031_ (_09777_, _09776_, _09775_);
  or _41032_ (_09778_, _09777_, _09695_);
  or _41033_ (_09779_, _09708_, word_in[14]);
  and _41034_ (_09780_, _09779_, _09778_);
  or _41035_ (_09781_, _09780_, _09683_);
  nor _41036_ (_09782_, _09684_, _08774_);
  nor _41037_ (_09783_, _09782_, _09682_);
  and _41038_ (_09784_, _09783_, _09781_);
  and _41039_ (_09785_, _09682_, word_in[30]);
  or _41040_ (_26844_[6], _09785_, _09784_);
  or _41041_ (_09786_, _09684_, _08033_);
  nor _41042_ (_09787_, _09687_, _07813_);
  and _41043_ (_09788_, _09687_, _08019_);
  or _41044_ (_09789_, _09788_, _09787_);
  and _41045_ (_09790_, _09789_, _09693_);
  and _41046_ (_09792_, _09695_, word_in[15]);
  or _41047_ (_09793_, _09792_, _09683_);
  or _41048_ (_09794_, _09793_, _09790_);
  and _41049_ (_09795_, _09794_, _09786_);
  or _41050_ (_09796_, _09795_, _09682_);
  or _41051_ (_09797_, _09701_, word_in[31]);
  and _41052_ (_26844_[7], _09797_, _09796_);
  and _41053_ (_09798_, _08043_, _23778_);
  and _41054_ (_09799_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or _41055_ (_27210_, _09799_, _09798_);
  and _41056_ (_09800_, _09466_, _07780_);
  and _41057_ (_09801_, _08011_, _07770_);
  not _41058_ (_09802_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _41059_ (_09803_, _09456_, _08014_);
  nor _41060_ (_09804_, _09803_, _09802_);
  and _41061_ (_09805_, _09803_, _08402_);
  nor _41062_ (_09806_, _09805_, _09804_);
  nor _41063_ (_09807_, _09806_, _09801_);
  and _41064_ (_09808_, _08815_, _07887_);
  and _41065_ (_09809_, _09801_, word_in[8]);
  or _41066_ (_09810_, _09809_, _09808_);
  or _41067_ (_09811_, _09810_, _09807_);
  not _41068_ (_09812_, _09808_);
  or _41069_ (_09813_, _09812_, _08678_);
  and _41070_ (_09814_, _09813_, _09811_);
  or _41071_ (_09815_, _09814_, _09800_);
  not _41072_ (_09816_, _09800_);
  or _41073_ (_09817_, _09816_, word_in[24]);
  and _41074_ (_26845_[0], _09817_, _09815_);
  not _41075_ (_09819_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _41076_ (_09820_, _09803_, _09819_);
  and _41077_ (_09822_, _09803_, _08428_);
  or _41078_ (_09824_, _09822_, _09820_);
  or _41079_ (_09825_, _09824_, _09801_);
  not _41080_ (_09826_, _09801_);
  or _41081_ (_09827_, _09826_, word_in[9]);
  and _41082_ (_09828_, _09827_, _09825_);
  or _41083_ (_09829_, _09828_, _09808_);
  nor _41084_ (_09830_, _09812_, _08422_);
  nor _41085_ (_09831_, _09830_, _09800_);
  and _41086_ (_09832_, _09831_, _09829_);
  and _41087_ (_09833_, _09800_, _08973_);
  or _41088_ (_26845_[1], _09833_, _09832_);
  not _41089_ (_09834_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _41090_ (_09835_, _09803_, _09834_);
  and _41091_ (_09836_, _09803_, _08591_);
  nor _41092_ (_09838_, _09836_, _09835_);
  nor _41093_ (_09840_, _09838_, _09801_);
  and _41094_ (_09841_, _09801_, word_in[10]);
  or _41095_ (_09842_, _09841_, _09808_);
  or _41096_ (_09844_, _09842_, _09840_);
  or _41097_ (_09845_, _09812_, _08715_);
  and _41098_ (_09846_, _09845_, _09844_);
  and _41099_ (_09847_, _09846_, _09816_);
  and _41100_ (_09848_, _09800_, word_in[26]);
  or _41101_ (_26845_[2], _09848_, _09847_);
  not _41102_ (_09849_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _41103_ (_09850_, _09803_, _09849_);
  and _41104_ (_09851_, _09803_, _08604_);
  nor _41105_ (_09852_, _09851_, _09850_);
  nor _41106_ (_09853_, _09852_, _09801_);
  and _41107_ (_09855_, _09801_, word_in[11]);
  or _41108_ (_09856_, _09855_, _09808_);
  or _41109_ (_09857_, _09856_, _09853_);
  or _41110_ (_09858_, _09812_, _08728_);
  and _41111_ (_09859_, _09858_, _09857_);
  and _41112_ (_09861_, _09859_, _09816_);
  and _41113_ (_09862_, _09800_, word_in[27]);
  or _41114_ (_26845_[3], _09862_, _09861_);
  not _41115_ (_09863_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _41116_ (_09864_, _09803_, _09863_);
  and _41117_ (_09865_, _09803_, _08619_);
  nor _41118_ (_09866_, _09865_, _09864_);
  nor _41119_ (_09867_, _09866_, _09801_);
  and _41120_ (_09868_, _09801_, word_in[12]);
  or _41121_ (_09869_, _09868_, _09808_);
  or _41122_ (_09870_, _09869_, _09867_);
  or _41123_ (_09871_, _09812_, _08744_);
  and _41124_ (_09872_, _09871_, _09870_);
  or _41125_ (_09873_, _09872_, _09800_);
  or _41126_ (_09874_, _09816_, word_in[28]);
  and _41127_ (_26845_[4], _09874_, _09873_);
  not _41128_ (_09875_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _41129_ (_09876_, _09803_, _09875_);
  and _41130_ (_09877_, _09803_, _08501_);
  or _41131_ (_09878_, _09877_, _09876_);
  or _41132_ (_09879_, _09878_, _09801_);
  or _41133_ (_09880_, _09826_, word_in[13]);
  and _41134_ (_09881_, _09880_, _09879_);
  or _41135_ (_09882_, _09881_, _09808_);
  nor _41136_ (_09883_, _09812_, _08758_);
  nor _41137_ (_09884_, _09883_, _09800_);
  and _41138_ (_09885_, _09884_, _09882_);
  and _41139_ (_09886_, _09800_, _08495_);
  or _41140_ (_26845_[5], _09886_, _09885_);
  not _41141_ (_09888_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _41142_ (_09889_, _09803_, _09888_);
  and _41143_ (_09890_, _09803_, _08648_);
  nor _41144_ (_09891_, _09890_, _09889_);
  nor _41145_ (_09892_, _09891_, _09801_);
  and _41146_ (_09893_, _09801_, word_in[14]);
  or _41147_ (_09894_, _09893_, _09808_);
  or _41148_ (_09895_, _09894_, _09892_);
  or _41149_ (_09896_, _09812_, _08774_);
  and _41150_ (_09897_, _09896_, _09895_);
  and _41151_ (_09898_, _09897_, _09816_);
  and _41152_ (_09899_, _09800_, word_in[30]);
  or _41153_ (_26845_[6], _09899_, _09898_);
  nor _41154_ (_09901_, _09803_, _07731_);
  and _41155_ (_09902_, _09803_, _08019_);
  or _41156_ (_09903_, _09902_, _09901_);
  or _41157_ (_09904_, _09903_, _09801_);
  nand _41158_ (_09905_, _09801_, _09188_);
  and _41159_ (_09907_, _09905_, _09904_);
  or _41160_ (_09908_, _09907_, _09808_);
  nor _41161_ (_09909_, _09812_, _08033_);
  nor _41162_ (_09910_, _09909_, _09800_);
  and _41163_ (_09911_, _09910_, _09908_);
  and _41164_ (_09912_, _09800_, _09072_);
  or _41165_ (_26845_[7], _09912_, _09911_);
  and _41166_ (_09913_, _24275_, _23754_);
  and _41167_ (_09914_, _09913_, _23747_);
  not _41168_ (_09915_, _09913_);
  and _41169_ (_09916_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or _41170_ (_02539_, _09916_, _09914_);
  and _41171_ (_09917_, _26112_, _26110_);
  nor _41172_ (_09918_, _09917_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _41173_ (_09920_, _09917_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _41174_ (_09921_, _09920_, _09918_);
  and _41175_ (_09922_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _41176_ (_09924_, _09922_, _26118_);
  nor _41177_ (_09925_, _09924_, _09921_);
  nor _41178_ (_09926_, _09925_, _24299_);
  and _41179_ (_09927_, _24299_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _41180_ (_09928_, _09927_, _09926_);
  and _41181_ (_09929_, _09928_, _24294_);
  and _41182_ (_09930_, _24293_, _23816_);
  or _41183_ (_09931_, _09930_, _09929_);
  and _41184_ (_02555_, _09931_, _22762_);
  and _41185_ (_09932_, _24371_, _23747_);
  and _41186_ (_09933_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or _41187_ (_02571_, _09933_, _09932_);
  not _41188_ (_09934_, _07948_);
  and _41189_ (_09935_, _08929_, _09934_);
  and _41190_ (_09936_, _09935_, _07790_);
  not _41191_ (_09937_, _09936_);
  and _41192_ (_09938_, _08008_, _07751_);
  not _41193_ (_09939_, _09938_);
  and _41194_ (_09941_, _08010_, _08244_);
  not _41195_ (_09942_, _09941_);
  and _41196_ (_09943_, _08396_, _08016_);
  and _41197_ (_09944_, _09943_, word_in[0]);
  not _41198_ (_09946_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _41199_ (_09947_, _09943_, _09946_);
  or _41200_ (_09948_, _09947_, _09944_);
  and _41201_ (_09949_, _09948_, _09942_);
  and _41202_ (_09951_, _09941_, word_in[8]);
  or _41203_ (_09953_, _09951_, _09949_);
  and _41204_ (_09955_, _09953_, _09939_);
  and _41205_ (_09957_, _09938_, _08678_);
  or _41206_ (_09959_, _09957_, _09955_);
  and _41207_ (_09960_, _09959_, _09937_);
  and _41208_ (_09961_, _09936_, _08954_);
  or _41209_ (_26846_[0], _09961_, _09960_);
  or _41210_ (_09962_, _09939_, _08422_);
  not _41211_ (_09963_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _41212_ (_09965_, _09943_, _09963_);
  and _41213_ (_09967_, _09943_, _08428_);
  or _41214_ (_09968_, _09967_, _09965_);
  or _41215_ (_09969_, _09968_, _09941_);
  or _41216_ (_09970_, _09942_, word_in[9]);
  and _41217_ (_09971_, _09970_, _09969_);
  or _41218_ (_09972_, _09971_, _09938_);
  and _41219_ (_09973_, _09972_, _09962_);
  or _41220_ (_09975_, _09973_, _09936_);
  or _41221_ (_09977_, _09937_, _08973_);
  and _41222_ (_26846_[1], _09977_, _09975_);
  or _41223_ (_09978_, _09939_, _08715_);
  not _41224_ (_09979_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _41225_ (_09980_, _09943_, _09979_);
  and _41226_ (_09982_, _09943_, _08591_);
  or _41227_ (_09983_, _09982_, _09980_);
  or _41228_ (_09984_, _09983_, _09941_);
  or _41229_ (_09985_, _09942_, word_in[10]);
  and _41230_ (_09986_, _09985_, _09984_);
  or _41231_ (_09987_, _09986_, _09938_);
  and _41232_ (_09989_, _09987_, _09978_);
  or _41233_ (_09990_, _09989_, _09936_);
  or _41234_ (_09992_, _09937_, _08993_);
  and _41235_ (_26846_[2], _09992_, _09990_);
  or _41236_ (_09993_, _09939_, _08728_);
  not _41237_ (_09994_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _41238_ (_09995_, _09943_, _09994_);
  and _41239_ (_09996_, _09943_, _08604_);
  or _41240_ (_09997_, _09996_, _09995_);
  or _41241_ (_09998_, _09997_, _09941_);
  or _41242_ (_09999_, _09942_, word_in[11]);
  and _41243_ (_10000_, _09999_, _09998_);
  or _41244_ (_10001_, _10000_, _09938_);
  and _41245_ (_10002_, _10001_, _09993_);
  or _41246_ (_10003_, _10002_, _09936_);
  or _41247_ (_10004_, _09937_, _08461_);
  and _41248_ (_26846_[3], _10004_, _10003_);
  or _41249_ (_10006_, _09939_, _08744_);
  not _41250_ (_10008_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _41251_ (_10009_, _09943_, _10008_);
  and _41252_ (_10010_, _09943_, _08619_);
  or _41253_ (_10011_, _10010_, _10009_);
  or _41254_ (_10012_, _10011_, _09941_);
  or _41255_ (_10014_, _09942_, word_in[12]);
  and _41256_ (_10016_, _10014_, _10012_);
  or _41257_ (_10017_, _10016_, _09938_);
  and _41258_ (_10018_, _10017_, _10006_);
  or _41259_ (_10019_, _10018_, _09936_);
  or _41260_ (_10020_, _09937_, _08481_);
  and _41261_ (_26846_[4], _10020_, _10019_);
  or _41262_ (_10022_, _09939_, _08758_);
  not _41263_ (_10023_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _41264_ (_10024_, _09943_, _10023_);
  and _41265_ (_10025_, _09943_, _08501_);
  or _41266_ (_10026_, _10025_, _10024_);
  or _41267_ (_10027_, _10026_, _09941_);
  or _41268_ (_10028_, _09942_, word_in[13]);
  and _41269_ (_10029_, _10028_, _10027_);
  or _41270_ (_10030_, _10029_, _09938_);
  and _41271_ (_10031_, _10030_, _10022_);
  or _41272_ (_10032_, _10031_, _09936_);
  or _41273_ (_10033_, _09937_, _08495_);
  and _41274_ (_26846_[5], _10033_, _10032_);
  or _41275_ (_10034_, _09939_, _08774_);
  not _41276_ (_10035_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _41277_ (_10037_, _09943_, _10035_);
  and _41278_ (_10038_, _09943_, _08648_);
  or _41279_ (_10040_, _10038_, _10037_);
  or _41280_ (_10041_, _10040_, _09941_);
  or _41281_ (_10042_, _09942_, word_in[14]);
  and _41282_ (_10043_, _10042_, _10041_);
  or _41283_ (_10044_, _10043_, _09938_);
  and _41284_ (_10045_, _10044_, _10034_);
  or _41285_ (_10046_, _10045_, _09936_);
  or _41286_ (_10047_, _09937_, _08510_);
  and _41287_ (_26846_[6], _10047_, _10046_);
  or _41288_ (_10049_, _09939_, _08033_);
  nor _41289_ (_10051_, _09943_, _07866_);
  and _41290_ (_10052_, _09943_, _08019_);
  or _41291_ (_10053_, _10052_, _10051_);
  or _41292_ (_10054_, _10053_, _09941_);
  nand _41293_ (_10056_, _09941_, _09188_);
  and _41294_ (_10057_, _10056_, _10054_);
  or _41295_ (_10058_, _10057_, _09938_);
  and _41296_ (_10059_, _10058_, _10049_);
  or _41297_ (_10060_, _10059_, _09936_);
  or _41298_ (_10061_, _09937_, _09072_);
  and _41299_ (_26846_[7], _10061_, _10060_);
  and _41300_ (_10062_, _05042_, _23824_);
  and _41301_ (_10063_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or _41302_ (_27135_, _10063_, _10062_);
  and _41303_ (_10064_, _08008_, _07754_);
  not _41304_ (_10065_, _10064_);
  and _41305_ (_10066_, _08553_, _07860_);
  and _41306_ (_10067_, _08557_, _08016_);
  and _41307_ (_10068_, _10067_, word_in[0]);
  not _41308_ (_10069_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _41309_ (_10070_, _10067_, _10069_);
  nor _41310_ (_10071_, _10070_, _10068_);
  nor _41311_ (_10072_, _10071_, _10066_);
  and _41312_ (_10073_, _10066_, word_in[8]);
  or _41313_ (_10075_, _10073_, _10072_);
  and _41314_ (_10076_, _10075_, _10065_);
  and _41315_ (_10077_, _09935_, _07751_);
  and _41316_ (_10078_, _10064_, _08678_);
  or _41317_ (_10079_, _10078_, _10077_);
  or _41318_ (_10080_, _10079_, _10076_);
  not _41319_ (_10081_, _10077_);
  or _41320_ (_10082_, _10081_, word_in[24]);
  and _41321_ (_26847_[0], _10082_, _10080_);
  not _41322_ (_10084_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _41323_ (_10086_, _10067_, _10084_);
  and _41324_ (_10087_, _10067_, word_in[1]);
  or _41325_ (_10088_, _10087_, _10086_);
  or _41326_ (_10090_, _10088_, _10066_);
  not _41327_ (_10091_, _10066_);
  or _41328_ (_10092_, _10091_, word_in[9]);
  and _41329_ (_10093_, _10092_, _10090_);
  or _41330_ (_10094_, _10093_, _10064_);
  or _41331_ (_10095_, _10065_, _08422_);
  and _41332_ (_10096_, _10095_, _10094_);
  and _41333_ (_10098_, _10096_, _10081_);
  and _41334_ (_10099_, _10077_, word_in[25]);
  or _41335_ (_26847_[1], _10099_, _10098_);
  or _41336_ (_10101_, _10065_, _08715_);
  not _41337_ (_10102_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _41338_ (_10103_, _10067_, _10102_);
  and _41339_ (_10105_, _10067_, word_in[2]);
  or _41340_ (_10106_, _10105_, _10103_);
  or _41341_ (_10107_, _10106_, _10066_);
  or _41342_ (_10109_, _10091_, word_in[10]);
  and _41343_ (_10111_, _10109_, _10107_);
  or _41344_ (_10112_, _10111_, _10064_);
  and _41345_ (_10113_, _10112_, _10101_);
  or _41346_ (_10115_, _10113_, _10077_);
  or _41347_ (_10116_, _10081_, word_in[26]);
  and _41348_ (_26847_[2], _10116_, _10115_);
  or _41349_ (_10117_, _10065_, _08728_);
  not _41350_ (_10118_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _41351_ (_10119_, _10067_, _10118_);
  and _41352_ (_10120_, _10067_, word_in[3]);
  or _41353_ (_10121_, _10120_, _10119_);
  or _41354_ (_10122_, _10121_, _10066_);
  or _41355_ (_10123_, _10091_, word_in[11]);
  and _41356_ (_10124_, _10123_, _10122_);
  or _41357_ (_10126_, _10124_, _10064_);
  and _41358_ (_10127_, _10126_, _10117_);
  and _41359_ (_10129_, _10127_, _10081_);
  and _41360_ (_10131_, _10077_, word_in[27]);
  or _41361_ (_26847_[3], _10131_, _10129_);
  or _41362_ (_10134_, _10065_, _08744_);
  not _41363_ (_10135_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _41364_ (_10136_, _10067_, _10135_);
  and _41365_ (_10137_, _10067_, word_in[4]);
  or _41366_ (_10139_, _10137_, _10136_);
  or _41367_ (_10140_, _10139_, _10066_);
  or _41368_ (_10141_, _10091_, word_in[12]);
  and _41369_ (_10142_, _10141_, _10140_);
  or _41370_ (_10144_, _10142_, _10064_);
  and _41371_ (_10145_, _10144_, _10134_);
  and _41372_ (_10146_, _10145_, _10081_);
  and _41373_ (_10148_, _10077_, word_in[28]);
  or _41374_ (_26847_[4], _10148_, _10146_);
  and _41375_ (_10149_, _10067_, word_in[5]);
  not _41376_ (_10150_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _41377_ (_10151_, _10067_, _10150_);
  nor _41378_ (_10152_, _10151_, _10149_);
  nor _41379_ (_10153_, _10152_, _10066_);
  and _41380_ (_10154_, _10066_, word_in[13]);
  or _41381_ (_10155_, _10154_, _10153_);
  and _41382_ (_10156_, _10155_, _10065_);
  and _41383_ (_10158_, _10064_, _08758_);
  or _41384_ (_10159_, _10158_, _10077_);
  or _41385_ (_10160_, _10159_, _10156_);
  or _41386_ (_10162_, _10081_, word_in[29]);
  and _41387_ (_26847_[5], _10162_, _10160_);
  or _41388_ (_10164_, _10091_, word_in[14]);
  not _41389_ (_10166_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _41390_ (_10167_, _10067_, _10166_);
  and _41391_ (_10168_, _10067_, word_in[6]);
  or _41392_ (_10170_, _10168_, _10167_);
  or _41393_ (_10171_, _10170_, _10066_);
  and _41394_ (_10173_, _10171_, _10065_);
  and _41395_ (_10174_, _10173_, _10164_);
  and _41396_ (_10175_, _10064_, _08774_);
  or _41397_ (_10176_, _10175_, _10077_);
  or _41398_ (_10177_, _10176_, _10174_);
  or _41399_ (_10178_, _10081_, word_in[30]);
  and _41400_ (_26847_[6], _10178_, _10177_);
  or _41401_ (_10180_, _10065_, _08033_);
  nor _41402_ (_10181_, _10067_, _07717_);
  and _41403_ (_10183_, _10067_, word_in[7]);
  or _41404_ (_10184_, _10183_, _10181_);
  or _41405_ (_10185_, _10184_, _10066_);
  nand _41406_ (_10187_, _10066_, _09188_);
  and _41407_ (_10189_, _10187_, _10185_);
  or _41408_ (_10190_, _10189_, _10064_);
  and _41409_ (_10191_, _10190_, _10180_);
  and _41410_ (_10193_, _10191_, _10081_);
  and _41411_ (_10195_, _10077_, word_in[31]);
  or _41412_ (_26847_[7], _10195_, _10193_);
  and _41413_ (_10198_, _02359_, _23778_);
  and _41414_ (_10199_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  or _41415_ (_27154_, _10199_, _10198_);
  and _41416_ (_10200_, _09935_, _07754_);
  and _41417_ (_10202_, _08008_, _07780_);
  not _41418_ (_10203_, _10202_);
  or _41419_ (_10204_, _10203_, _08678_);
  and _41420_ (_10205_, _08683_, _07860_);
  not _41421_ (_10207_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _41422_ (_10208_, _08688_, _08016_);
  nor _41423_ (_10209_, _10208_, _10207_);
  and _41424_ (_10210_, _10208_, _08402_);
  or _41425_ (_10211_, _10210_, _10209_);
  or _41426_ (_10213_, _10211_, _10205_);
  not _41427_ (_10214_, _10205_);
  or _41428_ (_10215_, _10214_, word_in[8]);
  and _41429_ (_10216_, _10215_, _10213_);
  or _41430_ (_10217_, _10216_, _10202_);
  and _41431_ (_10218_, _10217_, _10204_);
  or _41432_ (_10219_, _10218_, _10200_);
  not _41433_ (_10220_, _10200_);
  or _41434_ (_10222_, _10220_, word_in[24]);
  and _41435_ (_26848_[0], _10222_, _10219_);
  not _41436_ (_10223_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor _41437_ (_10224_, _10208_, _10223_);
  and _41438_ (_10226_, _10208_, _08428_);
  or _41439_ (_10228_, _10226_, _10224_);
  or _41440_ (_10229_, _10228_, _10205_);
  or _41441_ (_10230_, _10214_, word_in[9]);
  and _41442_ (_10232_, _10230_, _10229_);
  or _41443_ (_10233_, _10232_, _10202_);
  or _41444_ (_10234_, _10203_, _08422_);
  and _41445_ (_10235_, _10234_, _10233_);
  or _41446_ (_10237_, _10235_, _10200_);
  or _41447_ (_10238_, _10220_, word_in[25]);
  and _41448_ (_26848_[1], _10238_, _10237_);
  not _41449_ (_10241_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor _41450_ (_10242_, _10208_, _10241_);
  and _41451_ (_10243_, _10208_, _08591_);
  or _41452_ (_10244_, _10243_, _10242_);
  or _41453_ (_10245_, _10244_, _10205_);
  or _41454_ (_10246_, _10214_, word_in[10]);
  and _41455_ (_10247_, _10246_, _10245_);
  or _41456_ (_10248_, _10247_, _10202_);
  nor _41457_ (_10249_, _10203_, _08715_);
  nor _41458_ (_10250_, _10249_, _10200_);
  and _41459_ (_10251_, _10250_, _10248_);
  and _41460_ (_10252_, _10200_, word_in[26]);
  or _41461_ (_26848_[2], _10252_, _10251_);
  or _41462_ (_10254_, _10203_, _08728_);
  not _41463_ (_10255_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor _41464_ (_10256_, _10208_, _10255_);
  and _41465_ (_10257_, _10208_, _08604_);
  or _41466_ (_10259_, _10257_, _10256_);
  or _41467_ (_10261_, _10259_, _10205_);
  or _41468_ (_10262_, _10214_, word_in[11]);
  and _41469_ (_10263_, _10262_, _10261_);
  or _41470_ (_10264_, _10263_, _10202_);
  and _41471_ (_10265_, _10264_, _10254_);
  and _41472_ (_10266_, _10265_, _10220_);
  and _41473_ (_10267_, _10200_, word_in[27]);
  or _41474_ (_26848_[3], _10267_, _10266_);
  or _41475_ (_10268_, _10203_, _08744_);
  not _41476_ (_10269_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor _41477_ (_10270_, _10208_, _10269_);
  and _41478_ (_10271_, _10208_, _08619_);
  or _41479_ (_10272_, _10271_, _10270_);
  or _41480_ (_10273_, _10272_, _10205_);
  or _41481_ (_10274_, _10214_, word_in[12]);
  and _41482_ (_10275_, _10274_, _10273_);
  or _41483_ (_10276_, _10275_, _10202_);
  and _41484_ (_10277_, _10276_, _10268_);
  or _41485_ (_10278_, _10277_, _10200_);
  or _41486_ (_10279_, _10220_, word_in[28]);
  and _41487_ (_26848_[4], _10279_, _10278_);
  or _41488_ (_10281_, _10203_, _08758_);
  not _41489_ (_10282_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor _41490_ (_10283_, _10208_, _10282_);
  and _41491_ (_10284_, _10208_, _08501_);
  or _41492_ (_10285_, _10284_, _10283_);
  or _41493_ (_10286_, _10285_, _10205_);
  or _41494_ (_10288_, _10214_, word_in[13]);
  and _41495_ (_10290_, _10288_, _10286_);
  or _41496_ (_10292_, _10290_, _10202_);
  and _41497_ (_10294_, _10292_, _10281_);
  or _41498_ (_10295_, _10294_, _10200_);
  or _41499_ (_10296_, _10220_, word_in[29]);
  and _41500_ (_26848_[5], _10296_, _10295_);
  not _41501_ (_10298_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor _41502_ (_10299_, _10208_, _10298_);
  and _41503_ (_10300_, _10208_, _08648_);
  or _41504_ (_10302_, _10300_, _10299_);
  or _41505_ (_10303_, _10302_, _10205_);
  or _41506_ (_10305_, _10214_, word_in[14]);
  and _41507_ (_10306_, _10305_, _10303_);
  or _41508_ (_10307_, _10306_, _10202_);
  nor _41509_ (_10309_, _10203_, _08774_);
  nor _41510_ (_10311_, _10309_, _10200_);
  and _41511_ (_10312_, _10311_, _10307_);
  and _41512_ (_10313_, _10200_, word_in[30]);
  or _41513_ (_26848_[6], _10313_, _10312_);
  nor _41514_ (_10315_, _10208_, _07861_);
  and _41515_ (_10316_, _10208_, _08019_);
  or _41516_ (_10318_, _10316_, _10315_);
  or _41517_ (_10319_, _10318_, _10205_);
  nand _41518_ (_10320_, _10205_, _09188_);
  and _41519_ (_10321_, _10320_, _10319_);
  or _41520_ (_10322_, _10321_, _10202_);
  nor _41521_ (_10323_, _10203_, _08033_);
  nor _41522_ (_10324_, _10323_, _10200_);
  and _41523_ (_10325_, _10324_, _10322_);
  and _41524_ (_10326_, _10200_, word_in[31]);
  or _41525_ (_26848_[7], _10326_, _10325_);
  and _41526_ (_10327_, _05180_, _23946_);
  and _41527_ (_10328_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or _41528_ (_27132_, _10328_, _10327_);
  and _41529_ (_10331_, _06506_, _24282_);
  not _41530_ (_10332_, _10331_);
  and _41531_ (_10333_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  and _41532_ (_10334_, _10331_, _23778_);
  or _41533_ (_26981_, _10334_, _10333_);
  and _41534_ (_10335_, _05180_, _23778_);
  and _41535_ (_10337_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or _41536_ (_27130_, _10337_, _10335_);
  and _41537_ (_10339_, _08167_, _24050_);
  and _41538_ (_10340_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  or _41539_ (_27129_, _10340_, _10339_);
  and _41540_ (_10343_, _08167_, _23898_);
  and _41541_ (_10344_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  or _41542_ (_27128_, _10344_, _10343_);
  and _41543_ (_10347_, _01809_, _23986_);
  and _41544_ (_10348_, _10347_, _23946_);
  not _41545_ (_10350_, _10347_);
  and _41546_ (_10351_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  or _41547_ (_27127_, _10351_, _10348_);
  and _41548_ (_10352_, _10347_, _23747_);
  and _41549_ (_10354_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  or _41550_ (_27126_, _10354_, _10352_);
  and _41551_ (_10356_, _04797_, _24050_);
  and _41552_ (_10357_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or _41553_ (_27124_, _10357_, _10356_);
  and _41554_ (_10358_, _04797_, _23649_);
  and _41555_ (_10359_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or _41556_ (_27123_, _10359_, _10358_);
  and _41557_ (_10361_, _01810_, _24050_);
  and _41558_ (_10362_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or _41559_ (_27122_, _10362_, _10361_);
  and _41560_ (_10363_, _01810_, _23649_);
  and _41561_ (_10365_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or _41562_ (_27121_, _10365_, _10363_);
  and _41563_ (_10366_, _08954_, _08029_);
  and _41564_ (_10367_, _08017_, word_in[0]);
  not _41565_ (_10369_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor _41566_ (_10371_, _08017_, _10369_);
  nor _41567_ (_10372_, _10371_, _10367_);
  nor _41568_ (_10373_, _10372_, _08012_);
  and _41569_ (_10374_, _08012_, word_in[8]);
  or _41570_ (_10376_, _10374_, _10373_);
  and _41571_ (_10378_, _10376_, _08031_);
  and _41572_ (_10380_, _08678_, _08009_);
  or _41573_ (_10381_, _10380_, _10378_);
  and _41574_ (_10383_, _10381_, _08030_);
  or _41575_ (_26849_[0], _10383_, _10366_);
  and _41576_ (_10385_, _01810_, _23778_);
  and _41577_ (_10386_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or _41578_ (_27120_, _10386_, _10385_);
  and _41579_ (_10387_, _08017_, word_in[1]);
  not _41580_ (_10388_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor _41581_ (_10389_, _08017_, _10388_);
  nor _41582_ (_10391_, _10389_, _10387_);
  nor _41583_ (_10392_, _10391_, _08012_);
  and _41584_ (_10393_, _08012_, word_in[9]);
  or _41585_ (_10394_, _10393_, _10392_);
  and _41586_ (_10396_, _10394_, _08031_);
  and _41587_ (_10398_, _08422_, _08009_);
  or _41588_ (_10400_, _10398_, _10396_);
  and _41589_ (_10402_, _10400_, _08030_);
  and _41590_ (_10404_, _08029_, word_in[25]);
  or _41591_ (_26849_[1], _10404_, _10402_);
  and _41592_ (_10405_, _02284_, _23707_);
  and _41593_ (_10407_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or _41594_ (_27119_, _10407_, _10405_);
  and _41595_ (_10408_, _08017_, word_in[2]);
  not _41596_ (_10410_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _41597_ (_10411_, _08017_, _10410_);
  nor _41598_ (_10412_, _10411_, _10408_);
  nor _41599_ (_10414_, _10412_, _08012_);
  and _41600_ (_10415_, _08012_, word_in[10]);
  or _41601_ (_10417_, _10415_, _10414_);
  and _41602_ (_10418_, _10417_, _08031_);
  and _41603_ (_10419_, _08715_, _08009_);
  or _41604_ (_10420_, _10419_, _10418_);
  and _41605_ (_10421_, _10420_, _08030_);
  and _41606_ (_10422_, _08993_, _08029_);
  or _41607_ (_26849_[2], _10422_, _10421_);
  and _41608_ (_10423_, _02284_, _23946_);
  and _41609_ (_10424_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  or _41610_ (_27118_, _10424_, _10423_);
  and _41611_ (_10425_, _08017_, word_in[3]);
  not _41612_ (_10426_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor _41613_ (_10427_, _08017_, _10426_);
  nor _41614_ (_10428_, _10427_, _10425_);
  nor _41615_ (_10429_, _10428_, _08012_);
  and _41616_ (_10430_, _08012_, word_in[11]);
  or _41617_ (_10432_, _10430_, _10429_);
  and _41618_ (_10433_, _10432_, _08031_);
  and _41619_ (_10434_, _08728_, _08009_);
  or _41620_ (_10435_, _10434_, _10433_);
  and _41621_ (_10437_, _10435_, _08030_);
  and _41622_ (_10438_, _08029_, word_in[27]);
  or _41623_ (_26849_[3], _10438_, _10437_);
  and _41624_ (_10439_, _08481_, _08029_);
  and _41625_ (_10440_, _08017_, word_in[4]);
  not _41626_ (_10441_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor _41627_ (_10442_, _08017_, _10441_);
  nor _41628_ (_10443_, _10442_, _10440_);
  nor _41629_ (_10444_, _10443_, _08012_);
  and _41630_ (_10445_, _08012_, word_in[12]);
  or _41631_ (_10446_, _10445_, _10444_);
  and _41632_ (_10447_, _10446_, _08031_);
  and _41633_ (_10448_, _08744_, _08009_);
  or _41634_ (_10449_, _10448_, _10447_);
  and _41635_ (_10450_, _10449_, _08030_);
  or _41636_ (_26849_[4], _10450_, _10439_);
  and _41637_ (_10451_, _08017_, word_in[5]);
  not _41638_ (_10453_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor _41639_ (_10455_, _08017_, _10453_);
  nor _41640_ (_10456_, _10455_, _10451_);
  nor _41641_ (_10457_, _10456_, _08012_);
  and _41642_ (_10458_, _08012_, word_in[13]);
  or _41643_ (_10459_, _10458_, _10457_);
  and _41644_ (_10460_, _10459_, _08031_);
  and _41645_ (_10461_, _08758_, _08009_);
  or _41646_ (_10462_, _10461_, _10460_);
  and _41647_ (_10463_, _10462_, _08030_);
  and _41648_ (_10464_, _08029_, word_in[29]);
  or _41649_ (_26849_[5], _10464_, _10463_);
  and _41650_ (_10465_, _08510_, _08029_);
  and _41651_ (_10466_, _08017_, word_in[6]);
  not _41652_ (_10467_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor _41653_ (_10468_, _08017_, _10467_);
  nor _41654_ (_10469_, _10468_, _10466_);
  nor _41655_ (_10470_, _10469_, _08012_);
  and _41656_ (_10472_, _08012_, word_in[14]);
  or _41657_ (_10473_, _10472_, _10470_);
  and _41658_ (_10474_, _10473_, _08031_);
  and _41659_ (_10475_, _08774_, _08009_);
  or _41660_ (_10476_, _10475_, _10474_);
  and _41661_ (_10477_, _10476_, _08030_);
  or _41662_ (_26849_[6], _10477_, _10465_);
  and _41663_ (_10478_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and _41664_ (_10479_, _08351_, _23946_);
  or _41665_ (_02826_, _10479_, _10478_);
  and _41666_ (_10480_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  and _41667_ (_10481_, _08375_, _23946_);
  or _41668_ (_02844_, _10481_, _10480_);
  and _41669_ (_10482_, _02302_, _23649_);
  and _41670_ (_10483_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or _41671_ (_02874_, _10483_, _10482_);
  and _41672_ (_10484_, _02302_, _23778_);
  and _41673_ (_10485_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or _41674_ (_02876_, _10485_, _10484_);
  and _41675_ (_10486_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  and _41676_ (_10487_, _08375_, _24050_);
  or _41677_ (_02880_, _10487_, _10486_);
  and _41678_ (_10488_, _02374_, _23946_);
  and _41679_ (_10489_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or _41680_ (_02882_, _10489_, _10488_);
  and _41681_ (_10490_, _03339_, _23747_);
  and _41682_ (_10491_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or _41683_ (_27113_, _10491_, _10490_);
  and _41684_ (_10492_, _03339_, _23898_);
  and _41685_ (_10493_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or _41686_ (_27111_, _10493_, _10492_);
  and _41687_ (_10494_, _24766_, _24282_);
  not _41688_ (_10495_, _10494_);
  and _41689_ (_10496_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and _41690_ (_10497_, _10494_, _23778_);
  or _41691_ (_02893_, _10497_, _10496_);
  and _41692_ (_10498_, _04917_, _23649_);
  and _41693_ (_10499_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or _41694_ (_27109_, _10499_, _10498_);
  and _41695_ (_10501_, _04917_, _23824_);
  and _41696_ (_10502_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or _41697_ (_02906_, _10502_, _10501_);
  and _41698_ (_10503_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  and _41699_ (_10504_, _10494_, _23898_);
  or _41700_ (_02908_, _10504_, _10503_);
  and _41701_ (_10505_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  and _41702_ (_10506_, _10494_, _23747_);
  or _41703_ (_02911_, _10506_, _10505_);
  and _41704_ (_10507_, _07471_, _24050_);
  and _41705_ (_10508_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  or _41706_ (_02923_, _10508_, _10507_);
  and _41707_ (_10509_, _07673_, word_in[0]);
  nand _41708_ (_10510_, _07570_, _08556_);
  or _41709_ (_10512_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _41710_ (_10513_, _10512_, _10510_);
  and _41711_ (_10514_, _10513_, _07624_);
  or _41712_ (_10515_, _10514_, _07577_);
  nand _41713_ (_10517_, _07570_, _09080_);
  or _41714_ (_10518_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _41715_ (_10519_, _10518_, _10517_);
  and _41716_ (_10520_, _10519_, _07591_);
  nand _41717_ (_10521_, _07570_, _09333_);
  or _41718_ (_10522_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _41719_ (_10523_, _10522_, _10521_);
  and _41720_ (_10524_, _10523_, _07608_);
  nand _41721_ (_10525_, _07570_, _08809_);
  or _41722_ (_10526_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _41723_ (_10527_, _10526_, _10525_);
  and _41724_ (_10528_, _10527_, _07597_);
  or _41725_ (_10529_, _10528_, _10524_);
  or _41726_ (_10530_, _10529_, _10520_);
  or _41727_ (_10531_, _10530_, _10515_);
  nand _41728_ (_10532_, _07570_, _09570_);
  or _41729_ (_10533_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _41730_ (_10534_, _10533_, _10532_);
  and _41731_ (_10535_, _10534_, _07624_);
  or _41732_ (_10536_, _10535_, _07648_);
  nand _41733_ (_10537_, _07570_, _10069_);
  or _41734_ (_10538_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _41735_ (_10539_, _10538_, _10537_);
  and _41736_ (_10541_, _10539_, _07591_);
  nand _41737_ (_10542_, _07570_, _10369_);
  or _41738_ (_10543_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _41739_ (_10544_, _10543_, _10542_);
  and _41740_ (_10545_, _10544_, _07608_);
  nand _41741_ (_10546_, _07570_, _09802_);
  or _41742_ (_10547_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _41743_ (_10548_, _10547_, _10546_);
  and _41744_ (_10549_, _10548_, _07597_);
  or _41745_ (_10551_, _10549_, _10545_);
  or _41746_ (_10552_, _10551_, _10541_);
  or _41747_ (_10553_, _10552_, _10536_);
  and _41748_ (_10554_, _10553_, _10531_);
  and _41749_ (_10555_, _10554_, _07672_);
  or _41750_ (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _10555_, _10509_);
  and _41751_ (_10556_, _07673_, word_in[1]);
  nand _41752_ (_10557_, _07570_, _08575_);
  or _41753_ (_10558_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _41754_ (_10560_, _10558_, _10557_);
  and _41755_ (_10561_, _10560_, _07624_);
  or _41756_ (_10562_, _10561_, _07577_);
  nand _41757_ (_10563_, _07570_, _09098_);
  or _41758_ (_10564_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _41759_ (_10565_, _10564_, _10563_);
  and _41760_ (_10566_, _10565_, _07591_);
  nand _41761_ (_10567_, _07570_, _09352_);
  or _41762_ (_10568_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _41763_ (_10570_, _10568_, _10567_);
  and _41764_ (_10571_, _10570_, _07608_);
  nand _41765_ (_10572_, _07570_, _08830_);
  or _41766_ (_10573_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _41767_ (_10575_, _10573_, _10572_);
  and _41768_ (_10576_, _10575_, _07597_);
  or _41769_ (_10577_, _10576_, _10571_);
  or _41770_ (_10578_, _10577_, _10566_);
  or _41771_ (_10579_, _10578_, _10562_);
  nand _41772_ (_10580_, _07570_, _09586_);
  or _41773_ (_10581_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _41774_ (_10582_, _10581_, _10580_);
  and _41775_ (_10583_, _10582_, _07624_);
  or _41776_ (_10584_, _10583_, _07648_);
  nand _41777_ (_10585_, _07570_, _10084_);
  or _41778_ (_10586_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _41779_ (_10587_, _10586_, _10585_);
  and _41780_ (_10588_, _10587_, _07591_);
  nand _41781_ (_10589_, _07570_, _10388_);
  or _41782_ (_10590_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _41783_ (_10591_, _10590_, _10589_);
  and _41784_ (_10592_, _10591_, _07608_);
  nand _41785_ (_10593_, _07570_, _09819_);
  or _41786_ (_10594_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _41787_ (_10595_, _10594_, _10593_);
  and _41788_ (_10596_, _10595_, _07597_);
  or _41789_ (_10597_, _10596_, _10592_);
  or _41790_ (_10598_, _10597_, _10588_);
  or _41791_ (_10600_, _10598_, _10584_);
  and _41792_ (_10601_, _10600_, _10579_);
  and _41793_ (_10602_, _10601_, _07672_);
  or _41794_ (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _10602_, _10556_);
  and _41795_ (_10603_, _07673_, word_in[2]);
  nand _41796_ (_10605_, _07570_, _08844_);
  or _41797_ (_10607_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _41798_ (_10608_, _10607_, _10605_);
  and _41799_ (_10609_, _10608_, _07597_);
  or _41800_ (_10610_, _10609_, _07577_);
  nand _41801_ (_10611_, _07570_, _09113_);
  or _41802_ (_10612_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _41803_ (_10613_, _10612_, _10611_);
  and _41804_ (_10614_, _10613_, _07591_);
  nand _41805_ (_10615_, _07570_, _09371_);
  or _41806_ (_10616_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _41807_ (_10617_, _10616_, _10615_);
  and _41808_ (_10618_, _10617_, _07608_);
  nand _41809_ (_10619_, _07570_, _08589_);
  or _41810_ (_10620_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _41811_ (_10621_, _10620_, _10619_);
  and _41812_ (_10622_, _10621_, _07624_);
  or _41813_ (_10624_, _10622_, _10618_);
  or _41814_ (_10626_, _10624_, _10614_);
  or _41815_ (_10627_, _10626_, _10610_);
  nand _41816_ (_10629_, _07570_, _09834_);
  or _41817_ (_10630_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _41818_ (_10631_, _10630_, _10629_);
  and _41819_ (_10632_, _10631_, _07597_);
  or _41820_ (_10633_, _10632_, _07648_);
  nand _41821_ (_10634_, _07570_, _10410_);
  or _41822_ (_10635_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _41823_ (_10636_, _10635_, _10634_);
  and _41824_ (_10637_, _10636_, _07608_);
  nand _41825_ (_10638_, _07570_, _10102_);
  or _41826_ (_10639_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _41827_ (_10640_, _10639_, _10638_);
  and _41828_ (_10642_, _10640_, _07591_);
  or _41829_ (_10643_, _10642_, _10637_);
  nand _41830_ (_10644_, _07570_, _09598_);
  or _41831_ (_10645_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _41832_ (_10647_, _10645_, _10644_);
  and _41833_ (_10648_, _10647_, _07624_);
  or _41834_ (_10649_, _10648_, _10643_);
  or _41835_ (_10651_, _10649_, _10633_);
  and _41836_ (_10653_, _10651_, _10627_);
  and _41837_ (_10654_, _10653_, _07672_);
  or _41838_ (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _10654_, _10603_);
  and _41839_ (_10655_, _07673_, word_in[3]);
  nand _41840_ (_10656_, _07570_, _08857_);
  or _41841_ (_10658_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _41842_ (_10659_, _10658_, _10656_);
  and _41843_ (_10661_, _10659_, _07597_);
  or _41844_ (_10662_, _10661_, _07577_);
  nand _41845_ (_10663_, _07570_, _09128_);
  or _41846_ (_10664_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _41847_ (_10665_, _10664_, _10663_);
  and _41848_ (_10666_, _10665_, _07591_);
  nand _41849_ (_10667_, _07570_, _09389_);
  or _41850_ (_10668_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _41851_ (_10669_, _10668_, _10667_);
  and _41852_ (_10670_, _10669_, _07608_);
  nand _41853_ (_10671_, _07570_, _08602_);
  or _41854_ (_10672_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _41855_ (_10673_, _10672_, _10671_);
  and _41856_ (_10674_, _10673_, _07624_);
  or _41857_ (_10675_, _10674_, _10670_);
  or _41858_ (_10676_, _10675_, _10666_);
  or _41859_ (_10678_, _10676_, _10662_);
  nand _41860_ (_10680_, _07570_, _09849_);
  or _41861_ (_10681_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _41862_ (_10682_, _10681_, _10680_);
  and _41863_ (_10683_, _10682_, _07597_);
  or _41864_ (_10684_, _10683_, _07648_);
  nand _41865_ (_10685_, _07570_, _10426_);
  or _41866_ (_10686_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _41867_ (_10687_, _10686_, _10685_);
  and _41868_ (_10688_, _10687_, _07608_);
  nand _41869_ (_10689_, _07570_, _10118_);
  or _41870_ (_10690_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and _41871_ (_10691_, _10690_, _10689_);
  and _41872_ (_10692_, _10691_, _07591_);
  or _41873_ (_10693_, _10692_, _10688_);
  nand _41874_ (_10694_, _07570_, _09613_);
  or _41875_ (_10695_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and _41876_ (_10696_, _10695_, _10694_);
  and _41877_ (_10697_, _10696_, _07624_);
  or _41878_ (_10698_, _10697_, _10693_);
  or _41879_ (_10699_, _10698_, _10684_);
  and _41880_ (_10700_, _10699_, _10678_);
  and _41881_ (_10702_, _10700_, _07672_);
  or _41882_ (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _10702_, _10655_);
  and _41883_ (_10703_, _07673_, word_in[4]);
  nand _41884_ (_10704_, _07570_, _08617_);
  or _41885_ (_10705_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _41886_ (_10707_, _10705_, _10704_);
  and _41887_ (_10708_, _10707_, _07624_);
  or _41888_ (_10709_, _10708_, _07577_);
  nand _41889_ (_10711_, _07570_, _09141_);
  or _41890_ (_10712_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _41891_ (_10713_, _10712_, _10711_);
  and _41892_ (_10714_, _10713_, _07591_);
  nand _41893_ (_10715_, _07570_, _09402_);
  or _41894_ (_10716_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _41895_ (_10717_, _10716_, _10715_);
  and _41896_ (_10719_, _10717_, _07608_);
  nand _41897_ (_10720_, _07570_, _08870_);
  or _41898_ (_10721_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _41899_ (_10722_, _10721_, _10720_);
  and _41900_ (_10723_, _10722_, _07597_);
  or _41901_ (_10724_, _10723_, _10719_);
  or _41902_ (_10725_, _10724_, _10714_);
  or _41903_ (_10726_, _10725_, _10709_);
  nand _41904_ (_10727_, _07570_, _09627_);
  or _41905_ (_10728_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and _41906_ (_10729_, _10728_, _10727_);
  and _41907_ (_10730_, _10729_, _07624_);
  or _41908_ (_10732_, _10730_, _07648_);
  nand _41909_ (_10733_, _07570_, _10135_);
  or _41910_ (_10734_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and _41911_ (_10736_, _10734_, _10733_);
  and _41912_ (_10738_, _10736_, _07591_);
  nand _41913_ (_10739_, _07570_, _10441_);
  or _41914_ (_10740_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _41915_ (_10741_, _10740_, _10739_);
  and _41916_ (_10743_, _10741_, _07608_);
  nand _41917_ (_10744_, _07570_, _09863_);
  or _41918_ (_10746_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _41919_ (_10747_, _10746_, _10744_);
  and _41920_ (_10749_, _10747_, _07597_);
  or _41921_ (_10751_, _10749_, _10743_);
  or _41922_ (_10752_, _10751_, _10738_);
  or _41923_ (_10753_, _10752_, _10732_);
  and _41924_ (_10754_, _10753_, _10726_);
  and _41925_ (_10756_, _10754_, _07672_);
  or _41926_ (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _10756_, _10703_);
  and _41927_ (_10758_, _07673_, word_in[5]);
  nand _41928_ (_10759_, _07570_, _08630_);
  or _41929_ (_10760_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _41930_ (_10761_, _10760_, _10759_);
  and _41931_ (_10762_, _10761_, _07624_);
  or _41932_ (_10763_, _10762_, _07577_);
  nand _41933_ (_10764_, _07570_, _09153_);
  or _41934_ (_10765_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _41935_ (_10766_, _10765_, _10764_);
  and _41936_ (_10767_, _10766_, _07591_);
  nand _41937_ (_10768_, _07570_, _09415_);
  or _41938_ (_10769_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _41939_ (_10771_, _10769_, _10768_);
  and _41940_ (_10772_, _10771_, _07608_);
  nand _41941_ (_10773_, _07570_, _08883_);
  or _41942_ (_10774_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _41943_ (_10776_, _10774_, _10773_);
  and _41944_ (_10777_, _10776_, _07597_);
  or _41945_ (_10778_, _10777_, _10772_);
  or _41946_ (_10781_, _10778_, _10767_);
  or _41947_ (_10782_, _10781_, _10763_);
  nand _41948_ (_10783_, _07570_, _09641_);
  or _41949_ (_10785_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _41950_ (_10786_, _10785_, _10783_);
  and _41951_ (_10787_, _10786_, _07624_);
  or _41952_ (_10789_, _10787_, _07648_);
  nand _41953_ (_10790_, _07570_, _10150_);
  or _41954_ (_10792_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _41955_ (_10793_, _10792_, _10790_);
  and _41956_ (_10794_, _10793_, _07591_);
  nand _41957_ (_10795_, _07570_, _10453_);
  or _41958_ (_10796_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _41959_ (_10798_, _10796_, _10795_);
  and _41960_ (_10800_, _10798_, _07608_);
  nand _41961_ (_10801_, _07570_, _09875_);
  or _41962_ (_10802_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _41963_ (_10803_, _10802_, _10801_);
  and _41964_ (_10804_, _10803_, _07597_);
  or _41965_ (_10805_, _10804_, _10800_);
  or _41966_ (_10807_, _10805_, _10794_);
  or _41967_ (_10808_, _10807_, _10789_);
  and _41968_ (_10809_, _10808_, _10782_);
  and _41969_ (_10811_, _10809_, _07672_);
  or _41970_ (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _10811_, _10758_);
  and _41971_ (_10812_, _07673_, word_in[6]);
  nand _41972_ (_10814_, _07570_, _08898_);
  or _41973_ (_10815_, _07570_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _41974_ (_10816_, _10815_, _10814_);
  and _41975_ (_10817_, _10816_, _07597_);
  or _41976_ (_10818_, _10817_, _07577_);
  nand _41977_ (_10819_, _07570_, _09166_);
  or _41978_ (_10820_, _07570_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _41979_ (_10821_, _10820_, _10819_);
  and _41980_ (_10822_, _10821_, _07591_);
  nand _41981_ (_10823_, _07570_, _09428_);
  or _41982_ (_10824_, _07570_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _41983_ (_10825_, _10824_, _10823_);
  and _41984_ (_10827_, _10825_, _07608_);
  nand _41985_ (_10828_, _07570_, _08646_);
  or _41986_ (_10831_, _07570_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _41987_ (_10833_, _10831_, _10828_);
  and _41988_ (_10835_, _10833_, _07624_);
  or _41989_ (_10836_, _10835_, _10827_);
  or _41990_ (_10837_, _10836_, _10822_);
  or _41991_ (_10839_, _10837_, _10818_);
  nand _41992_ (_10840_, _07570_, _09888_);
  or _41993_ (_10841_, _07570_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _41994_ (_10842_, _10841_, _10840_);
  and _41995_ (_10843_, _10842_, _07597_);
  or _41996_ (_10845_, _10843_, _07648_);
  nand _41997_ (_10846_, _07570_, _10467_);
  or _41998_ (_10847_, _07570_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _41999_ (_10848_, _10847_, _10846_);
  and _42000_ (_10849_, _10848_, _07608_);
  nand _42001_ (_10850_, _07570_, _10166_);
  or _42002_ (_10851_, _07570_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _42003_ (_10852_, _10851_, _10850_);
  and _42004_ (_10853_, _10852_, _07591_);
  or _42005_ (_10854_, _10853_, _10849_);
  nand _42006_ (_10857_, _07570_, _09654_);
  or _42007_ (_10858_, _07570_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _42008_ (_10859_, _10858_, _10857_);
  and _42009_ (_10860_, _10859_, _07624_);
  or _42010_ (_10861_, _10860_, _10854_);
  or _42011_ (_10862_, _10861_, _10845_);
  and _42012_ (_10863_, _10862_, _10839_);
  and _42013_ (_10865_, _10863_, _07672_);
  or _42014_ (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _10865_, _10812_);
  and _42015_ (_10866_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  and _42016_ (_10867_, _10494_, _23649_);
  or _42017_ (_27024_, _10867_, _10866_);
  and _42018_ (_10868_, _07810_, word_in[8]);
  nand _42019_ (_10869_, _07570_, _08686_);
  or _42020_ (_10870_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _42021_ (_10871_, _10870_, _10869_);
  and _42022_ (_10872_, _10871_, _07812_);
  nand _42023_ (_10874_, _07570_, _08393_);
  or _42024_ (_10875_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _42025_ (_10877_, _10875_, _10874_);
  and _42026_ (_10878_, _10877_, _07811_);
  or _42027_ (_10879_, _10878_, _10872_);
  and _42028_ (_10881_, _10879_, _07766_);
  nand _42029_ (_10882_, _07570_, _09686_);
  or _42030_ (_10883_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _42031_ (_10884_, _10883_, _10882_);
  and _42032_ (_10885_, _10884_, _07812_);
  nand _42033_ (_10887_, _07570_, _09453_);
  or _42034_ (_10889_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _42035_ (_10890_, _10889_, _10887_);
  and _42036_ (_10893_, _10890_, _07811_);
  or _42037_ (_10894_, _10893_, _10885_);
  and _42038_ (_10896_, _10894_, _07770_);
  nand _42039_ (_10898_, _07570_, _09200_);
  or _42040_ (_10899_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _42041_ (_10900_, _10899_, _10898_);
  and _42042_ (_10901_, _10900_, _07812_);
  nand _42043_ (_10903_, _07570_, _08938_);
  or _42044_ (_10904_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _42045_ (_10905_, _10904_, _10903_);
  and _42046_ (_10906_, _10905_, _07811_);
  or _42047_ (_10907_, _10906_, _10901_);
  and _42048_ (_10908_, _10907_, _07845_);
  nand _42049_ (_10909_, _07570_, _10207_);
  or _42050_ (_10910_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _42051_ (_10911_, _10910_, _10909_);
  and _42052_ (_10912_, _10911_, _07812_);
  nand _42053_ (_10913_, _07570_, _09946_);
  or _42054_ (_10914_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _42055_ (_10916_, _10914_, _10913_);
  and _42056_ (_10917_, _10916_, _07811_);
  or _42057_ (_10918_, _10917_, _10912_);
  and _42058_ (_10919_, _10918_, _07860_);
  or _42059_ (_10921_, _10919_, _10908_);
  or _42060_ (_10922_, _10921_, _10896_);
  nor _42061_ (_10923_, _10922_, _10881_);
  nor _42062_ (_10924_, _10923_, _07810_);
  or _42063_ (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _10924_, _10868_);
  and _42064_ (_10925_, _07810_, word_in[9]);
  nand _42065_ (_10926_, _07570_, _08702_);
  or _42066_ (_10927_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _42067_ (_10929_, _10927_, _10926_);
  and _42068_ (_10931_, _10929_, _07812_);
  nand _42069_ (_10932_, _07570_, _08425_);
  or _42070_ (_10933_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _42071_ (_10934_, _10933_, _10932_);
  and _42072_ (_10935_, _10934_, _07811_);
  or _42073_ (_10936_, _10935_, _10931_);
  and _42074_ (_10937_, _10936_, _07766_);
  nand _42075_ (_10939_, _07570_, _09703_);
  or _42076_ (_10941_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _42077_ (_10942_, _10941_, _10939_);
  and _42078_ (_10943_, _10942_, _07812_);
  nand _42079_ (_10944_, _07570_, _09474_);
  or _42080_ (_10946_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _42081_ (_10948_, _10946_, _10944_);
  and _42082_ (_10949_, _10948_, _07811_);
  or _42083_ (_10950_, _10949_, _10943_);
  and _42084_ (_10951_, _10950_, _07770_);
  nand _42085_ (_10953_, _07570_, _09222_);
  or _42086_ (_10954_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _42087_ (_10956_, _10954_, _10953_);
  and _42088_ (_10957_, _10956_, _07812_);
  nand _42089_ (_10959_, _07570_, _08957_);
  or _42090_ (_10961_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and _42091_ (_10962_, _10961_, _10959_);
  and _42092_ (_10963_, _10962_, _07811_);
  or _42093_ (_10964_, _10963_, _10957_);
  and _42094_ (_10965_, _10964_, _07845_);
  nand _42095_ (_10967_, _07570_, _10223_);
  or _42096_ (_10969_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _42097_ (_10970_, _10969_, _10967_);
  and _42098_ (_10971_, _10970_, _07812_);
  nand _42099_ (_10972_, _07570_, _09963_);
  or _42100_ (_10974_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _42101_ (_10976_, _10974_, _10972_);
  and _42102_ (_10977_, _10976_, _07811_);
  or _42103_ (_10978_, _10977_, _10971_);
  and _42104_ (_10979_, _10978_, _07860_);
  or _42105_ (_10981_, _10979_, _10965_);
  or _42106_ (_10983_, _10981_, _10951_);
  nor _42107_ (_10984_, _10983_, _10937_);
  nor _42108_ (_10985_, _10984_, _07810_);
  or _42109_ (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _10985_, _10925_);
  and _42110_ (_10986_, _07810_, word_in[10]);
  nand _42111_ (_10987_, _07570_, _08717_);
  or _42112_ (_10988_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _42113_ (_10989_, _10988_, _10987_);
  and _42114_ (_10990_, _10989_, _07812_);
  nand _42115_ (_10991_, _07570_, _08450_);
  or _42116_ (_10992_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _42117_ (_10993_, _10992_, _10991_);
  and _42118_ (_10994_, _10993_, _07811_);
  or _42119_ (_10995_, _10994_, _10990_);
  and _42120_ (_10996_, _10995_, _07766_);
  nand _42121_ (_10997_, _07570_, _09716_);
  or _42122_ (_10998_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _42123_ (_10999_, _10998_, _10997_);
  and _42124_ (_11000_, _10999_, _07812_);
  nand _42125_ (_11001_, _07570_, _09486_);
  or _42126_ (_11002_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _42127_ (_11003_, _11002_, _11001_);
  and _42128_ (_11004_, _11003_, _07811_);
  or _42129_ (_11005_, _11004_, _11000_);
  and _42130_ (_11006_, _11005_, _07770_);
  nand _42131_ (_11007_, _07570_, _09236_);
  or _42132_ (_11008_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _42133_ (_11009_, _11008_, _11007_);
  and _42134_ (_11010_, _11009_, _07812_);
  nand _42135_ (_11011_, _07570_, _08979_);
  or _42136_ (_11012_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and _42137_ (_11013_, _11012_, _11011_);
  and _42138_ (_11014_, _11013_, _07811_);
  or _42139_ (_11015_, _11014_, _11010_);
  and _42140_ (_11016_, _11015_, _07845_);
  nand _42141_ (_11017_, _07570_, _10241_);
  or _42142_ (_11018_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _42143_ (_11019_, _11018_, _11017_);
  and _42144_ (_11020_, _11019_, _07812_);
  nand _42145_ (_11021_, _07570_, _09979_);
  or _42146_ (_11022_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and _42147_ (_11023_, _11022_, _11021_);
  and _42148_ (_11024_, _11023_, _07811_);
  or _42149_ (_11025_, _11024_, _11020_);
  and _42150_ (_11026_, _11025_, _07860_);
  or _42151_ (_11027_, _11026_, _11016_);
  or _42152_ (_11028_, _11027_, _11006_);
  nor _42153_ (_11029_, _11028_, _10996_);
  nor _42154_ (_11030_, _11029_, _07810_);
  or _42155_ (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _11030_, _10986_);
  and _42156_ (_11031_, _07810_, word_in[11]);
  nand _42157_ (_11032_, _07570_, _08730_);
  or _42158_ (_11033_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _42159_ (_11034_, _11033_, _11032_);
  and _42160_ (_11035_, _11034_, _07812_);
  nand _42161_ (_11036_, _07570_, _08467_);
  or _42162_ (_11037_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and _42163_ (_11038_, _11037_, _11036_);
  and _42164_ (_11039_, _11038_, _07811_);
  or _42165_ (_11040_, _11039_, _11035_);
  and _42166_ (_11041_, _11040_, _07766_);
  nand _42167_ (_11042_, _07570_, _09732_);
  or _42168_ (_11043_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _42169_ (_11044_, _11043_, _11042_);
  and _42170_ (_11045_, _11044_, _07812_);
  nand _42171_ (_11046_, _07570_, _09499_);
  or _42172_ (_11047_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _42173_ (_11048_, _11047_, _11046_);
  and _42174_ (_11049_, _11048_, _07811_);
  or _42175_ (_11050_, _11049_, _11045_);
  and _42176_ (_11052_, _11050_, _07770_);
  nand _42177_ (_11054_, _07570_, _09248_);
  or _42178_ (_11055_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _42179_ (_11056_, _11055_, _11054_);
  and _42180_ (_11058_, _11056_, _07812_);
  nand _42181_ (_11059_, _07570_, _08996_);
  or _42182_ (_11060_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and _42183_ (_11061_, _11060_, _11059_);
  and _42184_ (_11063_, _11061_, _07811_);
  or _42185_ (_11064_, _11063_, _11058_);
  and _42186_ (_11065_, _11064_, _07845_);
  nand _42187_ (_11066_, _07570_, _10255_);
  or _42188_ (_11067_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _42189_ (_11068_, _11067_, _11066_);
  and _42190_ (_11069_, _11068_, _07812_);
  nand _42191_ (_11070_, _07570_, _09994_);
  or _42192_ (_11072_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _42193_ (_11073_, _11072_, _11070_);
  and _42194_ (_11075_, _11073_, _07811_);
  or _42195_ (_11076_, _11075_, _11069_);
  and _42196_ (_11078_, _11076_, _07860_);
  or _42197_ (_11079_, _11078_, _11065_);
  or _42198_ (_11081_, _11079_, _11052_);
  nor _42199_ (_11082_, _11081_, _11041_);
  nor _42200_ (_11084_, _11082_, _07810_);
  or _42201_ (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _11084_, _11031_);
  and _42202_ (_11087_, _07810_, word_in[12]);
  nand _42203_ (_11088_, _07570_, _08746_);
  or _42204_ (_11089_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _42205_ (_11090_, _11089_, _11088_);
  and _42206_ (_11093_, _11090_, _07812_);
  nand _42207_ (_11095_, _07570_, _08485_);
  or _42208_ (_11096_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _42209_ (_11097_, _11096_, _11095_);
  and _42210_ (_11098_, _11097_, _07811_);
  or _42211_ (_11099_, _11098_, _11093_);
  and _42212_ (_11101_, _11099_, _07766_);
  nand _42213_ (_11103_, _07570_, _09746_);
  or _42214_ (_11105_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _42215_ (_11107_, _11105_, _11103_);
  and _42216_ (_11108_, _11107_, _07812_);
  nand _42217_ (_11110_, _07570_, _09512_);
  or _42218_ (_11112_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _42219_ (_11113_, _11112_, _11110_);
  and _42220_ (_11114_, _11113_, _07811_);
  or _42221_ (_11115_, _11114_, _11108_);
  and _42222_ (_11116_, _11115_, _07770_);
  nand _42223_ (_11118_, _07570_, _09262_);
  or _42224_ (_11120_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _42225_ (_11121_, _11120_, _11118_);
  and _42226_ (_11122_, _11121_, _07812_);
  nand _42227_ (_11123_, _07570_, _09013_);
  or _42228_ (_11125_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _42229_ (_11126_, _11125_, _11123_);
  and _42230_ (_11128_, _11126_, _07811_);
  or _42231_ (_11129_, _11128_, _11122_);
  and _42232_ (_11130_, _11129_, _07845_);
  nand _42233_ (_11131_, _07570_, _10269_);
  or _42234_ (_11133_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _42235_ (_11135_, _11133_, _11131_);
  and _42236_ (_11137_, _11135_, _07812_);
  nand _42237_ (_11138_, _07570_, _10008_);
  or _42238_ (_11140_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and _42239_ (_11142_, _11140_, _11138_);
  and _42240_ (_11143_, _11142_, _07811_);
  or _42241_ (_11144_, _11143_, _11137_);
  and _42242_ (_11145_, _11144_, _07860_);
  or _42243_ (_11146_, _11145_, _11130_);
  or _42244_ (_11148_, _11146_, _11116_);
  nor _42245_ (_11150_, _11148_, _11101_);
  nor _42246_ (_11151_, _11150_, _07810_);
  or _42247_ (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _11151_, _11087_);
  and _42248_ (_11152_, _07810_, word_in[13]);
  nand _42249_ (_11154_, _07570_, _08760_);
  or _42250_ (_11155_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _42251_ (_11157_, _11155_, _11154_);
  and _42252_ (_11158_, _11157_, _07812_);
  nand _42253_ (_11160_, _07570_, _08499_);
  or _42254_ (_11162_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _42255_ (_11163_, _11162_, _11160_);
  and _42256_ (_11165_, _11163_, _07811_);
  or _42257_ (_11166_, _11165_, _11158_);
  and _42258_ (_11167_, _11166_, _07766_);
  nand _42259_ (_11168_, _07570_, _09760_);
  or _42260_ (_11169_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _42261_ (_11170_, _11169_, _11168_);
  and _42262_ (_11171_, _11170_, _07812_);
  nand _42263_ (_11172_, _07570_, _09525_);
  or _42264_ (_11173_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _42265_ (_11174_, _11173_, _11172_);
  and _42266_ (_11176_, _11174_, _07811_);
  or _42267_ (_11177_, _11176_, _11171_);
  and _42268_ (_11178_, _11177_, _07770_);
  nand _42269_ (_11179_, _07570_, _09279_);
  or _42270_ (_11180_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _42271_ (_11181_, _11180_, _11179_);
  and _42272_ (_11182_, _11181_, _07812_);
  nand _42273_ (_11184_, _07570_, _09029_);
  or _42274_ (_11185_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and _42275_ (_11186_, _11185_, _11184_);
  and _42276_ (_11187_, _11186_, _07811_);
  or _42277_ (_11188_, _11187_, _11182_);
  and _42278_ (_11190_, _11188_, _07845_);
  nand _42279_ (_11191_, _07570_, _10282_);
  or _42280_ (_11192_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _42281_ (_11194_, _11192_, _11191_);
  and _42282_ (_11196_, _11194_, _07812_);
  nand _42283_ (_11197_, _07570_, _10023_);
  or _42284_ (_11198_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _42285_ (_11199_, _11198_, _11197_);
  and _42286_ (_11201_, _11199_, _07811_);
  or _42287_ (_11202_, _11201_, _11196_);
  and _42288_ (_11204_, _11202_, _07860_);
  or _42289_ (_11205_, _11204_, _11190_);
  or _42290_ (_11206_, _11205_, _11178_);
  nor _42291_ (_11208_, _11206_, _11167_);
  nor _42292_ (_11209_, _11208_, _07810_);
  or _42293_ (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _11209_, _11152_);
  and _42294_ (_11210_, _07810_, word_in[14]);
  nand _42295_ (_11211_, _07570_, _08776_);
  or _42296_ (_11212_, _07570_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _42297_ (_11213_, _11212_, _11211_);
  and _42298_ (_11214_, _11213_, _07812_);
  nand _42299_ (_11215_, _07570_, _08515_);
  or _42300_ (_11217_, _07570_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _42301_ (_11218_, _11217_, _11215_);
  and _42302_ (_11219_, _11218_, _07811_);
  or _42303_ (_11220_, _11219_, _11214_);
  and _42304_ (_11221_, _11220_, _07766_);
  nand _42305_ (_11223_, _07570_, _09774_);
  or _42306_ (_11224_, _07570_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _42307_ (_11225_, _11224_, _11223_);
  and _42308_ (_11226_, _11225_, _07812_);
  nand _42309_ (_11227_, _07570_, _09537_);
  or _42310_ (_11229_, _07570_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _42311_ (_11231_, _11229_, _11227_);
  and _42312_ (_11232_, _11231_, _07811_);
  or _42313_ (_11233_, _11232_, _11226_);
  and _42314_ (_11234_, _11233_, _07770_);
  nand _42315_ (_11235_, _07570_, _09293_);
  or _42316_ (_11237_, _07570_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _42317_ (_11238_, _11237_, _11235_);
  and _42318_ (_11239_, _11238_, _07812_);
  nand _42319_ (_11240_, _07570_, _09043_);
  or _42320_ (_11241_, _07570_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _42321_ (_11243_, _11241_, _11240_);
  and _42322_ (_11245_, _11243_, _07811_);
  or _42323_ (_11247_, _11245_, _11239_);
  and _42324_ (_11248_, _11247_, _07845_);
  nand _42325_ (_11249_, _07570_, _10298_);
  or _42326_ (_11250_, _07570_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _42327_ (_11251_, _11250_, _11249_);
  and _42328_ (_11253_, _11251_, _07812_);
  nand _42329_ (_11254_, _07570_, _10035_);
  or _42330_ (_11256_, _07570_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _42331_ (_11257_, _11256_, _11254_);
  and _42332_ (_11259_, _11257_, _07811_);
  or _42333_ (_11260_, _11259_, _11253_);
  and _42334_ (_11261_, _11260_, _07860_);
  or _42335_ (_11263_, _11261_, _11248_);
  or _42336_ (_11264_, _11263_, _11234_);
  nor _42337_ (_11266_, _11264_, _11221_);
  nor _42338_ (_11268_, _11266_, _07810_);
  or _42339_ (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _11268_, _11210_);
  and _42340_ (_11269_, _07471_, _23898_);
  and _42341_ (_11271_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  or _42342_ (_02972_, _11271_, _11269_);
  and _42343_ (_11272_, _07914_, word_in[16]);
  and _42344_ (_11274_, _10523_, _07591_);
  and _42345_ (_11275_, _10527_, _07624_);
  or _42346_ (_11276_, _11275_, _11274_);
  and _42347_ (_11277_, _10519_, _07597_);
  and _42348_ (_11278_, _10513_, _07608_);
  or _42349_ (_11279_, _11278_, _11277_);
  or _42350_ (_11281_, _11279_, _11276_);
  or _42351_ (_11282_, _11281_, _07881_);
  and _42352_ (_11283_, _10548_, _07624_);
  and _42353_ (_11284_, _10534_, _07608_);
  or _42354_ (_11285_, _11284_, _11283_);
  and _42355_ (_11287_, _10544_, _07591_);
  and _42356_ (_11288_, _10539_, _07597_);
  or _42357_ (_11290_, _11288_, _11287_);
  or _42358_ (_11291_, _11290_, _11285_);
  or _42359_ (_11292_, _11291_, _07915_);
  nand _42360_ (_11293_, _11292_, _11282_);
  nor _42361_ (_11294_, _11293_, _07914_);
  or _42362_ (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _11294_, _11272_);
  and _42363_ (_11295_, _07914_, word_in[17]);
  and _42364_ (_11297_, _10575_, _07624_);
  and _42365_ (_11298_, _10565_, _07597_);
  or _42366_ (_11300_, _11298_, _11297_);
  and _42367_ (_11301_, _10570_, _07591_);
  and _42368_ (_11302_, _10560_, _07608_);
  or _42369_ (_11303_, _11302_, _11301_);
  or _42370_ (_11304_, _11303_, _11300_);
  or _42371_ (_11305_, _11304_, _07881_);
  and _42372_ (_11306_, _10591_, _07591_);
  and _42373_ (_11308_, _10587_, _07597_);
  or _42374_ (_11309_, _11308_, _11306_);
  and _42375_ (_11310_, _10595_, _07624_);
  and _42376_ (_11311_, _10582_, _07608_);
  or _42377_ (_11313_, _11311_, _11310_);
  or _42378_ (_11314_, _11313_, _11309_);
  or _42379_ (_11316_, _11314_, _07915_);
  nand _42380_ (_11318_, _11316_, _11305_);
  nor _42381_ (_11320_, _11318_, _07914_);
  or _42382_ (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _11320_, _11295_);
  and _42383_ (_11321_, _07914_, word_in[18]);
  and _42384_ (_11323_, _10617_, _07591_);
  and _42385_ (_11324_, _10608_, _07624_);
  or _42386_ (_11325_, _11324_, _11323_);
  and _42387_ (_11326_, _10613_, _07597_);
  and _42388_ (_11327_, _10621_, _07608_);
  or _42389_ (_11328_, _11327_, _11326_);
  or _42390_ (_11330_, _11328_, _11325_);
  or _42391_ (_11332_, _11330_, _07881_);
  and _42392_ (_11333_, _10631_, _07624_);
  and _42393_ (_11334_, _10640_, _07597_);
  or _42394_ (_11336_, _11334_, _11333_);
  and _42395_ (_11337_, _10636_, _07591_);
  and _42396_ (_11338_, _10647_, _07608_);
  or _42397_ (_11339_, _11338_, _11337_);
  or _42398_ (_11340_, _11339_, _11336_);
  or _42399_ (_11342_, _11340_, _07915_);
  nand _42400_ (_11343_, _11342_, _11332_);
  nor _42401_ (_11344_, _11343_, _07914_);
  or _42402_ (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _11344_, _11321_);
  and _42403_ (_11345_, _07914_, word_in[19]);
  and _42404_ (_11347_, _10659_, _07624_);
  and _42405_ (_11348_, _10665_, _07597_);
  or _42406_ (_11350_, _11348_, _11347_);
  and _42407_ (_11351_, _10669_, _07591_);
  and _42408_ (_11352_, _10673_, _07608_);
  or _42409_ (_11354_, _11352_, _11351_);
  or _42410_ (_11355_, _11354_, _11350_);
  or _42411_ (_11357_, _11355_, _07881_);
  and _42412_ (_11359_, _10682_, _07624_);
  and _42413_ (_11360_, _10691_, _07597_);
  or _42414_ (_11361_, _11360_, _11359_);
  and _42415_ (_11362_, _10687_, _07591_);
  and _42416_ (_11363_, _10696_, _07608_);
  or _42417_ (_11365_, _11363_, _11362_);
  or _42418_ (_11366_, _11365_, _11361_);
  or _42419_ (_11367_, _11366_, _07915_);
  nand _42420_ (_11369_, _11367_, _11357_);
  nor _42421_ (_11370_, _11369_, _07914_);
  or _42422_ (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _11370_, _11345_);
  and _42423_ (_11371_, _07914_, word_in[20]);
  and _42424_ (_11372_, _10722_, _07624_);
  and _42425_ (_11373_, _10713_, _07597_);
  or _42426_ (_11375_, _11373_, _11372_);
  and _42427_ (_11377_, _10717_, _07591_);
  and _42428_ (_11378_, _10707_, _07608_);
  or _42429_ (_11379_, _11378_, _11377_);
  or _42430_ (_11380_, _11379_, _11375_);
  or _42431_ (_11381_, _11380_, _07881_);
  and _42432_ (_11382_, _10741_, _07591_);
  and _42433_ (_11383_, _10747_, _07624_);
  or _42434_ (_11384_, _11383_, _11382_);
  and _42435_ (_11385_, _10736_, _07597_);
  and _42436_ (_11386_, _10729_, _07608_);
  or _42437_ (_11387_, _11386_, _11385_);
  or _42438_ (_11389_, _11387_, _11384_);
  or _42439_ (_11390_, _11389_, _07915_);
  nand _42440_ (_11391_, _11390_, _11381_);
  nor _42441_ (_11392_, _11391_, _07914_);
  or _42442_ (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _11392_, _11371_);
  and _42443_ (_11393_, _07914_, word_in[21]);
  and _42444_ (_11395_, _10766_, _07597_);
  and _42445_ (_11397_, _10761_, _07608_);
  or _42446_ (_11398_, _11397_, _11395_);
  and _42447_ (_11399_, _10771_, _07591_);
  and _42448_ (_11401_, _10776_, _07624_);
  or _42449_ (_11402_, _11401_, _11399_);
  or _42450_ (_11403_, _11402_, _11398_);
  or _42451_ (_11405_, _11403_, _07881_);
  and _42452_ (_11407_, _10793_, _07597_);
  and _42453_ (_11409_, _10786_, _07608_);
  or _42454_ (_11411_, _11409_, _11407_);
  and _42455_ (_11412_, _10798_, _07591_);
  and _42456_ (_11415_, _10803_, _07624_);
  or _42457_ (_11416_, _11415_, _11412_);
  or _42458_ (_11417_, _11416_, _11411_);
  or _42459_ (_11419_, _11417_, _07915_);
  nand _42460_ (_11420_, _11419_, _11405_);
  nor _42461_ (_11421_, _11420_, _07914_);
  or _42462_ (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _11421_, _11393_);
  and _42463_ (_11422_, _07914_, word_in[22]);
  and _42464_ (_11423_, _10825_, _07591_);
  and _42465_ (_11424_, _10816_, _07624_);
  or _42466_ (_11426_, _11424_, _11423_);
  and _42467_ (_11427_, _10821_, _07597_);
  and _42468_ (_11428_, _10833_, _07608_);
  or _42469_ (_11429_, _11428_, _11427_);
  or _42470_ (_11430_, _11429_, _11426_);
  or _42471_ (_11431_, _11430_, _07881_);
  and _42472_ (_11432_, _10848_, _07591_);
  and _42473_ (_11433_, _10842_, _07624_);
  or _42474_ (_11434_, _11433_, _11432_);
  and _42475_ (_11435_, _10852_, _07597_);
  and _42476_ (_11436_, _10859_, _07608_);
  or _42477_ (_11437_, _11436_, _11435_);
  or _42478_ (_11438_, _11437_, _11434_);
  or _42479_ (_11439_, _11438_, _07915_);
  nand _42480_ (_11440_, _11439_, _11431_);
  nor _42481_ (_11441_, _11440_, _07914_);
  or _42482_ (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _11441_, _11422_);
  and _42483_ (_11442_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  and _42484_ (_11443_, _10494_, _23707_);
  or _42485_ (_02996_, _11443_, _11442_);
  and _42486_ (_11444_, _07975_, word_in[24]);
  and _42487_ (_11445_, _10877_, _07812_);
  and _42488_ (_11446_, _10871_, _07811_);
  or _42489_ (_11447_, _11446_, _11445_);
  and _42490_ (_11448_, _11447_, _07949_);
  and _42491_ (_11449_, _10890_, _07812_);
  and _42492_ (_11450_, _10884_, _07811_);
  or _42493_ (_11451_, _11450_, _11449_);
  and _42494_ (_11452_, _11451_, _07951_);
  and _42495_ (_11453_, _10905_, _07812_);
  and _42496_ (_11455_, _10900_, _07811_);
  or _42497_ (_11457_, _11455_, _11453_);
  and _42498_ (_11459_, _11457_, _07984_);
  and _42499_ (_11461_, _10916_, _07812_);
  and _42500_ (_11462_, _10911_, _07811_);
  or _42501_ (_11464_, _11462_, _11461_);
  and _42502_ (_11465_, _11464_, _07992_);
  or _42503_ (_11466_, _11465_, _11459_);
  or _42504_ (_11467_, _11466_, _11452_);
  nor _42505_ (_11469_, _11467_, _11448_);
  nor _42506_ (_11470_, _11469_, _07975_);
  or _42507_ (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _11470_, _11444_);
  and _42508_ (_11472_, _07975_, word_in[25]);
  and _42509_ (_11474_, _10934_, _07812_);
  and _42510_ (_11475_, _10929_, _07811_);
  or _42511_ (_11476_, _11475_, _11474_);
  and _42512_ (_11477_, _11476_, _07949_);
  and _42513_ (_11479_, _10948_, _07812_);
  and _42514_ (_11480_, _10942_, _07811_);
  or _42515_ (_11481_, _11480_, _11479_);
  and _42516_ (_11484_, _11481_, _07951_);
  and _42517_ (_11486_, _10962_, _07812_);
  and _42518_ (_11488_, _10956_, _07811_);
  or _42519_ (_11490_, _11488_, _11486_);
  and _42520_ (_11492_, _11490_, _07984_);
  and _42521_ (_11494_, _10976_, _07812_);
  and _42522_ (_11495_, _10970_, _07811_);
  or _42523_ (_11496_, _11495_, _11494_);
  and _42524_ (_11498_, _11496_, _07992_);
  or _42525_ (_11500_, _11498_, _11492_);
  or _42526_ (_11501_, _11500_, _11484_);
  nor _42527_ (_11503_, _11501_, _11477_);
  nor _42528_ (_11504_, _11503_, _07975_);
  or _42529_ (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _11504_, _11472_);
  and _42530_ (_11507_, _07975_, word_in[26]);
  and _42531_ (_11508_, _10993_, _07812_);
  and _42532_ (_11509_, _10989_, _07811_);
  or _42533_ (_11511_, _11509_, _11508_);
  and _42534_ (_11513_, _11511_, _07949_);
  and _42535_ (_11514_, _11003_, _07812_);
  and _42536_ (_11516_, _10999_, _07811_);
  or _42537_ (_11517_, _11516_, _11514_);
  and _42538_ (_11518_, _11517_, _07951_);
  and _42539_ (_11520_, _11013_, _07812_);
  and _42540_ (_11521_, _11009_, _07811_);
  or _42541_ (_11523_, _11521_, _11520_);
  and _42542_ (_11525_, _11523_, _07984_);
  and _42543_ (_11527_, _11023_, _07812_);
  and _42544_ (_11529_, _11019_, _07811_);
  or _42545_ (_11530_, _11529_, _11527_);
  and _42546_ (_11531_, _11530_, _07992_);
  or _42547_ (_11533_, _11531_, _11525_);
  or _42548_ (_11535_, _11533_, _11518_);
  nor _42549_ (_11536_, _11535_, _11513_);
  nor _42550_ (_11537_, _11536_, _07975_);
  or _42551_ (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _11537_, _11507_);
  and _42552_ (_11540_, _07975_, word_in[27]);
  and _42553_ (_11542_, _11038_, _07812_);
  and _42554_ (_11544_, _11034_, _07811_);
  or _42555_ (_11546_, _11544_, _11542_);
  and _42556_ (_11547_, _11546_, _07949_);
  and _42557_ (_11549_, _11048_, _07812_);
  and _42558_ (_11550_, _11044_, _07811_);
  or _42559_ (_11551_, _11550_, _11549_);
  and _42560_ (_11552_, _11551_, _07951_);
  and _42561_ (_11553_, _11061_, _07812_);
  and _42562_ (_11554_, _11056_, _07811_);
  or _42563_ (_11555_, _11554_, _11553_);
  and _42564_ (_11556_, _11555_, _07984_);
  and _42565_ (_11557_, _11073_, _07812_);
  and _42566_ (_11559_, _11068_, _07811_);
  or _42567_ (_11560_, _11559_, _11557_);
  and _42568_ (_11561_, _11560_, _07992_);
  or _42569_ (_11563_, _11561_, _11556_);
  or _42570_ (_11564_, _11563_, _11552_);
  nor _42571_ (_11566_, _11564_, _11547_);
  nor _42572_ (_11567_, _11566_, _07975_);
  or _42573_ (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _11567_, _11540_);
  and _42574_ (_11570_, _07975_, word_in[28]);
  and _42575_ (_11571_, _11097_, _07812_);
  and _42576_ (_11572_, _11090_, _07811_);
  or _42577_ (_11573_, _11572_, _11571_);
  and _42578_ (_11574_, _11573_, _07949_);
  and _42579_ (_11575_, _11113_, _07812_);
  and _42580_ (_11576_, _11107_, _07811_);
  or _42581_ (_11578_, _11576_, _11575_);
  and _42582_ (_11579_, _11578_, _07951_);
  and _42583_ (_11580_, _11126_, _07812_);
  and _42584_ (_11581_, _11121_, _07811_);
  or _42585_ (_11582_, _11581_, _11580_);
  and _42586_ (_11584_, _11582_, _07984_);
  and _42587_ (_11585_, _11142_, _07812_);
  and _42588_ (_11586_, _11135_, _07811_);
  or _42589_ (_11587_, _11586_, _11585_);
  and _42590_ (_11588_, _11587_, _07992_);
  or _42591_ (_11589_, _11588_, _11584_);
  or _42592_ (_11590_, _11589_, _11579_);
  nor _42593_ (_11592_, _11590_, _11574_);
  nor _42594_ (_11593_, _11592_, _07975_);
  or _42595_ (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _11593_, _11570_);
  and _42596_ (_11594_, _07975_, word_in[29]);
  and _42597_ (_11596_, _11163_, _07812_);
  and _42598_ (_11597_, _11157_, _07811_);
  or _42599_ (_11598_, _11597_, _11596_);
  and _42600_ (_11599_, _11598_, _07949_);
  and _42601_ (_11600_, _11174_, _07812_);
  and _42602_ (_11601_, _11170_, _07811_);
  or _42603_ (_11602_, _11601_, _11600_);
  and _42604_ (_11603_, _11602_, _07951_);
  and _42605_ (_11605_, _11186_, _07812_);
  and _42606_ (_11606_, _11181_, _07811_);
  or _42607_ (_11607_, _11606_, _11605_);
  and _42608_ (_11608_, _11607_, _07984_);
  and _42609_ (_11610_, _11199_, _07812_);
  and _42610_ (_11611_, _11194_, _07811_);
  or _42611_ (_11612_, _11611_, _11610_);
  and _42612_ (_11614_, _11612_, _07992_);
  or _42613_ (_11616_, _11614_, _11608_);
  or _42614_ (_11618_, _11616_, _11603_);
  nor _42615_ (_11619_, _11618_, _11599_);
  nor _42616_ (_11620_, _11619_, _07975_);
  or _42617_ (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _11620_, _11594_);
  and _42618_ (_11623_, _07975_, word_in[30]);
  and _42619_ (_11624_, _11231_, _07812_);
  and _42620_ (_11626_, _11225_, _07811_);
  or _42621_ (_11627_, _11626_, _11624_);
  and _42622_ (_11629_, _11627_, _07951_);
  and _42623_ (_11630_, _11218_, _07812_);
  and _42624_ (_11631_, _11213_, _07811_);
  or _42625_ (_11632_, _11631_, _11630_);
  and _42626_ (_11633_, _11632_, _07949_);
  and _42627_ (_11634_, _11243_, _07812_);
  and _42628_ (_11635_, _11238_, _07811_);
  or _42629_ (_11636_, _11635_, _11634_);
  and _42630_ (_11638_, _11636_, _07984_);
  and _42631_ (_11639_, _11257_, _07812_);
  and _42632_ (_11640_, _11251_, _07811_);
  or _42633_ (_11641_, _11640_, _11639_);
  and _42634_ (_11642_, _11641_, _07992_);
  or _42635_ (_11644_, _11642_, _11638_);
  or _42636_ (_11646_, _11644_, _11633_);
  nor _42637_ (_11647_, _11646_, _11629_);
  nor _42638_ (_11648_, _11647_, _07975_);
  or _42639_ (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _11648_, _11623_);
  and _42640_ (_11649_, _05445_, _23707_);
  and _42641_ (_11650_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  or _42642_ (_03046_, _11650_, _11649_);
  and _42643_ (_11652_, _25078_, _24766_);
  not _42644_ (_11653_, _11652_);
  and _42645_ (_11654_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and _42646_ (_11655_, _11652_, _23778_);
  or _42647_ (_03052_, _11655_, _11654_);
  and _42648_ (_11657_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and _42649_ (_11658_, _11652_, _23824_);
  or _42650_ (_03069_, _11658_, _11657_);
  and _42651_ (_11660_, _05445_, _23824_);
  and _42652_ (_11661_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  or _42653_ (_03108_, _11661_, _11660_);
  and _42654_ (_11664_, _02374_, _23778_);
  and _42655_ (_11666_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  or _42656_ (_03114_, _11666_, _11664_);
  and _42657_ (_11667_, _24086_, _23898_);
  and _42658_ (_11668_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or _42659_ (_03117_, _11668_, _11667_);
  and _42660_ (_11669_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and _42661_ (_11670_, _11652_, _23747_);
  or _42662_ (_03123_, _11670_, _11669_);
  and _42663_ (_11671_, _07536_, _23946_);
  and _42664_ (_11672_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  or _42665_ (_03125_, _11672_, _11671_);
  and _42666_ (_11673_, _07536_, _23898_);
  and _42667_ (_11674_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  or _42668_ (_03129_, _11674_, _11673_);
  and _42669_ (_11675_, _07536_, _23747_);
  and _42670_ (_11676_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  or _42671_ (_03139_, _11676_, _11675_);
  and _42672_ (_11678_, _02345_, _23824_);
  and _42673_ (_11679_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or _42674_ (_27191_, _11679_, _11678_);
  and _42675_ (_11680_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and _42676_ (_11682_, _11652_, _24050_);
  or _42677_ (_03144_, _11682_, _11680_);
  nor _42678_ (_26887_[1], _00094_, rst);
  and _42679_ (_11685_, _05180_, _23824_);
  and _42680_ (_11686_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or _42681_ (_03160_, _11686_, _11685_);
  and _42682_ (_11688_, _08167_, _23747_);
  and _42683_ (_11689_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  or _42684_ (_03164_, _11689_, _11688_);
  and _42685_ (_11691_, _10347_, _23707_);
  and _42686_ (_11692_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  or _42687_ (_03168_, _11692_, _11691_);
  and _42688_ (_11693_, _24766_, _23656_);
  not _42689_ (_11695_, _11693_);
  and _42690_ (_11697_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and _42691_ (_11699_, _11693_, _23898_);
  or _42692_ (_03175_, _11699_, _11697_);
  and _42693_ (_11700_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and _42694_ (_11701_, _11693_, _23747_);
  or _42695_ (_03177_, _11701_, _11700_);
  and _42696_ (_11702_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and _42697_ (_11703_, _11693_, _23946_);
  or _42698_ (_03194_, _11703_, _11702_);
  and _42699_ (_11705_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and _42700_ (_11706_, _11693_, _23707_);
  or _42701_ (_03199_, _11706_, _11705_);
  and _42702_ (_11708_, _02284_, _23898_);
  and _42703_ (_11709_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  or _42704_ (_27116_, _11709_, _11708_);
  and _42705_ (_11712_, _04811_, _23898_);
  and _42706_ (_11713_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  or _42707_ (_03209_, _11713_, _11712_);
  and _42708_ (_11714_, _02302_, _24050_);
  and _42709_ (_11716_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or _42710_ (_03211_, _11716_, _11714_);
  and _42711_ (_11717_, _02302_, _23824_);
  and _42712_ (_11719_, _02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or _42713_ (_03222_, _11719_, _11717_);
  and _42714_ (_11720_, _02374_, _23707_);
  and _42715_ (_11722_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  or _42716_ (_03225_, _11722_, _11720_);
  and _42717_ (_11725_, _03339_, _23946_);
  and _42718_ (_11727_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or _42719_ (_03227_, _11727_, _11725_);
  and _42720_ (_11729_, _24766_, _23752_);
  not _42721_ (_11730_, _11729_);
  and _42722_ (_11731_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  and _42723_ (_11732_, _11729_, _23778_);
  or _42724_ (_03231_, _11732_, _11731_);
  and _42725_ (_11735_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  and _42726_ (_11736_, _11729_, _23824_);
  or _42727_ (_03233_, _11736_, _11735_);
  and _42728_ (_11737_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  and _42729_ (_11739_, _11729_, _23946_);
  or _42730_ (_03244_, _11739_, _11737_);
  and _42731_ (_11740_, _04917_, _24050_);
  and _42732_ (_11741_, _04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or _42733_ (_27110_, _11741_, _11740_);
  and _42734_ (_11742_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  and _42735_ (_11743_, _11729_, _24050_);
  or _42736_ (_27026_, _11743_, _11742_);
  and _42737_ (_11744_, _07471_, _23747_);
  and _42738_ (_11745_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  or _42739_ (_03270_, _11745_, _11744_);
  and _42740_ (_11746_, _24766_, _24329_);
  not _42741_ (_11747_, _11746_);
  and _42742_ (_11748_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and _42743_ (_11749_, _11746_, _23778_);
  or _42744_ (_03282_, _11749_, _11748_);
  and _42745_ (_11750_, _05445_, _23649_);
  and _42746_ (_11751_, _05447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  or _42747_ (_03287_, _11751_, _11750_);
  and _42748_ (_11752_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and _42749_ (_11753_, _11746_, _23898_);
  or _42750_ (_03289_, _11753_, _11752_);
  and _42751_ (_11756_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and _42752_ (_11757_, _11746_, _23649_);
  or _42753_ (_03291_, _11757_, _11756_);
  and _42754_ (_11760_, _02374_, _23824_);
  and _42755_ (_11761_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  or _42756_ (_03294_, _11761_, _11760_);
  and _42757_ (_11763_, _09913_, _23946_);
  and _42758_ (_11764_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or _42759_ (_03304_, _11764_, _11763_);
  and _42760_ (_11765_, _07536_, _23707_);
  and _42761_ (_11766_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  or _42762_ (_03310_, _11766_, _11765_);
  and _42763_ (_11767_, _05180_, _24050_);
  and _42764_ (_11768_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or _42765_ (_27133_, _11768_, _11767_);
  and _42766_ (_11769_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and _42767_ (_11770_, _11746_, _23946_);
  or _42768_ (_03326_, _11770_, _11769_);
  and _42769_ (_11771_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and _42770_ (_11772_, _11746_, _23707_);
  or _42771_ (_27030_, _11772_, _11771_);
  and _42772_ (_11773_, _08167_, _23707_);
  and _42773_ (_11774_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or _42774_ (_03333_, _11774_, _11773_);
  and _42775_ (_11775_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  and _42776_ (_11776_, _04748_, _23778_);
  or _42777_ (_03341_, _11776_, _11775_);
  and _42778_ (_11777_, _10347_, _23778_);
  and _42779_ (_11778_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  or _42780_ (_03346_, _11778_, _11777_);
  and _42781_ (_11779_, _04797_, _23778_);
  and _42782_ (_11780_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or _42783_ (_03357_, _11780_, _11779_);
  and _42784_ (_11781_, _01810_, _23898_);
  and _42785_ (_11782_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or _42786_ (_03362_, _11782_, _11781_);
  and _42787_ (_11784_, _24371_, _23649_);
  and _42788_ (_11785_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or _42789_ (_03365_, _11785_, _11784_);
  and _42790_ (_11786_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  and _42791_ (_11788_, _06888_, _23707_);
  or _42792_ (_03371_, _11788_, _11786_);
  and _42793_ (_11789_, _07471_, _23707_);
  and _42794_ (_11790_, _07473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or _42795_ (_03391_, _11790_, _11789_);
  and _42796_ (_11794_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  and _42797_ (_11796_, _06888_, _24050_);
  or _42798_ (_03398_, _11796_, _11794_);
  and _42799_ (_11798_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and _42800_ (_11799_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or _42801_ (_11800_, _11799_, _11798_);
  and _42802_ (_11801_, _11800_, _02445_);
  and _42803_ (_11802_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and _42804_ (_11804_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or _42805_ (_11805_, _11804_, _11802_);
  and _42806_ (_11806_, _11805_, _02393_);
  or _42807_ (_11807_, _11806_, _11801_);
  or _42808_ (_11808_, _11807_, _02459_);
  and _42809_ (_11809_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and _42810_ (_11810_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or _42811_ (_11811_, _11810_, _11809_);
  and _42812_ (_11812_, _11811_, _02445_);
  and _42813_ (_11813_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and _42814_ (_11814_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or _42815_ (_11815_, _11814_, _11813_);
  and _42816_ (_11816_, _11815_, _02393_);
  or _42817_ (_11818_, _11816_, _11812_);
  or _42818_ (_11819_, _11818_, _02421_);
  and _42819_ (_11820_, _11819_, _02458_);
  and _42820_ (_11821_, _11820_, _11808_);
  or _42821_ (_11822_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or _42822_ (_11823_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and _42823_ (_11824_, _11823_, _02393_);
  and _42824_ (_11825_, _11824_, _11822_);
  or _42825_ (_11826_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or _42826_ (_11827_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and _42827_ (_11829_, _11827_, _02445_);
  and _42828_ (_11831_, _11829_, _11826_);
  or _42829_ (_11832_, _11831_, _11825_);
  or _42830_ (_11833_, _11832_, _02459_);
  or _42831_ (_11835_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or _42832_ (_11836_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and _42833_ (_11837_, _11836_, _02393_);
  and _42834_ (_11838_, _11837_, _11835_);
  or _42835_ (_11839_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or _42836_ (_11840_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and _42837_ (_11841_, _11840_, _02445_);
  and _42838_ (_11842_, _11841_, _11839_);
  or _42839_ (_11843_, _11842_, _11838_);
  or _42840_ (_11844_, _11843_, _02421_);
  and _42841_ (_11845_, _11844_, _02414_);
  and _42842_ (_11846_, _11845_, _11833_);
  or _42843_ (_11847_, _11846_, _11821_);
  or _42844_ (_11848_, _11847_, _02398_);
  and _42845_ (_11850_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and _42846_ (_11851_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or _42847_ (_11852_, _11851_, _02393_);
  or _42848_ (_11854_, _11852_, _11850_);
  and _42849_ (_11856_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and _42850_ (_11858_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or _42851_ (_11860_, _11858_, _02445_);
  or _42852_ (_11861_, _11860_, _11856_);
  and _42853_ (_11862_, _11861_, _11854_);
  or _42854_ (_11864_, _11862_, _02459_);
  and _42855_ (_11865_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and _42856_ (_11866_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or _42857_ (_11868_, _11866_, _02393_);
  or _42858_ (_11869_, _11868_, _11865_);
  and _42859_ (_11870_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and _42860_ (_11871_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or _42861_ (_11873_, _11871_, _02445_);
  or _42862_ (_11874_, _11873_, _11870_);
  and _42863_ (_11875_, _11874_, _11869_);
  or _42864_ (_11876_, _11875_, _02421_);
  and _42865_ (_11877_, _11876_, _02458_);
  and _42866_ (_11879_, _11877_, _11864_);
  or _42867_ (_11880_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or _42868_ (_11881_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and _42869_ (_11883_, _11881_, _11880_);
  or _42870_ (_11885_, _11883_, _02445_);
  or _42871_ (_11886_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or _42872_ (_11887_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and _42873_ (_11888_, _11887_, _11886_);
  or _42874_ (_11889_, _11888_, _02393_);
  and _42875_ (_11890_, _11889_, _11885_);
  or _42876_ (_11892_, _11890_, _02459_);
  or _42877_ (_11893_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or _42878_ (_11894_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and _42879_ (_11895_, _11894_, _11893_);
  or _42880_ (_11896_, _11895_, _02445_);
  or _42881_ (_11897_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or _42882_ (_11898_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and _42883_ (_11899_, _11898_, _11897_);
  or _42884_ (_11900_, _11899_, _02393_);
  and _42885_ (_11901_, _11900_, _11896_);
  or _42886_ (_11902_, _11901_, _02421_);
  and _42887_ (_11903_, _11902_, _02414_);
  and _42888_ (_11904_, _11903_, _11892_);
  or _42889_ (_11905_, _11904_, _11879_);
  or _42890_ (_11906_, _11905_, _02496_);
  and _42891_ (_11907_, _11906_, _02546_);
  and _42892_ (_11908_, _11907_, _11848_);
  and _42893_ (_11909_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and _42894_ (_11910_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or _42895_ (_11912_, _11910_, _11909_);
  and _42896_ (_11913_, _11912_, _02393_);
  and _42897_ (_11914_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and _42898_ (_11915_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or _42899_ (_11916_, _11915_, _11914_);
  and _42900_ (_11917_, _11916_, _02445_);
  or _42901_ (_11918_, _11917_, _11913_);
  and _42902_ (_11919_, _11918_, _02421_);
  and _42903_ (_11920_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and _42904_ (_11921_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or _42905_ (_11922_, _11921_, _11920_);
  and _42906_ (_11923_, _11922_, _02393_);
  and _42907_ (_11925_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and _42908_ (_11926_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or _42909_ (_11927_, _11926_, _11925_);
  and _42910_ (_11928_, _11927_, _02445_);
  or _42911_ (_11929_, _11928_, _11923_);
  and _42912_ (_11930_, _11929_, _02459_);
  or _42913_ (_11931_, _11930_, _11919_);
  and _42914_ (_11932_, _11931_, _02458_);
  or _42915_ (_11933_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or _42916_ (_11934_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and _42917_ (_11935_, _11934_, _11933_);
  and _42918_ (_11936_, _11935_, _02393_);
  or _42919_ (_11937_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or _42920_ (_11938_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and _42921_ (_11939_, _11938_, _11937_);
  and _42922_ (_11940_, _11939_, _02445_);
  or _42923_ (_11941_, _11940_, _11936_);
  and _42924_ (_11942_, _11941_, _02421_);
  or _42925_ (_11943_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or _42926_ (_11944_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and _42927_ (_11945_, _11944_, _11943_);
  and _42928_ (_11946_, _11945_, _02393_);
  or _42929_ (_11947_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or _42930_ (_11948_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and _42931_ (_11949_, _11948_, _11947_);
  and _42932_ (_11950_, _11949_, _02445_);
  or _42933_ (_11951_, _11950_, _11946_);
  and _42934_ (_11952_, _11951_, _02459_);
  or _42935_ (_11953_, _11952_, _11942_);
  and _42936_ (_11955_, _11953_, _02414_);
  or _42937_ (_11956_, _11955_, _11932_);
  and _42938_ (_11957_, _11956_, _02398_);
  and _42939_ (_11958_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  and _42940_ (_11959_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  or _42941_ (_11960_, _11959_, _11958_);
  and _42942_ (_11961_, _11960_, _02393_);
  and _42943_ (_11963_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  and _42944_ (_11965_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  or _42945_ (_11966_, _11965_, _11963_);
  and _42946_ (_11967_, _11966_, _02445_);
  or _42947_ (_11968_, _11967_, _11961_);
  and _42948_ (_11969_, _11968_, _02421_);
  and _42949_ (_11970_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  and _42950_ (_11971_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  or _42951_ (_11972_, _11971_, _11970_);
  and _42952_ (_11973_, _11972_, _02393_);
  and _42953_ (_11974_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  and _42954_ (_11975_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  or _42955_ (_11976_, _11975_, _11974_);
  and _42956_ (_11977_, _11976_, _02445_);
  or _42957_ (_11978_, _11977_, _11973_);
  and _42958_ (_11979_, _11978_, _02459_);
  or _42959_ (_11980_, _11979_, _11969_);
  and _42960_ (_11981_, _11980_, _02458_);
  or _42961_ (_11982_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  or _42962_ (_11983_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  and _42963_ (_11984_, _11983_, _11982_);
  and _42964_ (_11985_, _11984_, _02393_);
  or _42965_ (_11986_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  or _42966_ (_11988_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  and _42967_ (_11989_, _11988_, _11986_);
  and _42968_ (_11990_, _11989_, _02445_);
  or _42969_ (_11991_, _11990_, _11985_);
  and _42970_ (_11992_, _11991_, _02421_);
  or _42971_ (_11993_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  or _42972_ (_11994_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  and _42973_ (_11995_, _11994_, _11993_);
  and _42974_ (_11996_, _11995_, _02393_);
  or _42975_ (_11997_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  or _42976_ (_11999_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  and _42977_ (_12000_, _11999_, _11997_);
  and _42978_ (_12001_, _12000_, _02445_);
  or _42979_ (_12003_, _12001_, _11996_);
  and _42980_ (_12004_, _12003_, _02459_);
  or _42981_ (_12005_, _12004_, _11992_);
  and _42982_ (_12006_, _12005_, _02414_);
  or _42983_ (_12007_, _12006_, _11981_);
  and _42984_ (_12008_, _12007_, _02496_);
  or _42985_ (_12010_, _12008_, _11957_);
  and _42986_ (_12011_, _12010_, _02400_);
  or _42987_ (_12012_, _12011_, _11908_);
  and _42988_ (_12013_, _12012_, _02646_);
  or _42989_ (_12014_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or _42990_ (_12015_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and _42991_ (_12016_, _12015_, _02445_);
  and _42992_ (_12017_, _12016_, _12014_);
  or _42993_ (_12018_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or _42994_ (_12019_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and _42995_ (_12020_, _12019_, _02393_);
  and _42996_ (_12021_, _12020_, _12018_);
  or _42997_ (_12023_, _12021_, _12017_);
  and _42998_ (_12025_, _12023_, _02459_);
  or _42999_ (_12027_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or _43000_ (_12029_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and _43001_ (_12030_, _12029_, _02445_);
  and _43002_ (_12031_, _12030_, _12027_);
  or _43003_ (_12032_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or _43004_ (_12033_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and _43005_ (_12034_, _12033_, _02393_);
  and _43006_ (_12036_, _12034_, _12032_);
  or _43007_ (_12038_, _12036_, _12031_);
  and _43008_ (_12039_, _12038_, _02421_);
  or _43009_ (_12041_, _12039_, _12025_);
  and _43010_ (_12043_, _12041_, _02414_);
  and _43011_ (_12045_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and _43012_ (_12046_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or _43013_ (_12047_, _12046_, _12045_);
  and _43014_ (_12049_, _12047_, _02393_);
  and _43015_ (_12051_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and _43016_ (_12053_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or _43017_ (_12055_, _12053_, _12051_);
  and _43018_ (_12057_, _12055_, _02445_);
  or _43019_ (_12058_, _12057_, _12049_);
  and _43020_ (_12059_, _12058_, _02459_);
  and _43021_ (_12061_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and _43022_ (_12062_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or _43023_ (_12064_, _12062_, _12061_);
  and _43024_ (_12065_, _12064_, _02393_);
  and _43025_ (_12067_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and _43026_ (_12069_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or _43027_ (_12071_, _12069_, _12067_);
  and _43028_ (_12073_, _12071_, _02445_);
  or _43029_ (_12074_, _12073_, _12065_);
  and _43030_ (_12075_, _12074_, _02421_);
  or _43031_ (_12076_, _12075_, _12059_);
  and _43032_ (_12077_, _12076_, _02458_);
  or _43033_ (_12078_, _12077_, _12043_);
  and _43034_ (_12079_, _12078_, _02496_);
  or _43035_ (_12080_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or _43036_ (_12081_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and _43037_ (_12082_, _12081_, _12080_);
  and _43038_ (_12083_, _12082_, _02393_);
  or _43039_ (_12084_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or _43040_ (_12085_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and _43041_ (_12087_, _12085_, _12084_);
  and _43042_ (_12088_, _12087_, _02445_);
  or _43043_ (_12089_, _12088_, _12083_);
  and _43044_ (_12090_, _12089_, _02459_);
  or _43045_ (_12091_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or _43046_ (_12092_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and _43047_ (_12093_, _12092_, _12091_);
  and _43048_ (_12094_, _12093_, _02393_);
  or _43049_ (_12095_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or _43050_ (_12096_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and _43051_ (_12097_, _12096_, _12095_);
  and _43052_ (_12098_, _12097_, _02445_);
  or _43053_ (_12099_, _12098_, _12094_);
  and _43054_ (_12100_, _12099_, _02421_);
  or _43055_ (_12102_, _12100_, _12090_);
  and _43056_ (_12103_, _12102_, _02414_);
  and _43057_ (_12104_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and _43058_ (_12106_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or _43059_ (_12108_, _12106_, _12104_);
  and _43060_ (_12110_, _12108_, _02393_);
  and _43061_ (_12112_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and _43062_ (_12114_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or _43063_ (_12115_, _12114_, _12112_);
  and _43064_ (_12117_, _12115_, _02445_);
  or _43065_ (_12118_, _12117_, _12110_);
  and _43066_ (_12119_, _12118_, _02459_);
  and _43067_ (_12120_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and _43068_ (_12121_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or _43069_ (_12122_, _12121_, _12120_);
  and _43070_ (_12123_, _12122_, _02393_);
  and _43071_ (_12124_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and _43072_ (_12125_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or _43073_ (_12126_, _12125_, _12124_);
  and _43074_ (_12127_, _12126_, _02445_);
  or _43075_ (_12128_, _12127_, _12123_);
  and _43076_ (_12129_, _12128_, _02421_);
  or _43077_ (_12130_, _12129_, _12119_);
  and _43078_ (_12131_, _12130_, _02458_);
  or _43079_ (_12132_, _12131_, _12103_);
  and _43080_ (_12133_, _12132_, _02398_);
  or _43081_ (_12134_, _12133_, _12079_);
  and _43082_ (_12135_, _12134_, _02400_);
  and _43083_ (_12136_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and _43084_ (_12137_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or _43085_ (_12138_, _12137_, _12136_);
  and _43086_ (_12140_, _12138_, _02393_);
  and _43087_ (_12141_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and _43088_ (_12142_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or _43089_ (_12143_, _12142_, _12141_);
  and _43090_ (_12144_, _12143_, _02445_);
  or _43091_ (_12145_, _12144_, _12140_);
  or _43092_ (_12146_, _12145_, _02459_);
  and _43093_ (_12147_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and _43094_ (_12148_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or _43095_ (_12149_, _12148_, _12147_);
  and _43096_ (_12150_, _12149_, _02393_);
  and _43097_ (_12151_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and _43098_ (_12152_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or _43099_ (_12153_, _12152_, _12151_);
  and _43100_ (_12154_, _12153_, _02445_);
  or _43101_ (_12155_, _12154_, _12150_);
  or _43102_ (_12156_, _12155_, _02421_);
  and _43103_ (_12157_, _12156_, _02458_);
  and _43104_ (_12158_, _12157_, _12146_);
  or _43105_ (_12159_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or _43106_ (_12160_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and _43107_ (_12161_, _12160_, _12159_);
  and _43108_ (_12162_, _12161_, _02393_);
  or _43109_ (_12163_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or _43110_ (_12164_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and _43111_ (_12165_, _12164_, _12163_);
  and _43112_ (_12166_, _12165_, _02445_);
  or _43113_ (_12167_, _12166_, _12162_);
  or _43114_ (_12168_, _12167_, _02459_);
  or _43115_ (_12169_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or _43116_ (_12171_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and _43117_ (_12172_, _12171_, _12169_);
  and _43118_ (_12173_, _12172_, _02393_);
  or _43119_ (_12174_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or _43120_ (_12175_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and _43121_ (_12176_, _12175_, _12174_);
  and _43122_ (_12177_, _12176_, _02445_);
  or _43123_ (_12178_, _12177_, _12173_);
  or _43124_ (_12179_, _12178_, _02421_);
  and _43125_ (_12180_, _12179_, _02414_);
  and _43126_ (_12181_, _12180_, _12168_);
  or _43127_ (_12182_, _12181_, _12158_);
  and _43128_ (_12183_, _12182_, _02398_);
  and _43129_ (_12184_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and _43130_ (_12186_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or _43131_ (_12187_, _12186_, _12184_);
  and _43132_ (_12188_, _12187_, _02393_);
  and _43133_ (_12189_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and _43134_ (_12190_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or _43135_ (_12191_, _12190_, _12189_);
  and _43136_ (_12193_, _12191_, _02445_);
  or _43137_ (_12194_, _12193_, _12188_);
  or _43138_ (_12195_, _12194_, _02459_);
  and _43139_ (_12196_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and _43140_ (_12197_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or _43141_ (_12198_, _12197_, _12196_);
  and _43142_ (_12199_, _12198_, _02393_);
  and _43143_ (_12200_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and _43144_ (_12201_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or _43145_ (_12202_, _12201_, _12200_);
  and _43146_ (_12203_, _12202_, _02445_);
  or _43147_ (_12204_, _12203_, _12199_);
  or _43148_ (_12205_, _12204_, _02421_);
  and _43149_ (_12206_, _12205_, _02458_);
  and _43150_ (_12207_, _12206_, _12195_);
  or _43151_ (_12208_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or _43152_ (_12209_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and _43153_ (_12210_, _12209_, _02445_);
  and _43154_ (_12211_, _12210_, _12208_);
  or _43155_ (_12212_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or _43156_ (_12213_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and _43157_ (_12214_, _12213_, _02393_);
  and _43158_ (_12215_, _12214_, _12212_);
  or _43159_ (_12216_, _12215_, _12211_);
  or _43160_ (_12217_, _12216_, _02459_);
  or _43161_ (_12218_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or _43162_ (_12219_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and _43163_ (_12220_, _12219_, _02445_);
  and _43164_ (_12221_, _12220_, _12218_);
  or _43165_ (_12222_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or _43166_ (_12225_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and _43167_ (_12227_, _12225_, _02393_);
  and _43168_ (_12229_, _12227_, _12222_);
  or _43169_ (_12231_, _12229_, _12221_);
  or _43170_ (_12233_, _12231_, _02421_);
  and _43171_ (_12235_, _12233_, _02414_);
  and _43172_ (_12236_, _12235_, _12217_);
  or _43173_ (_12238_, _12236_, _12207_);
  and _43174_ (_12240_, _12238_, _02496_);
  or _43175_ (_12242_, _12240_, _12183_);
  and _43176_ (_12244_, _12242_, _02546_);
  or _43177_ (_12246_, _12244_, _12135_);
  and _43178_ (_12248_, _12246_, _02405_);
  or _43179_ (_12250_, _12248_, _12013_);
  and _43180_ (_12251_, _12250_, _26777_);
  and _43181_ (_12253_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and _43182_ (_12255_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or _43183_ (_12257_, _12255_, _12253_);
  and _43184_ (_12259_, _12257_, _02393_);
  and _43185_ (_12261_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and _43186_ (_12262_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or _43187_ (_12263_, _12262_, _12261_);
  and _43188_ (_12265_, _12263_, _02445_);
  or _43189_ (_12267_, _12265_, _12259_);
  and _43190_ (_12269_, _12267_, _02421_);
  and _43191_ (_12270_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and _43192_ (_12271_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or _43193_ (_12272_, _12271_, _12270_);
  and _43194_ (_12274_, _12272_, _02393_);
  and _43195_ (_12275_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and _43196_ (_12276_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or _43197_ (_12278_, _12276_, _12275_);
  and _43198_ (_12279_, _12278_, _02445_);
  or _43199_ (_12281_, _12279_, _12274_);
  and _43200_ (_12283_, _12281_, _02459_);
  or _43201_ (_12285_, _12283_, _12269_);
  and _43202_ (_12286_, _12285_, _02458_);
  or _43203_ (_12287_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or _43204_ (_12289_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and _43205_ (_12291_, _12289_, _12287_);
  and _43206_ (_12293_, _12291_, _02393_);
  or _43207_ (_12295_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or _43208_ (_12296_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and _43209_ (_12297_, _12296_, _12295_);
  and _43210_ (_12298_, _12297_, _02445_);
  or _43211_ (_12299_, _12298_, _12293_);
  and _43212_ (_12300_, _12299_, _02421_);
  or _43213_ (_12301_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or _43214_ (_12302_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and _43215_ (_12303_, _12302_, _12301_);
  and _43216_ (_12304_, _12303_, _02393_);
  or _43217_ (_12305_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or _43218_ (_12306_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and _43219_ (_12307_, _12306_, _12305_);
  and _43220_ (_12308_, _12307_, _02445_);
  or _43221_ (_12309_, _12308_, _12304_);
  and _43222_ (_12310_, _12309_, _02459_);
  or _43223_ (_12311_, _12310_, _12300_);
  and _43224_ (_12312_, _12311_, _02414_);
  or _43225_ (_12313_, _12312_, _12286_);
  and _43226_ (_12314_, _12313_, _02398_);
  and _43227_ (_12315_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and _43228_ (_12316_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or _43229_ (_12317_, _12316_, _12315_);
  and _43230_ (_12318_, _12317_, _02393_);
  and _43231_ (_12319_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and _43232_ (_12320_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or _43233_ (_12321_, _12320_, _12319_);
  and _43234_ (_12322_, _12321_, _02445_);
  or _43235_ (_12323_, _12322_, _12318_);
  and _43236_ (_12324_, _12323_, _02421_);
  and _43237_ (_12325_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and _43238_ (_12326_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _43239_ (_12327_, _12326_, _12325_);
  and _43240_ (_12328_, _12327_, _02393_);
  and _43241_ (_12329_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and _43242_ (_12330_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or _43243_ (_12331_, _12330_, _12329_);
  and _43244_ (_12332_, _12331_, _02445_);
  or _43245_ (_12333_, _12332_, _12328_);
  and _43246_ (_12334_, _12333_, _02459_);
  or _43247_ (_12335_, _12334_, _12324_);
  and _43248_ (_12336_, _12335_, _02458_);
  or _43249_ (_12337_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _43250_ (_12338_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and _43251_ (_12339_, _12338_, _02445_);
  and _43252_ (_12340_, _12339_, _12337_);
  or _43253_ (_12341_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or _43254_ (_12342_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and _43255_ (_12343_, _12342_, _02393_);
  and _43256_ (_12345_, _12343_, _12341_);
  or _43257_ (_12346_, _12345_, _12340_);
  and _43258_ (_12347_, _12346_, _02421_);
  or _43259_ (_12348_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _43260_ (_12349_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and _43261_ (_12350_, _12349_, _02445_);
  and _43262_ (_12351_, _12350_, _12348_);
  or _43263_ (_12352_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or _43264_ (_12353_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and _43265_ (_12354_, _12353_, _02393_);
  and _43266_ (_12355_, _12354_, _12352_);
  or _43267_ (_12356_, _12355_, _12351_);
  and _43268_ (_12357_, _12356_, _02459_);
  or _43269_ (_12358_, _12357_, _12347_);
  and _43270_ (_12359_, _12358_, _02414_);
  or _43271_ (_12360_, _12359_, _12336_);
  and _43272_ (_12361_, _12360_, _02496_);
  or _43273_ (_12362_, _12361_, _12314_);
  and _43274_ (_12363_, _12362_, _02400_);
  and _43275_ (_12364_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and _43276_ (_12365_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or _43277_ (_12366_, _12365_, _12364_);
  and _43278_ (_12367_, _12366_, _02393_);
  and _43279_ (_12368_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  and _43280_ (_12369_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or _43281_ (_12370_, _12369_, _12368_);
  and _43282_ (_12371_, _12370_, _02445_);
  or _43283_ (_12372_, _12371_, _12367_);
  or _43284_ (_12373_, _12372_, _02459_);
  and _43285_ (_12374_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and _43286_ (_12375_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or _43287_ (_12376_, _12375_, _12374_);
  and _43288_ (_12377_, _12376_, _02393_);
  and _43289_ (_12378_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and _43290_ (_12379_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or _43291_ (_12380_, _12379_, _12378_);
  and _43292_ (_12381_, _12380_, _02445_);
  or _43293_ (_12382_, _12381_, _12377_);
  or _43294_ (_12383_, _12382_, _02421_);
  and _43295_ (_12384_, _12383_, _02458_);
  and _43296_ (_12385_, _12384_, _12373_);
  or _43297_ (_12386_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or _43298_ (_12387_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and _43299_ (_12388_, _12387_, _02445_);
  and _43300_ (_12389_, _12388_, _12386_);
  or _43301_ (_12390_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or _43302_ (_12391_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and _43303_ (_12392_, _12391_, _02393_);
  and _43304_ (_12393_, _12392_, _12390_);
  or _43305_ (_12394_, _12393_, _12389_);
  or _43306_ (_12396_, _12394_, _02459_);
  or _43307_ (_12397_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or _43308_ (_12398_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and _43309_ (_12399_, _12398_, _02445_);
  and _43310_ (_12400_, _12399_, _12397_);
  or _43311_ (_12401_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or _43312_ (_12402_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  and _43313_ (_12403_, _12402_, _02393_);
  and _43314_ (_12404_, _12403_, _12401_);
  or _43315_ (_12405_, _12404_, _12400_);
  or _43316_ (_12406_, _12405_, _02421_);
  and _43317_ (_12407_, _12406_, _02414_);
  and _43318_ (_12408_, _12407_, _12396_);
  or _43319_ (_12409_, _12408_, _12385_);
  and _43320_ (_12410_, _12409_, _02496_);
  and _43321_ (_12411_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and _43322_ (_12412_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or _43323_ (_12413_, _12412_, _12411_);
  and _43324_ (_12414_, _12413_, _02393_);
  and _43325_ (_12415_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and _43326_ (_12416_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or _43327_ (_12417_, _12416_, _12415_);
  and _43328_ (_12418_, _12417_, _02445_);
  or _43329_ (_12419_, _12418_, _12414_);
  or _43330_ (_12420_, _12419_, _02459_);
  and _43331_ (_12421_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and _43332_ (_12422_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or _43333_ (_12423_, _12422_, _12421_);
  and _43334_ (_12424_, _12423_, _02393_);
  and _43335_ (_12425_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  and _43336_ (_12426_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or _43337_ (_12427_, _12426_, _12425_);
  and _43338_ (_12428_, _12427_, _02445_);
  or _43339_ (_12429_, _12428_, _12424_);
  or _43340_ (_12430_, _12429_, _02421_);
  and _43341_ (_12431_, _12430_, _02458_);
  and _43342_ (_12432_, _12431_, _12420_);
  or _43343_ (_12433_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or _43344_ (_12434_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and _43345_ (_12435_, _12434_, _12433_);
  and _43346_ (_12436_, _12435_, _02393_);
  or _43347_ (_12437_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or _43348_ (_12438_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  and _43349_ (_12439_, _12438_, _12437_);
  and _43350_ (_12440_, _12439_, _02445_);
  or _43351_ (_12441_, _12440_, _12436_);
  or _43352_ (_12442_, _12441_, _02459_);
  or _43353_ (_12443_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or _43354_ (_12444_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and _43355_ (_12445_, _12444_, _12443_);
  and _43356_ (_12446_, _12445_, _02393_);
  or _43357_ (_12447_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or _43358_ (_12448_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and _43359_ (_12449_, _12448_, _12447_);
  and _43360_ (_12450_, _12449_, _02445_);
  or _43361_ (_12451_, _12450_, _12446_);
  or _43362_ (_12452_, _12451_, _02421_);
  and _43363_ (_12453_, _12452_, _02414_);
  and _43364_ (_12454_, _12453_, _12442_);
  or _43365_ (_12455_, _12454_, _12432_);
  and _43366_ (_12456_, _12455_, _02398_);
  or _43367_ (_12457_, _12456_, _12410_);
  and _43368_ (_12458_, _12457_, _02546_);
  or _43369_ (_12459_, _12458_, _12363_);
  and _43370_ (_12460_, _12459_, _02646_);
  or _43371_ (_12461_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or _43372_ (_12462_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and _43373_ (_12463_, _12462_, _02445_);
  and _43374_ (_12464_, _12463_, _12461_);
  or _43375_ (_12465_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or _43376_ (_12466_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and _43377_ (_12467_, _12466_, _02393_);
  and _43378_ (_12468_, _12467_, _12465_);
  or _43379_ (_12469_, _12468_, _12464_);
  and _43380_ (_12470_, _12469_, _02459_);
  or _43381_ (_12471_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or _43382_ (_12472_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and _43383_ (_12473_, _12472_, _02445_);
  and _43384_ (_12474_, _12473_, _12471_);
  or _43385_ (_12475_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or _43386_ (_12476_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  and _43387_ (_12478_, _12476_, _02393_);
  and _43388_ (_12479_, _12478_, _12475_);
  or _43389_ (_12480_, _12479_, _12474_);
  and _43390_ (_12481_, _12480_, _02421_);
  or _43391_ (_12482_, _12481_, _12470_);
  and _43392_ (_12483_, _12482_, _02414_);
  and _43393_ (_12484_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and _43394_ (_12485_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or _43395_ (_12486_, _12485_, _12484_);
  and _43396_ (_12487_, _12486_, _02393_);
  and _43397_ (_12488_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and _43398_ (_12489_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or _43399_ (_12490_, _12489_, _12488_);
  and _43400_ (_12491_, _12490_, _02445_);
  or _43401_ (_12492_, _12491_, _12487_);
  and _43402_ (_12493_, _12492_, _02459_);
  and _43403_ (_12494_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and _43404_ (_12495_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or _43405_ (_12496_, _12495_, _12494_);
  and _43406_ (_12497_, _12496_, _02393_);
  and _43407_ (_12498_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and _43408_ (_12499_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or _43409_ (_12500_, _12499_, _12498_);
  and _43410_ (_12501_, _12500_, _02445_);
  or _43411_ (_12502_, _12501_, _12497_);
  and _43412_ (_12503_, _12502_, _02421_);
  or _43413_ (_12504_, _12503_, _12493_);
  and _43414_ (_12505_, _12504_, _02458_);
  or _43415_ (_12506_, _12505_, _12483_);
  and _43416_ (_12508_, _12506_, _02496_);
  or _43417_ (_12510_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or _43418_ (_12511_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  and _43419_ (_12512_, _12511_, _12510_);
  and _43420_ (_12513_, _12512_, _02393_);
  or _43421_ (_12514_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or _43422_ (_12515_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and _43423_ (_12516_, _12515_, _12514_);
  and _43424_ (_12517_, _12516_, _02445_);
  or _43425_ (_12518_, _12517_, _12513_);
  and _43426_ (_12519_, _12518_, _02459_);
  or _43427_ (_12520_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or _43428_ (_12521_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and _43429_ (_12522_, _12521_, _12520_);
  and _43430_ (_12523_, _12522_, _02393_);
  or _43431_ (_12524_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or _43432_ (_12525_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  and _43433_ (_12526_, _12525_, _12524_);
  and _43434_ (_12527_, _12526_, _02445_);
  or _43435_ (_12528_, _12527_, _12523_);
  and _43436_ (_12530_, _12528_, _02421_);
  or _43437_ (_12531_, _12530_, _12519_);
  and _43438_ (_12532_, _12531_, _02414_);
  and _43439_ (_12533_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and _43440_ (_12534_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or _43441_ (_12535_, _12534_, _12533_);
  and _43442_ (_12536_, _12535_, _02393_);
  and _43443_ (_12537_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and _43444_ (_12538_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or _43445_ (_12539_, _12538_, _12537_);
  and _43446_ (_12541_, _12539_, _02445_);
  or _43447_ (_12542_, _12541_, _12536_);
  and _43448_ (_12544_, _12542_, _02459_);
  and _43449_ (_12546_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and _43450_ (_12547_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or _43451_ (_12548_, _12547_, _12546_);
  and _43452_ (_12549_, _12548_, _02393_);
  and _43453_ (_12550_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and _43454_ (_12551_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or _43455_ (_12552_, _12551_, _12550_);
  and _43456_ (_12553_, _12552_, _02445_);
  or _43457_ (_12554_, _12553_, _12549_);
  and _43458_ (_12555_, _12554_, _02421_);
  or _43459_ (_12556_, _12555_, _12544_);
  and _43460_ (_12557_, _12556_, _02458_);
  or _43461_ (_12558_, _12557_, _12532_);
  and _43462_ (_12559_, _12558_, _02398_);
  or _43463_ (_12560_, _12559_, _12508_);
  and _43464_ (_12561_, _12560_, _02400_);
  and _43465_ (_12562_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and _43466_ (_12563_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or _43467_ (_12564_, _12563_, _12562_);
  and _43468_ (_12566_, _12564_, _02393_);
  and _43469_ (_12567_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and _43470_ (_12568_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or _43471_ (_12570_, _12568_, _12567_);
  and _43472_ (_12571_, _12570_, _02445_);
  or _43473_ (_12572_, _12571_, _12566_);
  or _43474_ (_12573_, _12572_, _02459_);
  and _43475_ (_12574_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and _43476_ (_12575_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or _43477_ (_12576_, _12575_, _12574_);
  and _43478_ (_12577_, _12576_, _02393_);
  and _43479_ (_12578_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and _43480_ (_12579_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or _43481_ (_12580_, _12579_, _12578_);
  and _43482_ (_12581_, _12580_, _02445_);
  or _43483_ (_12582_, _12581_, _12577_);
  or _43484_ (_12583_, _12582_, _02421_);
  and _43485_ (_12584_, _12583_, _02458_);
  and _43486_ (_12585_, _12584_, _12573_);
  or _43487_ (_12587_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or _43488_ (_12588_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and _43489_ (_12589_, _12588_, _12587_);
  and _43490_ (_12590_, _12589_, _02393_);
  or _43491_ (_12591_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or _43492_ (_12592_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and _43493_ (_12593_, _12592_, _12591_);
  and _43494_ (_12594_, _12593_, _02445_);
  or _43495_ (_12595_, _12594_, _12590_);
  or _43496_ (_12596_, _12595_, _02459_);
  or _43497_ (_12597_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or _43498_ (_12598_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and _43499_ (_12599_, _12598_, _12597_);
  and _43500_ (_12600_, _12599_, _02393_);
  or _43501_ (_12601_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or _43502_ (_12602_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and _43503_ (_12603_, _12602_, _12601_);
  and _43504_ (_12604_, _12603_, _02445_);
  or _43505_ (_12605_, _12604_, _12600_);
  or _43506_ (_12606_, _12605_, _02421_);
  and _43507_ (_12607_, _12606_, _02414_);
  and _43508_ (_12608_, _12607_, _12596_);
  or _43509_ (_12609_, _12608_, _12585_);
  and _43510_ (_12610_, _12609_, _02398_);
  and _43511_ (_12611_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  and _43512_ (_12612_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or _43513_ (_12614_, _12612_, _12611_);
  and _43514_ (_12616_, _12614_, _02393_);
  and _43515_ (_12618_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and _43516_ (_12619_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or _43517_ (_12620_, _12619_, _12618_);
  and _43518_ (_12621_, _12620_, _02445_);
  or _43519_ (_12622_, _12621_, _12616_);
  or _43520_ (_12623_, _12622_, _02459_);
  and _43521_ (_12624_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and _43522_ (_12625_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or _43523_ (_12626_, _12625_, _12624_);
  and _43524_ (_12627_, _12626_, _02393_);
  and _43525_ (_12628_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and _43526_ (_12629_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or _43527_ (_12630_, _12629_, _12628_);
  and _43528_ (_12631_, _12630_, _02445_);
  or _43529_ (_12633_, _12631_, _12627_);
  or _43530_ (_12634_, _12633_, _02421_);
  and _43531_ (_12635_, _12634_, _02458_);
  and _43532_ (_12636_, _12635_, _12623_);
  or _43533_ (_12637_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or _43534_ (_12638_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and _43535_ (_12639_, _12638_, _02445_);
  and _43536_ (_12640_, _12639_, _12637_);
  or _43537_ (_12641_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or _43538_ (_12642_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and _43539_ (_12643_, _12642_, _02393_);
  and _43540_ (_12644_, _12643_, _12641_);
  or _43541_ (_12645_, _12644_, _12640_);
  or _43542_ (_12646_, _12645_, _02459_);
  or _43543_ (_12647_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or _43544_ (_12648_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and _43545_ (_12649_, _12648_, _02445_);
  and _43546_ (_12650_, _12649_, _12647_);
  or _43547_ (_12651_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or _43548_ (_12652_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  and _43549_ (_12653_, _12652_, _02393_);
  and _43550_ (_12654_, _12653_, _12651_);
  or _43551_ (_12655_, _12654_, _12650_);
  or _43552_ (_12656_, _12655_, _02421_);
  and _43553_ (_12657_, _12656_, _02414_);
  and _43554_ (_12658_, _12657_, _12646_);
  or _43555_ (_12659_, _12658_, _12636_);
  and _43556_ (_12660_, _12659_, _02496_);
  or _43557_ (_12661_, _12660_, _12610_);
  and _43558_ (_12662_, _12661_, _02546_);
  or _43559_ (_12663_, _12662_, _12561_);
  and _43560_ (_12664_, _12663_, _02405_);
  or _43561_ (_12665_, _12664_, _12460_);
  and _43562_ (_12666_, _12665_, _02444_);
  or _43563_ (_12667_, _12666_, _12251_);
  or _43564_ (_12668_, _12667_, _02443_);
  or _43565_ (_12669_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and _43566_ (_12670_, _12669_, _22762_);
  and _43567_ (_03400_, _12670_, _12668_);
  not _43568_ (_12671_, _02077_);
  or _43569_ (_12673_, _12671_, _23892_);
  not _43570_ (_12675_, _02073_);
  and _43571_ (_12676_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _43572_ (_12677_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _43573_ (_12678_, _12677_, _12676_);
  or _43574_ (_12680_, _12678_, _02077_);
  and _43575_ (_12682_, _12680_, _12675_);
  and _43576_ (_12683_, _12682_, _12673_);
  and _43577_ (_12684_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _43578_ (_12685_, _12684_, _12683_);
  and _43579_ (_03406_, _12685_, _22762_);
  or _43580_ (_12686_, _12675_, _23642_);
  not _43581_ (_12687_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor _43582_ (_12688_, _02078_, _12687_);
  and _43583_ (_12689_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _43584_ (_12690_, _12689_, _12688_);
  or _43585_ (_12691_, _12690_, _02073_);
  and _43586_ (_12692_, _12691_, _22762_);
  and _43587_ (_03409_, _12692_, _12686_);
  and _43588_ (_12693_, _02284_, _23824_);
  and _43589_ (_12694_, _02286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  or _43590_ (_27117_, _12694_, _12693_);
  and _43591_ (_12695_, _03339_, _24050_);
  and _43592_ (_12696_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or _43593_ (_03418_, _12696_, _12695_);
  and _43594_ (_12697_, _02374_, _23747_);
  and _43595_ (_12698_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  or _43596_ (_03433_, _12698_, _12697_);
  and _43597_ (_12699_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  and _43598_ (_12700_, _06888_, _23778_);
  or _43599_ (_03436_, _12700_, _12699_);
  and _43600_ (_12701_, _05180_, _23707_);
  and _43601_ (_12702_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or _43602_ (_03439_, _12702_, _12701_);
  and _43603_ (_12703_, _04797_, _23898_);
  and _43604_ (_12705_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or _43605_ (_03441_, _12705_, _12703_);
  or _43606_ (_12707_, _02009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _43607_ (_12708_, _02009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _43608_ (_12709_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _43609_ (_12710_, _12709_, _01996_);
  nand _43610_ (_12712_, _12710_, _12708_);
  and _43611_ (_12713_, _12712_, _12707_);
  or _43612_ (_12714_, _12713_, _02001_);
  or _43613_ (_12715_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _43614_ (_12716_, _12715_, _01979_);
  and _43615_ (_12718_, _12716_, _12714_);
  and _43616_ (_12719_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _43617_ (_12721_, _01977_, _24685_);
  or _43618_ (_12722_, _12721_, _12719_);
  or _43619_ (_12723_, _12722_, _12718_);
  and _43620_ (_03444_, _12723_, _22762_);
  and _43621_ (_12724_, _08360_, _24050_);
  and _43622_ (_12725_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  or _43623_ (_03448_, _12725_, _12724_);
  and _43624_ (_12726_, _08198_, _23946_);
  and _43625_ (_12727_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or _43626_ (_03453_, _12727_, _12726_);
  and _43627_ (_12728_, _06886_, _23986_);
  not _43628_ (_12729_, _12728_);
  and _43629_ (_12730_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  and _43630_ (_12732_, _12728_, _23707_);
  or _43631_ (_03463_, _12732_, _12730_);
  and _43632_ (_12733_, _23986_, _23664_);
  and _43633_ (_12734_, _12733_, _23649_);
  not _43634_ (_12735_, _12733_);
  and _43635_ (_12737_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  or _43636_ (_27085_, _12737_, _12734_);
  and _43637_ (_12738_, _01977_, _23642_);
  and _43638_ (_12739_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _43639_ (_12740_, _12739_, _02041_);
  nand _43640_ (_12742_, _02009_, _01983_);
  nor _43641_ (_12743_, _12742_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _43642_ (_12744_, _12742_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _43643_ (_12745_, _12744_, _02001_);
  or _43644_ (_12746_, _12745_, _12743_);
  or _43645_ (_12747_, _12746_, _12740_);
  or _43646_ (_12748_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _43647_ (_12749_, _12748_, _01979_);
  and _43648_ (_12750_, _12749_, _12747_);
  and _43649_ (_12751_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _43650_ (_12752_, _12751_, _12750_);
  or _43651_ (_12753_, _12752_, _12738_);
  and _43652_ (_03477_, _12753_, _22762_);
  not _43653_ (_12754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _43654_ (_12755_, _02025_, _12754_);
  nand _43655_ (_12756_, _12755_, _02041_);
  not _43656_ (_12757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand _43657_ (_12758_, _02009_, _01989_);
  and _43658_ (_12759_, _12758_, _12757_);
  nor _43659_ (_12760_, _12758_, _12757_);
  or _43660_ (_12761_, _12760_, _12759_);
  and _43661_ (_12762_, _12761_, _02002_);
  nand _43662_ (_12763_, _12762_, _12756_);
  not _43663_ (_12764_, _01979_);
  and _43664_ (_12765_, _02001_, _12754_);
  nor _43665_ (_12766_, _12765_, _12764_);
  and _43666_ (_12767_, _12766_, _12763_);
  and _43667_ (_12768_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _43668_ (_12769_, _12768_, _12767_);
  and _43669_ (_12770_, _01978_, _23816_);
  or _43670_ (_12771_, _12770_, _12769_);
  and _43671_ (_03486_, _12771_, _22762_);
  and _43672_ (_12772_, _08307_, _24291_);
  nand _43673_ (_12773_, _12772_, _23594_);
  not _43674_ (_12774_, _08313_);
  or _43675_ (_12775_, _12772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _43676_ (_12776_, _12775_, _12774_);
  and _43677_ (_12777_, _12776_, _12773_);
  and _43678_ (_12778_, _08313_, _23816_);
  or _43679_ (_12779_, _12778_, _12777_);
  and _43680_ (_03500_, _12779_, _22762_);
  and _43681_ (_12780_, _08799_, _23778_);
  and _43682_ (_12781_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  or _43683_ (_03505_, _12781_, _12780_);
  and _43684_ (_12782_, _24282_, _23664_);
  and _43685_ (_12783_, _12782_, _23824_);
  not _43686_ (_12784_, _12782_);
  and _43687_ (_12785_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or _43688_ (_03509_, _12785_, _12783_);
  and _43689_ (_12786_, _24010_, _23664_);
  and _43690_ (_12787_, _12786_, _23707_);
  not _43691_ (_12788_, _12786_);
  and _43692_ (_12789_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  or _43693_ (_03518_, _12789_, _12787_);
  and _43694_ (_12790_, _08360_, _23946_);
  and _43695_ (_12791_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or _43696_ (_03524_, _12791_, _12790_);
  and _43697_ (_12792_, _05350_, _23898_);
  and _43698_ (_12793_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  or _43699_ (_03539_, _12793_, _12792_);
  and _43700_ (_12794_, _09913_, _23898_);
  and _43701_ (_12795_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or _43702_ (_03557_, _12795_, _12794_);
  and _43703_ (_12796_, _25739_, _23747_);
  and _43704_ (_12797_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  or _43705_ (_03574_, _12797_, _12796_);
  and _43706_ (_12798_, _02370_, _23946_);
  and _43707_ (_12799_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or _43708_ (_03577_, _12799_, _12798_);
  and _43709_ (_12800_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  and _43710_ (_12801_, _06888_, _23824_);
  or _43711_ (_27013_, _12801_, _12800_);
  and _43712_ (_12802_, _04811_, _23778_);
  and _43713_ (_12803_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  or _43714_ (_27066_, _12803_, _12802_);
  and _43715_ (_12804_, _03300_, _23778_);
  and _43716_ (_12806_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or _43717_ (_03605_, _12806_, _12804_);
  and _43718_ (_12807_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  and _43719_ (_12808_, _06888_, _23898_);
  or _43720_ (_03608_, _12808_, _12807_);
  and _43721_ (_12809_, _23755_, _23707_);
  and _43722_ (_12810_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or _43723_ (_03613_, _12810_, _12809_);
  and _43724_ (_12811_, _26110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor _43725_ (_12812_, _12811_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _43726_ (_12813_, _12812_, _09917_);
  and _43727_ (_12814_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _43728_ (_12815_, _12814_, _26118_);
  nor _43729_ (_12816_, _12815_, _12813_);
  nor _43730_ (_12817_, _12816_, _24299_);
  and _43731_ (_12818_, _24299_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _43732_ (_12819_, _12818_, _12817_);
  and _43733_ (_12820_, _12819_, _24294_);
  and _43734_ (_12821_, _24293_, _23892_);
  or _43735_ (_12822_, _12821_, _12820_);
  and _43736_ (_03628_, _12822_, _22762_);
  and _43737_ (_12823_, _24226_, _23946_);
  and _43738_ (_12824_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or _43739_ (_03638_, _12824_, _12823_);
  and _43740_ (_12825_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  and _43741_ (_12826_, _25252_, _23778_);
  or _43742_ (_03656_, _12826_, _12825_);
  and _43743_ (_12827_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  and _43744_ (_12828_, _25542_, _23747_);
  or _43745_ (_03664_, _12828_, _12827_);
  and _43746_ (_12829_, _24201_, _24085_);
  not _43747_ (_12830_, _12829_);
  and _43748_ (_12831_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and _43749_ (_12832_, _12829_, _24050_);
  or _43750_ (_03676_, _12832_, _12831_);
  and _43751_ (_12833_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  and _43752_ (_12834_, _02245_, _23898_);
  or _43753_ (_27035_, _12834_, _12833_);
  and _43754_ (_12835_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  and _43755_ (_12836_, _12728_, _23824_);
  or _43756_ (_03680_, _12836_, _12835_);
  and _43757_ (_12837_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  and _43758_ (_12838_, _12728_, _23898_);
  or _43759_ (_03683_, _12838_, _12837_);
  and _43760_ (_12839_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  and _43761_ (_12840_, _04748_, _24050_);
  or _43762_ (_27032_, _12840_, _12839_);
  and _43763_ (_12841_, _05008_, _23649_);
  and _43764_ (_12842_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or _43765_ (_03701_, _12842_, _12841_);
  and _43766_ (_12843_, _05008_, _23898_);
  and _43767_ (_12844_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or _43768_ (_03703_, _12844_, _12843_);
  and _43769_ (_12845_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  and _43770_ (_12846_, _12728_, _23778_);
  or _43771_ (_03710_, _12846_, _12845_);
  and _43772_ (_12847_, _05288_, _23946_);
  and _43773_ (_12848_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  or _43774_ (_03713_, _12848_, _12847_);
  and _43775_ (_12849_, _05701_, _23747_);
  and _43776_ (_12850_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or _43777_ (_03724_, _12850_, _12849_);
  and _43778_ (_12851_, _01971_, _23649_);
  and _43779_ (_12852_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  or _43780_ (_03742_, _12852_, _12851_);
  and _43781_ (_12853_, _24050_, _23665_);
  and _43782_ (_12854_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  or _43783_ (_03748_, _12854_, _12853_);
  and _43784_ (_12855_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and _43785_ (_12856_, _06918_, _23649_);
  or _43786_ (_03751_, _12856_, _12855_);
  or _43787_ (_12857_, _04945_, _24591_);
  and _43788_ (_12858_, _24604_, _26582_);
  and _43789_ (_12859_, _26625_, _24599_);
  or _43790_ (_12860_, _12859_, _12858_);
  or _43791_ (_12861_, _12860_, _12857_);
  and _43792_ (_12862_, _25638_, _26582_);
  and _43793_ (_12863_, _24604_, _24445_);
  or _43794_ (_12864_, _12863_, _12862_);
  or _43795_ (_12865_, _04958_, _04982_);
  or _43796_ (_12866_, _12865_, _12864_);
  or _43797_ (_12867_, _12866_, _12861_);
  and _43798_ (_12868_, _24556_, _24541_);
  or _43799_ (_12869_, _05016_, _12868_);
  or _43800_ (_12870_, _12869_, _12867_);
  or _43801_ (_12871_, _04974_, _04970_);
  or _43802_ (_12872_, _12871_, _04943_);
  or _43803_ (_12873_, _24605_, _24586_);
  or _43804_ (_12874_, _12873_, _24600_);
  or _43805_ (_12875_, _02269_, _24537_);
  or _43806_ (_12876_, _12875_, _12874_);
  or _43807_ (_12877_, _12876_, _12872_);
  or _43808_ (_12878_, _12877_, _12870_);
  and _43809_ (_12879_, _12878_, _22768_);
  and _43810_ (_12880_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _43811_ (_12881_, _12880_, _05003_);
  or _43812_ (_12882_, _12881_, _12879_);
  and _43813_ (_26866_[0], _12882_, _22762_);
  and _43814_ (_12883_, _25748_, _24050_);
  and _43815_ (_12884_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or _43816_ (_03763_, _12884_, _12883_);
  and _43817_ (_12885_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  and _43818_ (_12886_, _12728_, _23946_);
  or _43819_ (_03765_, _12886_, _12885_);
  and _43820_ (_12887_, _05281_, _23946_);
  and _43821_ (_12888_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or _43822_ (_03768_, _12888_, _12887_);
  and _43823_ (_12889_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  and _43824_ (_12890_, _12728_, _23649_);
  or _43825_ (_03775_, _12890_, _12889_);
  and _43826_ (_12891_, _24331_, _23649_);
  and _43827_ (_12892_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or _43828_ (_03792_, _12892_, _12891_);
  and _43829_ (_12893_, _24081_, _23707_);
  and _43830_ (_12894_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or _43831_ (_03802_, _12894_, _12893_);
  and _43832_ (_12895_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  and _43833_ (_12896_, _25252_, _23946_);
  or _43834_ (_03809_, _12896_, _12895_);
  and _43835_ (_12897_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and _43836_ (_12898_, _25763_, _23649_);
  or _43837_ (_27041_, _12898_, _12897_);
  not _43838_ (_12899_, _25644_);
  and _43839_ (_12900_, _24598_, _24567_);
  nor _43840_ (_12901_, _12900_, _04981_);
  or _43841_ (_26862_[1], _12901_, _12899_);
  and _43842_ (_12902_, _12786_, _23778_);
  and _43843_ (_12903_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or _43844_ (_03846_, _12903_, _12902_);
  and _43845_ (_12904_, _09913_, _23824_);
  and _43846_ (_12905_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or _43847_ (_03849_, _12905_, _12904_);
  and _43848_ (_12906_, _06886_, _23069_);
  not _43849_ (_12907_, _12906_);
  and _43850_ (_12908_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and _43851_ (_12909_, _12906_, _23649_);
  or _43852_ (_03865_, _12909_, _12908_);
  and _43853_ (_12910_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  and _43854_ (_12911_, _25542_, _23649_);
  or _43855_ (_03871_, _12911_, _12910_);
  or _43856_ (_12912_, _04663_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _43857_ (_12913_, _04682_, _04666_);
  or _43858_ (_12914_, _12913_, _12912_);
  and _43859_ (_12915_, _12914_, _04694_);
  nor _43860_ (_12916_, _04693_, _24564_);
  or _43861_ (_12917_, _12916_, rst);
  or _43862_ (_26863_[0], _12917_, _12915_);
  and _43863_ (_12918_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and _43864_ (_12919_, _12906_, _23747_);
  or _43865_ (_03878_, _12919_, _12918_);
  and _43866_ (_12921_, _23833_, _23778_);
  and _43867_ (_12922_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or _43868_ (_03880_, _12922_, _12921_);
  and _43869_ (_12923_, _05125_, _23824_);
  and _43870_ (_12924_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  or _43871_ (_03883_, _12924_, _12923_);
  and _43872_ (_12925_, _08799_, _23707_);
  and _43873_ (_12926_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  or _43874_ (_03894_, _12926_, _12925_);
  and _43875_ (_12927_, _05336_, _23991_);
  not _43876_ (_12928_, _12927_);
  and _43877_ (_12929_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and _43878_ (_12930_, _12927_, _23747_);
  or _43879_ (_03936_, _12930_, _12929_);
  and _43880_ (_12931_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and _43881_ (_12932_, _12927_, _23778_);
  or _43882_ (_27103_, _12932_, _12931_);
  and _43883_ (_12933_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and _43884_ (_12934_, _12829_, _23946_);
  or _43885_ (_03969_, _12934_, _12933_);
  and _43886_ (_12935_, _05336_, _23903_);
  not _43887_ (_12936_, _12935_);
  and _43888_ (_12937_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and _43889_ (_12938_, _12935_, _23649_);
  or _43890_ (_27102_, _12938_, _12937_);
  and _43891_ (_12939_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and _43892_ (_12940_, _12906_, _23707_);
  or _43893_ (_03980_, _12940_, _12939_);
  and _43894_ (_12941_, _05336_, _24005_);
  not _43895_ (_12942_, _12941_);
  and _43896_ (_12943_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  and _43897_ (_12944_, _12941_, _24050_);
  or _43898_ (_03984_, _12944_, _12943_);
  and _43899_ (_12945_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  and _43900_ (_12946_, _12941_, _23649_);
  or _43901_ (_03987_, _12946_, _12945_);
  and _43902_ (_12947_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and _43903_ (_12948_, _12829_, _23649_);
  or _43904_ (_03995_, _12948_, _12947_);
  or _43905_ (_12949_, _24171_, _24043_);
  and _43906_ (_12951_, _24151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _43907_ (_12952_, _12951_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _43908_ (_12953_, _12951_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _43909_ (_12954_, _12953_, _12952_);
  nor _43910_ (_12955_, _24184_, _24132_);
  nor _43911_ (_12956_, _12955_, _24127_);
  and _43912_ (_12957_, _12956_, _12954_);
  not _43913_ (_12958_, _12956_);
  and _43914_ (_12959_, _12958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand _43915_ (_12960_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _43916_ (_12961_, _12960_, _24127_);
  or _43917_ (_12962_, _12961_, _12959_);
  or _43918_ (_12963_, _12962_, _12957_);
  or _43919_ (_12964_, _12963_, _24120_);
  and _43920_ (_12965_, _12964_, _22762_);
  and _43921_ (_03997_, _12965_, _12949_);
  and _43922_ (_12966_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and _43923_ (_12967_, _12906_, _24050_);
  or _43924_ (_04003_, _12967_, _12966_);
  and _43925_ (_12968_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and _43926_ (_12969_, _12906_, _23946_);
  or _43927_ (_04007_, _12969_, _12968_);
  and _43928_ (_12970_, _05336_, _23986_);
  not _43929_ (_12971_, _12970_);
  and _43930_ (_12972_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  and _43931_ (_12973_, _12970_, _23898_);
  or _43932_ (_27098_, _12973_, _12972_);
  and _43933_ (_12974_, _05336_, _23069_);
  not _43934_ (_12975_, _12974_);
  and _43935_ (_12976_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and _43936_ (_12977_, _12974_, _23649_);
  or _43937_ (_27096_, _12977_, _12976_);
  and _43938_ (_12978_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and _43939_ (_12979_, _06918_, _23898_);
  or _43940_ (_04025_, _12979_, _12978_);
  and _43941_ (_12980_, _05336_, _01808_);
  not _43942_ (_12981_, _12980_);
  and _43943_ (_12982_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and _43944_ (_12983_, _12980_, _23649_);
  or _43945_ (_04031_, _12983_, _12982_);
  and _43946_ (_12984_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and _43947_ (_12985_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or _43948_ (_12986_, _12985_, _12984_);
  and _43949_ (_12987_, _12986_, _02393_);
  and _43950_ (_12988_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and _43951_ (_12989_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or _43952_ (_12990_, _12989_, _12988_);
  and _43953_ (_12991_, _12990_, _02445_);
  or _43954_ (_12992_, _12991_, _12987_);
  and _43955_ (_12993_, _12992_, _02421_);
  and _43956_ (_12994_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and _43957_ (_12995_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or _43958_ (_12996_, _12995_, _12994_);
  and _43959_ (_12997_, _12996_, _02393_);
  and _43960_ (_12998_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and _43961_ (_12999_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or _43962_ (_13000_, _12999_, _12998_);
  and _43963_ (_13001_, _13000_, _02445_);
  or _43964_ (_13002_, _13001_, _12997_);
  and _43965_ (_13003_, _13002_, _02459_);
  or _43966_ (_13004_, _13003_, _12993_);
  and _43967_ (_13005_, _13004_, _02458_);
  or _43968_ (_13006_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or _43969_ (_13007_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and _43970_ (_13008_, _13007_, _13006_);
  and _43971_ (_13009_, _13008_, _02393_);
  or _43972_ (_13010_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or _43973_ (_13011_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and _43974_ (_13012_, _13011_, _13010_);
  and _43975_ (_13013_, _13012_, _02445_);
  or _43976_ (_13014_, _13013_, _13009_);
  and _43977_ (_13015_, _13014_, _02421_);
  or _43978_ (_13016_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or _43979_ (_13017_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and _43980_ (_13018_, _13017_, _13016_);
  and _43981_ (_13019_, _13018_, _02393_);
  or _43982_ (_13020_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or _43983_ (_13021_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and _43984_ (_13022_, _13021_, _13020_);
  and _43985_ (_13023_, _13022_, _02445_);
  or _43986_ (_13024_, _13023_, _13019_);
  and _43987_ (_13025_, _13024_, _02459_);
  or _43988_ (_13026_, _13025_, _13015_);
  and _43989_ (_13027_, _13026_, _02414_);
  or _43990_ (_13028_, _13027_, _13005_);
  and _43991_ (_13029_, _13028_, _02398_);
  and _43992_ (_13030_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and _43993_ (_13031_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or _43994_ (_13032_, _13031_, _13030_);
  and _43995_ (_13033_, _13032_, _02393_);
  and _43996_ (_13034_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and _43997_ (_13035_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or _43998_ (_13036_, _13035_, _13034_);
  and _43999_ (_13037_, _13036_, _02445_);
  or _44000_ (_13038_, _13037_, _13033_);
  and _44001_ (_13039_, _13038_, _02421_);
  and _44002_ (_13040_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and _44003_ (_13041_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or _44004_ (_13042_, _13041_, _13040_);
  and _44005_ (_13043_, _13042_, _02393_);
  and _44006_ (_13044_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and _44007_ (_13045_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or _44008_ (_13046_, _13045_, _13044_);
  and _44009_ (_13047_, _13046_, _02445_);
  or _44010_ (_13048_, _13047_, _13043_);
  and _44011_ (_13049_, _13048_, _02459_);
  or _44012_ (_13050_, _13049_, _13039_);
  and _44013_ (_13051_, _13050_, _02458_);
  or _44014_ (_13052_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or _44015_ (_13053_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and _44016_ (_13054_, _13053_, _02445_);
  and _44017_ (_13055_, _13054_, _13052_);
  or _44018_ (_13056_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or _44019_ (_13057_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and _44020_ (_13058_, _13057_, _02393_);
  and _44021_ (_13059_, _13058_, _13056_);
  or _44022_ (_13060_, _13059_, _13055_);
  and _44023_ (_13061_, _13060_, _02421_);
  or _44024_ (_13062_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or _44025_ (_13063_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and _44026_ (_13064_, _13063_, _02445_);
  and _44027_ (_13065_, _13064_, _13062_);
  or _44028_ (_13066_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or _44029_ (_13067_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and _44030_ (_13068_, _13067_, _02393_);
  and _44031_ (_13069_, _13068_, _13066_);
  or _44032_ (_13070_, _13069_, _13065_);
  and _44033_ (_13071_, _13070_, _02459_);
  or _44034_ (_13072_, _13071_, _13061_);
  and _44035_ (_13073_, _13072_, _02414_);
  or _44036_ (_13074_, _13073_, _13051_);
  and _44037_ (_13075_, _13074_, _02496_);
  or _44038_ (_13076_, _13075_, _13029_);
  and _44039_ (_13077_, _13076_, _02400_);
  and _44040_ (_13078_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and _44041_ (_13079_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or _44042_ (_13080_, _13079_, _13078_);
  and _44043_ (_13081_, _13080_, _02393_);
  and _44044_ (_13082_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and _44045_ (_13083_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or _44046_ (_13084_, _13083_, _13082_);
  and _44047_ (_13085_, _13084_, _02445_);
  or _44048_ (_13086_, _13085_, _13081_);
  or _44049_ (_13087_, _13086_, _02459_);
  and _44050_ (_13088_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and _44051_ (_13089_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or _44052_ (_13090_, _13089_, _13088_);
  and _44053_ (_13091_, _13090_, _02393_);
  and _44054_ (_13092_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and _44055_ (_13093_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or _44056_ (_13094_, _13093_, _13092_);
  and _44057_ (_13095_, _13094_, _02445_);
  or _44058_ (_13096_, _13095_, _13091_);
  or _44059_ (_13097_, _13096_, _02421_);
  and _44060_ (_13098_, _13097_, _02458_);
  and _44061_ (_13099_, _13098_, _13087_);
  or _44062_ (_13100_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or _44063_ (_13101_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and _44064_ (_13102_, _13101_, _02445_);
  and _44065_ (_13103_, _13102_, _13100_);
  or _44066_ (_13104_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or _44067_ (_13105_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and _44068_ (_13106_, _13105_, _02393_);
  and _44069_ (_13107_, _13106_, _13104_);
  or _44070_ (_13108_, _13107_, _13103_);
  or _44071_ (_13109_, _13108_, _02459_);
  or _44072_ (_13110_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or _44073_ (_13111_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and _44074_ (_13112_, _13111_, _02445_);
  and _44075_ (_13113_, _13112_, _13110_);
  or _44076_ (_13114_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or _44077_ (_13115_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and _44078_ (_13116_, _13115_, _02393_);
  and _44079_ (_13117_, _13116_, _13114_);
  or _44080_ (_13118_, _13117_, _13113_);
  or _44081_ (_13119_, _13118_, _02421_);
  and _44082_ (_13120_, _13119_, _02414_);
  and _44083_ (_13121_, _13120_, _13109_);
  or _44084_ (_13122_, _13121_, _13099_);
  and _44085_ (_13123_, _13122_, _02496_);
  and _44086_ (_13124_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and _44087_ (_13125_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or _44088_ (_13126_, _13125_, _13124_);
  and _44089_ (_13127_, _13126_, _02393_);
  and _44090_ (_13128_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and _44091_ (_13129_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or _44092_ (_13130_, _13129_, _13128_);
  and _44093_ (_13131_, _13130_, _02445_);
  or _44094_ (_13132_, _13131_, _13127_);
  or _44095_ (_13133_, _13132_, _02459_);
  and _44096_ (_13134_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and _44097_ (_13135_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or _44098_ (_13136_, _13135_, _13134_);
  and _44099_ (_13137_, _13136_, _02393_);
  and _44100_ (_13138_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and _44101_ (_13139_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or _44102_ (_13140_, _13139_, _13138_);
  and _44103_ (_13141_, _13140_, _02445_);
  or _44104_ (_13142_, _13141_, _13137_);
  or _44105_ (_13143_, _13142_, _02421_);
  and _44106_ (_13144_, _13143_, _02458_);
  and _44107_ (_13145_, _13144_, _13133_);
  or _44108_ (_13146_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or _44109_ (_13147_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and _44110_ (_13148_, _13147_, _13146_);
  and _44111_ (_13149_, _13148_, _02393_);
  or _44112_ (_13150_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or _44113_ (_13151_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and _44114_ (_13152_, _13151_, _13150_);
  and _44115_ (_13153_, _13152_, _02445_);
  or _44116_ (_13154_, _13153_, _13149_);
  or _44117_ (_13155_, _13154_, _02459_);
  or _44118_ (_13156_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or _44119_ (_13157_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and _44120_ (_13158_, _13157_, _13156_);
  and _44121_ (_13159_, _13158_, _02393_);
  or _44122_ (_13160_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or _44123_ (_13161_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and _44124_ (_13162_, _13161_, _13160_);
  and _44125_ (_13163_, _13162_, _02445_);
  or _44126_ (_13164_, _13163_, _13159_);
  or _44127_ (_13165_, _13164_, _02421_);
  and _44128_ (_13166_, _13165_, _02414_);
  and _44129_ (_13167_, _13166_, _13155_);
  or _44130_ (_13168_, _13167_, _13145_);
  and _44131_ (_13169_, _13168_, _02398_);
  or _44132_ (_13170_, _13169_, _13123_);
  and _44133_ (_13171_, _13170_, _02546_);
  or _44134_ (_13172_, _13171_, _13077_);
  and _44135_ (_13173_, _13172_, _02646_);
  or _44136_ (_13174_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or _44137_ (_13175_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and _44138_ (_13176_, _13175_, _02445_);
  and _44139_ (_13177_, _13176_, _13174_);
  or _44140_ (_13178_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or _44141_ (_13179_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and _44142_ (_13180_, _13179_, _02393_);
  and _44143_ (_13181_, _13180_, _13178_);
  or _44144_ (_13182_, _13181_, _13177_);
  and _44145_ (_13183_, _13182_, _02459_);
  or _44146_ (_13184_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or _44147_ (_13185_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and _44148_ (_13186_, _13185_, _02445_);
  and _44149_ (_13187_, _13186_, _13184_);
  or _44150_ (_13188_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or _44151_ (_13189_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and _44152_ (_13190_, _13189_, _02393_);
  and _44153_ (_13191_, _13190_, _13188_);
  or _44154_ (_13192_, _13191_, _13187_);
  and _44155_ (_13193_, _13192_, _02421_);
  or _44156_ (_13194_, _13193_, _13183_);
  and _44157_ (_13195_, _13194_, _02414_);
  and _44158_ (_13196_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and _44159_ (_13197_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or _44160_ (_13198_, _13197_, _13196_);
  and _44161_ (_13199_, _13198_, _02393_);
  and _44162_ (_13200_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and _44163_ (_13201_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or _44164_ (_13202_, _13201_, _13200_);
  and _44165_ (_13203_, _13202_, _02445_);
  or _44166_ (_13204_, _13203_, _13199_);
  and _44167_ (_13205_, _13204_, _02459_);
  and _44168_ (_13206_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  and _44169_ (_13207_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or _44170_ (_13208_, _13207_, _13206_);
  and _44171_ (_13209_, _13208_, _02393_);
  and _44172_ (_13210_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and _44173_ (_13211_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or _44174_ (_13212_, _13211_, _13210_);
  and _44175_ (_13213_, _13212_, _02445_);
  or _44176_ (_13214_, _13213_, _13209_);
  and _44177_ (_13215_, _13214_, _02421_);
  or _44178_ (_13216_, _13215_, _13205_);
  and _44179_ (_13217_, _13216_, _02458_);
  or _44180_ (_13218_, _13217_, _13195_);
  and _44181_ (_13219_, _13218_, _02496_);
  or _44182_ (_13220_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or _44183_ (_13221_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and _44184_ (_13222_, _13221_, _13220_);
  and _44185_ (_13223_, _13222_, _02393_);
  or _44186_ (_13224_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or _44187_ (_13225_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and _44188_ (_13226_, _13225_, _13224_);
  and _44189_ (_13227_, _13226_, _02445_);
  or _44190_ (_13228_, _13227_, _13223_);
  and _44191_ (_13229_, _13228_, _02459_);
  or _44192_ (_13230_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or _44193_ (_13231_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and _44194_ (_13232_, _13231_, _13230_);
  and _44195_ (_13233_, _13232_, _02393_);
  or _44196_ (_13234_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or _44197_ (_13235_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and _44198_ (_13236_, _13235_, _13234_);
  and _44199_ (_13237_, _13236_, _02445_);
  or _44200_ (_13238_, _13237_, _13233_);
  and _44201_ (_13239_, _13238_, _02421_);
  or _44202_ (_13240_, _13239_, _13229_);
  and _44203_ (_13241_, _13240_, _02414_);
  and _44204_ (_13242_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and _44205_ (_13243_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or _44206_ (_13244_, _13243_, _13242_);
  and _44207_ (_13245_, _13244_, _02393_);
  and _44208_ (_13246_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and _44209_ (_13247_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or _44210_ (_13248_, _13247_, _13246_);
  and _44211_ (_13249_, _13248_, _02445_);
  or _44212_ (_13250_, _13249_, _13245_);
  and _44213_ (_13251_, _13250_, _02459_);
  and _44214_ (_13252_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and _44215_ (_13253_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or _44216_ (_13254_, _13253_, _13252_);
  and _44217_ (_13255_, _13254_, _02393_);
  and _44218_ (_13256_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and _44219_ (_13257_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or _44220_ (_13258_, _13257_, _13256_);
  and _44221_ (_13259_, _13258_, _02445_);
  or _44222_ (_13260_, _13259_, _13255_);
  and _44223_ (_13261_, _13260_, _02421_);
  or _44224_ (_13262_, _13261_, _13251_);
  and _44225_ (_13263_, _13262_, _02458_);
  or _44226_ (_13264_, _13263_, _13241_);
  and _44227_ (_13265_, _13264_, _02398_);
  or _44228_ (_13266_, _13265_, _13219_);
  and _44229_ (_13267_, _13266_, _02400_);
  and _44230_ (_13268_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and _44231_ (_13269_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or _44232_ (_13270_, _13269_, _13268_);
  and _44233_ (_13271_, _13270_, _02393_);
  and _44234_ (_13272_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and _44235_ (_13273_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or _44236_ (_13274_, _13273_, _13272_);
  and _44237_ (_13275_, _13274_, _02445_);
  or _44238_ (_13276_, _13275_, _13271_);
  or _44239_ (_13277_, _13276_, _02459_);
  and _44240_ (_13278_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and _44241_ (_13279_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or _44242_ (_13280_, _13279_, _13278_);
  and _44243_ (_13281_, _13280_, _02393_);
  and _44244_ (_13282_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and _44245_ (_13283_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or _44246_ (_13284_, _13283_, _13282_);
  and _44247_ (_13285_, _13284_, _02445_);
  or _44248_ (_13286_, _13285_, _13281_);
  or _44249_ (_13287_, _13286_, _02421_);
  and _44250_ (_13288_, _13287_, _02458_);
  and _44251_ (_13289_, _13288_, _13277_);
  or _44252_ (_13290_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or _44253_ (_13291_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and _44254_ (_13292_, _13291_, _13290_);
  and _44255_ (_13293_, _13292_, _02393_);
  or _44256_ (_13294_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or _44257_ (_13295_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and _44258_ (_13296_, _13295_, _13294_);
  and _44259_ (_13297_, _13296_, _02445_);
  or _44260_ (_13298_, _13297_, _13293_);
  or _44261_ (_13299_, _13298_, _02459_);
  or _44262_ (_13300_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or _44263_ (_13301_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and _44264_ (_13302_, _13301_, _13300_);
  and _44265_ (_13303_, _13302_, _02393_);
  or _44266_ (_13304_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or _44267_ (_13305_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and _44268_ (_13306_, _13305_, _13304_);
  and _44269_ (_13307_, _13306_, _02445_);
  or _44270_ (_13308_, _13307_, _13303_);
  or _44271_ (_13309_, _13308_, _02421_);
  and _44272_ (_13310_, _13309_, _02414_);
  and _44273_ (_13311_, _13310_, _13299_);
  or _44274_ (_13312_, _13311_, _13289_);
  and _44275_ (_13313_, _13312_, _02398_);
  and _44276_ (_13314_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and _44277_ (_13315_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or _44278_ (_13316_, _13315_, _13314_);
  and _44279_ (_13317_, _13316_, _02393_);
  and _44280_ (_13318_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and _44281_ (_13319_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or _44282_ (_13320_, _13319_, _13318_);
  and _44283_ (_13321_, _13320_, _02445_);
  or _44284_ (_13322_, _13321_, _13317_);
  or _44285_ (_13323_, _13322_, _02459_);
  and _44286_ (_13324_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and _44287_ (_13325_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or _44288_ (_13326_, _13325_, _13324_);
  and _44289_ (_13327_, _13326_, _02393_);
  and _44290_ (_13328_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and _44291_ (_13329_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or _44292_ (_13330_, _13329_, _13328_);
  and _44293_ (_13331_, _13330_, _02445_);
  or _44294_ (_13332_, _13331_, _13327_);
  or _44295_ (_13333_, _13332_, _02421_);
  and _44296_ (_13334_, _13333_, _02458_);
  and _44297_ (_13335_, _13334_, _13323_);
  or _44298_ (_13336_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or _44299_ (_13337_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and _44300_ (_13338_, _13337_, _02445_);
  and _44301_ (_13339_, _13338_, _13336_);
  or _44302_ (_13340_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or _44303_ (_13341_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and _44304_ (_13342_, _13341_, _02393_);
  and _44305_ (_13343_, _13342_, _13340_);
  or _44306_ (_13344_, _13343_, _13339_);
  or _44307_ (_13345_, _13344_, _02459_);
  or _44308_ (_13346_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or _44309_ (_13347_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and _44310_ (_13348_, _13347_, _02445_);
  and _44311_ (_13349_, _13348_, _13346_);
  or _44312_ (_13350_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or _44313_ (_13351_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and _44314_ (_13352_, _13351_, _02393_);
  and _44315_ (_13353_, _13352_, _13350_);
  or _44316_ (_13354_, _13353_, _13349_);
  or _44317_ (_13355_, _13354_, _02421_);
  and _44318_ (_13356_, _13355_, _02414_);
  and _44319_ (_13357_, _13356_, _13345_);
  or _44320_ (_13358_, _13357_, _13335_);
  and _44321_ (_13359_, _13358_, _02496_);
  or _44322_ (_13360_, _13359_, _13313_);
  and _44323_ (_13361_, _13360_, _02546_);
  or _44324_ (_13362_, _13361_, _13267_);
  and _44325_ (_13363_, _13362_, _02405_);
  or _44326_ (_13364_, _13363_, _13173_);
  and _44327_ (_13365_, _13364_, _26777_);
  and _44328_ (_13366_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and _44329_ (_13367_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or _44330_ (_13368_, _13367_, _13366_);
  and _44331_ (_13369_, _13368_, _02393_);
  and _44332_ (_13370_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and _44333_ (_13371_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or _44334_ (_13372_, _13371_, _13370_);
  and _44335_ (_13373_, _13372_, _02445_);
  or _44336_ (_13374_, _13373_, _13369_);
  and _44337_ (_13375_, _13374_, _02421_);
  and _44338_ (_13376_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and _44339_ (_13377_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or _44340_ (_13378_, _13377_, _13376_);
  and _44341_ (_13379_, _13378_, _02393_);
  and _44342_ (_13380_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  and _44343_ (_13381_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or _44344_ (_13382_, _13381_, _13380_);
  and _44345_ (_13383_, _13382_, _02445_);
  or _44346_ (_13384_, _13383_, _13379_);
  and _44347_ (_13385_, _13384_, _02459_);
  or _44348_ (_13386_, _13385_, _02414_);
  or _44349_ (_13387_, _13386_, _13375_);
  or _44350_ (_13388_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or _44351_ (_13389_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  and _44352_ (_13390_, _13389_, _13388_);
  and _44353_ (_13391_, _13390_, _02393_);
  or _44354_ (_13392_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or _44355_ (_13393_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and _44356_ (_13394_, _13393_, _13392_);
  and _44357_ (_13395_, _13394_, _02445_);
  or _44358_ (_13396_, _13395_, _13391_);
  and _44359_ (_13397_, _13396_, _02421_);
  or _44360_ (_13398_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or _44361_ (_13399_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  and _44362_ (_13400_, _13399_, _13398_);
  and _44363_ (_13401_, _13400_, _02393_);
  or _44364_ (_13402_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or _44365_ (_13403_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and _44366_ (_13404_, _13403_, _13402_);
  and _44367_ (_13405_, _13404_, _02445_);
  or _44368_ (_13406_, _13405_, _13401_);
  and _44369_ (_13407_, _13406_, _02459_);
  or _44370_ (_13408_, _13407_, _02458_);
  or _44371_ (_13409_, _13408_, _13397_);
  and _44372_ (_13410_, _13409_, _13387_);
  or _44373_ (_13411_, _13410_, _02496_);
  and _44374_ (_13412_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and _44375_ (_13413_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or _44376_ (_13414_, _13413_, _13412_);
  and _44377_ (_13415_, _13414_, _02393_);
  and _44378_ (_13416_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and _44379_ (_13417_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or _44380_ (_13418_, _13417_, _13416_);
  and _44381_ (_13419_, _13418_, _02445_);
  or _44382_ (_13420_, _13419_, _13415_);
  and _44383_ (_13421_, _13420_, _02421_);
  and _44384_ (_13422_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and _44385_ (_13423_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _44386_ (_13424_, _13423_, _13422_);
  and _44387_ (_13425_, _13424_, _02393_);
  and _44388_ (_13426_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and _44389_ (_13427_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or _44390_ (_13428_, _13427_, _13426_);
  and _44391_ (_13429_, _13428_, _02445_);
  or _44392_ (_13430_, _13429_, _13425_);
  and _44393_ (_13431_, _13430_, _02459_);
  or _44394_ (_13432_, _13431_, _02414_);
  or _44395_ (_13433_, _13432_, _13421_);
  or _44396_ (_13434_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or _44397_ (_13435_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and _44398_ (_13436_, _13435_, _02445_);
  and _44399_ (_13437_, _13436_, _13434_);
  or _44400_ (_13438_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or _44401_ (_13439_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and _44402_ (_13440_, _13439_, _02393_);
  and _44403_ (_13441_, _13440_, _13438_);
  or _44404_ (_13442_, _13441_, _13437_);
  and _44405_ (_13443_, _13442_, _02421_);
  or _44406_ (_13444_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or _44407_ (_13445_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and _44408_ (_13446_, _13445_, _02445_);
  and _44409_ (_13447_, _13446_, _13444_);
  or _44410_ (_13448_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or _44411_ (_13449_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and _44412_ (_13450_, _13449_, _02393_);
  and _44413_ (_13451_, _13450_, _13448_);
  or _44414_ (_13452_, _13451_, _13447_);
  and _44415_ (_13453_, _13452_, _02459_);
  or _44416_ (_13454_, _13453_, _02458_);
  or _44417_ (_13455_, _13454_, _13443_);
  and _44418_ (_13456_, _13455_, _13433_);
  or _44419_ (_13457_, _13456_, _02398_);
  and _44420_ (_13458_, _13457_, _13411_);
  and _44421_ (_13459_, _13458_, _02400_);
  and _44422_ (_13460_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and _44423_ (_13461_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or _44424_ (_13462_, _13461_, _13460_);
  and _44425_ (_13463_, _13462_, _02393_);
  and _44426_ (_13464_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and _44427_ (_13465_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or _44428_ (_13466_, _13465_, _13464_);
  and _44429_ (_13467_, _13466_, _02445_);
  or _44430_ (_13468_, _13467_, _13463_);
  or _44431_ (_13469_, _13468_, _02459_);
  and _44432_ (_13470_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and _44433_ (_13471_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or _44434_ (_13472_, _13471_, _13470_);
  and _44435_ (_13473_, _13472_, _02393_);
  and _44436_ (_13474_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and _44437_ (_13475_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or _44438_ (_13476_, _13475_, _13474_);
  and _44439_ (_13477_, _13476_, _02445_);
  or _44440_ (_13478_, _13477_, _13473_);
  or _44441_ (_13479_, _13478_, _02421_);
  and _44442_ (_13480_, _13479_, _02458_);
  and _44443_ (_13481_, _13480_, _13469_);
  or _44444_ (_13482_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or _44445_ (_13483_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  and _44446_ (_13484_, _13483_, _02445_);
  and _44447_ (_13485_, _13484_, _13482_);
  or _44448_ (_13486_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or _44449_ (_13487_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and _44450_ (_13488_, _13487_, _02393_);
  and _44451_ (_13489_, _13488_, _13486_);
  or _44452_ (_13490_, _13489_, _13485_);
  or _44453_ (_13491_, _13490_, _02459_);
  or _44454_ (_13492_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or _44455_ (_13493_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  and _44456_ (_13494_, _13493_, _02445_);
  and _44457_ (_13495_, _13494_, _13492_);
  or _44458_ (_13496_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or _44459_ (_13497_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and _44460_ (_13498_, _13497_, _02393_);
  and _44461_ (_13499_, _13498_, _13496_);
  or _44462_ (_13500_, _13499_, _13495_);
  or _44463_ (_13501_, _13500_, _02421_);
  and _44464_ (_13502_, _13501_, _02414_);
  and _44465_ (_13503_, _13502_, _13491_);
  or _44466_ (_13504_, _13503_, _13481_);
  or _44467_ (_13505_, _13504_, _02398_);
  and _44468_ (_13506_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and _44469_ (_13507_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or _44470_ (_13508_, _13507_, _13506_);
  and _44471_ (_13509_, _13508_, _02393_);
  and _44472_ (_13510_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and _44473_ (_13511_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or _44474_ (_13512_, _13511_, _13510_);
  and _44475_ (_13513_, _13512_, _02445_);
  or _44476_ (_13514_, _13513_, _13509_);
  or _44477_ (_13515_, _13514_, _02459_);
  and _44478_ (_13516_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and _44479_ (_13517_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or _44480_ (_13518_, _13517_, _13516_);
  and _44481_ (_13519_, _13518_, _02393_);
  and _44482_ (_13520_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  and _44483_ (_13521_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or _44484_ (_13522_, _13521_, _13520_);
  and _44485_ (_13523_, _13522_, _02445_);
  or _44486_ (_13524_, _13523_, _13519_);
  or _44487_ (_13525_, _13524_, _02421_);
  and _44488_ (_13526_, _13525_, _02458_);
  and _44489_ (_13527_, _13526_, _13515_);
  or _44490_ (_13528_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or _44491_ (_13529_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and _44492_ (_13530_, _13529_, _13528_);
  and _44493_ (_13531_, _13530_, _02393_);
  or _44494_ (_13532_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or _44495_ (_13533_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and _44496_ (_13534_, _13533_, _13532_);
  and _44497_ (_13535_, _13534_, _02445_);
  or _44498_ (_13536_, _13535_, _13531_);
  or _44499_ (_13537_, _13536_, _02459_);
  or _44500_ (_13538_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or _44501_ (_13539_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and _44502_ (_13540_, _13539_, _13538_);
  and _44503_ (_13541_, _13540_, _02393_);
  or _44504_ (_13542_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or _44505_ (_13543_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and _44506_ (_13544_, _13543_, _13542_);
  and _44507_ (_13545_, _13544_, _02445_);
  or _44508_ (_13546_, _13545_, _13541_);
  or _44509_ (_13547_, _13546_, _02421_);
  and _44510_ (_13548_, _13547_, _02414_);
  and _44511_ (_13549_, _13548_, _13537_);
  or _44512_ (_13550_, _13549_, _13527_);
  or _44513_ (_13551_, _13550_, _02496_);
  and _44514_ (_13552_, _13551_, _13505_);
  and _44515_ (_13553_, _13552_, _02546_);
  or _44516_ (_13554_, _13553_, _13459_);
  and _44517_ (_13555_, _13554_, _02646_);
  and _44518_ (_13556_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and _44519_ (_13557_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or _44520_ (_13558_, _13557_, _13556_);
  and _44521_ (_13559_, _13558_, _02445_);
  and _44522_ (_13560_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and _44523_ (_13561_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or _44524_ (_13562_, _13561_, _13560_);
  and _44525_ (_13563_, _13562_, _02393_);
  or _44526_ (_13564_, _13563_, _13559_);
  or _44527_ (_13565_, _13564_, _02459_);
  and _44528_ (_13566_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and _44529_ (_13567_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or _44530_ (_13568_, _13567_, _13566_);
  and _44531_ (_13569_, _13568_, _02445_);
  and _44532_ (_13570_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and _44533_ (_13571_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or _44534_ (_13572_, _13571_, _13570_);
  and _44535_ (_13573_, _13572_, _02393_);
  or _44536_ (_13574_, _13573_, _13569_);
  or _44537_ (_13575_, _13574_, _02421_);
  and _44538_ (_13576_, _13575_, _02458_);
  and _44539_ (_13577_, _13576_, _13565_);
  or _44540_ (_13578_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or _44541_ (_13579_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and _44542_ (_13580_, _13579_, _02393_);
  and _44543_ (_13581_, _13580_, _13578_);
  or _44544_ (_13582_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or _44545_ (_13583_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and _44546_ (_13584_, _13583_, _02445_);
  and _44547_ (_13585_, _13584_, _13582_);
  or _44548_ (_13586_, _13585_, _13581_);
  or _44549_ (_13587_, _13586_, _02459_);
  or _44550_ (_13588_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or _44551_ (_13589_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  and _44552_ (_13590_, _13589_, _02393_);
  and _44553_ (_13591_, _13590_, _13588_);
  or _44554_ (_13592_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or _44555_ (_13593_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  and _44556_ (_13594_, _13593_, _02445_);
  and _44557_ (_13595_, _13594_, _13592_);
  or _44558_ (_13596_, _13595_, _13591_);
  or _44559_ (_13597_, _13596_, _02421_);
  and _44560_ (_13598_, _13597_, _02414_);
  and _44561_ (_13599_, _13598_, _13587_);
  or _44562_ (_13600_, _13599_, _13577_);
  or _44563_ (_13601_, _13600_, _02398_);
  and _44564_ (_13602_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and _44565_ (_13603_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or _44566_ (_13604_, _13603_, _02393_);
  or _44567_ (_13605_, _13604_, _13602_);
  and _44568_ (_13606_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and _44569_ (_13607_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or _44570_ (_13608_, _13607_, _02445_);
  or _44571_ (_13609_, _13608_, _13606_);
  and _44572_ (_13610_, _13609_, _13605_);
  or _44573_ (_13611_, _13610_, _02459_);
  and _44574_ (_13612_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and _44575_ (_13613_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or _44576_ (_13614_, _13613_, _02393_);
  or _44577_ (_13615_, _13614_, _13612_);
  and _44578_ (_13616_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and _44579_ (_13617_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or _44580_ (_13618_, _13617_, _02445_);
  or _44581_ (_13619_, _13618_, _13616_);
  and _44582_ (_13620_, _13619_, _13615_);
  or _44583_ (_13621_, _13620_, _02421_);
  and _44584_ (_13622_, _13621_, _02458_);
  and _44585_ (_13623_, _13622_, _13611_);
  or _44586_ (_13624_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or _44587_ (_13625_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and _44588_ (_13626_, _13625_, _13624_);
  or _44589_ (_13627_, _13626_, _02445_);
  or _44590_ (_13628_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or _44591_ (_13629_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and _44592_ (_13630_, _13629_, _13628_);
  or _44593_ (_13631_, _13630_, _02393_);
  and _44594_ (_13632_, _13631_, _13627_);
  or _44595_ (_13633_, _13632_, _02459_);
  or _44596_ (_13634_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or _44597_ (_13635_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and _44598_ (_13636_, _13635_, _13634_);
  or _44599_ (_13637_, _13636_, _02445_);
  or _44600_ (_13638_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or _44601_ (_13639_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and _44602_ (_13640_, _13639_, _13638_);
  or _44603_ (_13641_, _13640_, _02393_);
  and _44604_ (_13642_, _13641_, _13637_);
  or _44605_ (_13643_, _13642_, _02421_);
  and _44606_ (_13644_, _13643_, _02414_);
  and _44607_ (_13645_, _13644_, _13633_);
  or _44608_ (_13646_, _13645_, _13623_);
  or _44609_ (_13647_, _13646_, _02496_);
  and _44610_ (_13648_, _13647_, _02546_);
  and _44611_ (_13649_, _13648_, _13601_);
  and _44612_ (_13650_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  and _44613_ (_13651_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or _44614_ (_13652_, _13651_, _13650_);
  and _44615_ (_13653_, _13652_, _02393_);
  and _44616_ (_13654_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and _44617_ (_13655_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or _44618_ (_13656_, _13655_, _13654_);
  and _44619_ (_13657_, _13656_, _02445_);
  or _44620_ (_13658_, _13657_, _13653_);
  and _44621_ (_13659_, _13658_, _02421_);
  and _44622_ (_13660_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  and _44623_ (_13661_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or _44624_ (_13662_, _13661_, _13660_);
  and _44625_ (_13663_, _13662_, _02393_);
  and _44626_ (_13664_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  and _44627_ (_13665_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or _44628_ (_13666_, _13665_, _13664_);
  and _44629_ (_13667_, _13666_, _02445_);
  or _44630_ (_13668_, _13667_, _13663_);
  and _44631_ (_13669_, _13668_, _02459_);
  or _44632_ (_13670_, _13669_, _02414_);
  or _44633_ (_13671_, _13670_, _13659_);
  or _44634_ (_13672_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or _44635_ (_13673_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and _44636_ (_13674_, _13673_, _13672_);
  and _44637_ (_13675_, _13674_, _02393_);
  or _44638_ (_13676_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or _44639_ (_13677_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and _44640_ (_13678_, _13677_, _13676_);
  and _44641_ (_13679_, _13678_, _02445_);
  or _44642_ (_13680_, _13679_, _13675_);
  and _44643_ (_13681_, _13680_, _02421_);
  or _44644_ (_13682_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or _44645_ (_13683_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  and _44646_ (_13684_, _13683_, _13682_);
  and _44647_ (_13685_, _13684_, _02393_);
  or _44648_ (_13686_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or _44649_ (_13687_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and _44650_ (_13688_, _13687_, _13686_);
  and _44651_ (_13689_, _13688_, _02445_);
  or _44652_ (_13690_, _13689_, _13685_);
  and _44653_ (_13691_, _13690_, _02459_);
  or _44654_ (_13692_, _13691_, _02458_);
  or _44655_ (_13693_, _13692_, _13681_);
  and _44656_ (_13694_, _13693_, _13671_);
  or _44657_ (_13695_, _13694_, _02496_);
  and _44658_ (_13696_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  and _44659_ (_13697_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  or _44660_ (_13698_, _13697_, _13696_);
  and _44661_ (_13699_, _13698_, _02393_);
  and _44662_ (_13700_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  and _44663_ (_13701_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  or _44664_ (_13702_, _13701_, _13700_);
  and _44665_ (_13703_, _13702_, _02445_);
  or _44666_ (_13704_, _13703_, _13699_);
  and _44667_ (_13705_, _13704_, _02421_);
  and _44668_ (_13706_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  and _44669_ (_13707_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or _44670_ (_13708_, _13707_, _13706_);
  and _44671_ (_13709_, _13708_, _02393_);
  and _44672_ (_13710_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  and _44673_ (_13711_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  or _44674_ (_13712_, _13711_, _13710_);
  and _44675_ (_13713_, _13712_, _02445_);
  or _44676_ (_13714_, _13713_, _13709_);
  and _44677_ (_13715_, _13714_, _02459_);
  or _44678_ (_13716_, _13715_, _02414_);
  or _44679_ (_13717_, _13716_, _13705_);
  or _44680_ (_13718_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or _44681_ (_13719_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  and _44682_ (_13720_, _13719_, _13718_);
  and _44683_ (_13721_, _13720_, _02393_);
  or _44684_ (_13722_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  or _44685_ (_13723_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  and _44686_ (_13724_, _13723_, _13722_);
  and _44687_ (_13725_, _13724_, _02445_);
  or _44688_ (_13726_, _13725_, _13721_);
  and _44689_ (_13727_, _13726_, _02421_);
  or _44690_ (_13728_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  or _44691_ (_13729_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  and _44692_ (_13730_, _13729_, _13728_);
  and _44693_ (_13731_, _13730_, _02393_);
  or _44694_ (_13732_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  or _44695_ (_13733_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  and _44696_ (_13734_, _13733_, _13732_);
  and _44697_ (_13735_, _13734_, _02445_);
  or _44698_ (_13736_, _13735_, _13731_);
  and _44699_ (_13737_, _13736_, _02459_);
  or _44700_ (_13738_, _13737_, _02458_);
  or _44701_ (_13739_, _13738_, _13727_);
  and _44702_ (_13740_, _13739_, _13717_);
  or _44703_ (_13741_, _13740_, _02398_);
  and _44704_ (_13742_, _13741_, _13695_);
  and _44705_ (_13743_, _13742_, _02400_);
  or _44706_ (_13744_, _13743_, _13649_);
  and _44707_ (_13745_, _13744_, _02405_);
  or _44708_ (_13746_, _13745_, _13555_);
  and _44709_ (_13747_, _13746_, _02444_);
  or _44710_ (_13748_, _13747_, _13365_);
  or _44711_ (_13749_, _13748_, _02443_);
  or _44712_ (_13750_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and _44713_ (_13751_, _13750_, _22762_);
  and _44714_ (_04033_, _13751_, _13749_);
  and _44715_ (_13752_, _05336_, _24329_);
  not _44716_ (_13753_, _13752_);
  and _44717_ (_13754_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  and _44718_ (_13755_, _13752_, _23946_);
  or _44719_ (_04045_, _13755_, _13754_);
  and _44720_ (_13756_, _06886_, _01808_);
  not _44721_ (_13757_, _13756_);
  and _44722_ (_13758_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and _44723_ (_13759_, _13756_, _23946_);
  or _44724_ (_04049_, _13759_, _13758_);
  nand _44725_ (_13760_, _24352_, _22767_);
  or _44726_ (_13761_, _22767_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _44727_ (_13762_, _13761_, _22762_);
  and _44728_ (_26864_[3], _13762_, _13760_);
  and _44729_ (_13763_, _24201_, _24005_);
  not _44730_ (_13764_, _13763_);
  and _44731_ (_13765_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and _44732_ (_13766_, _13763_, _23707_);
  or _44733_ (_04080_, _13766_, _13765_);
  and _44734_ (_13767_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and _44735_ (_13768_, _13756_, _23707_);
  or _44736_ (_04090_, _13768_, _13767_);
  and _44737_ (_13769_, _05336_, _25078_);
  not _44738_ (_13770_, _13769_);
  and _44739_ (_13771_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  and _44740_ (_13772_, _13769_, _23747_);
  or _44741_ (_27091_, _13772_, _13771_);
  and _44742_ (_13773_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  and _44743_ (_13774_, _13769_, _23898_);
  or _44744_ (_04098_, _13774_, _13773_);
  and _44745_ (_13775_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and _44746_ (_13776_, _13756_, _24050_);
  or _44747_ (_04111_, _13776_, _13775_);
  and _44748_ (_13777_, _05336_, _24282_);
  not _44749_ (_13778_, _13777_);
  and _44750_ (_13779_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and _44751_ (_13780_, _13777_, _23824_);
  or _44752_ (_04114_, _13780_, _13779_);
  and _44753_ (_13781_, _10347_, _23649_);
  and _44754_ (_13782_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  or _44755_ (_04117_, _13782_, _13781_);
  and _44756_ (_13783_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  and _44757_ (_13784_, _13752_, _23824_);
  or _44758_ (_04120_, _13784_, _13783_);
  and _44759_ (_13785_, _05336_, _23752_);
  not _44760_ (_13786_, _13785_);
  and _44761_ (_13787_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and _44762_ (_13788_, _13785_, _23707_);
  or _44763_ (_04125_, _13788_, _13787_);
  and _44764_ (_13789_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and _44765_ (_13790_, _13785_, _23649_);
  or _44766_ (_04133_, _13790_, _13789_);
  and _44767_ (_13791_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and _44768_ (_13792_, _12935_, _24050_);
  or _44769_ (_04140_, _13792_, _13791_);
  or _44770_ (_13793_, _24436_, _23837_);
  or _44771_ (_13794_, _22767_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _44772_ (_13795_, _13794_, _22762_);
  and _44773_ (_26864_[2], _13795_, _13793_);
  nand _44774_ (_13796_, _24486_, _22767_);
  or _44775_ (_13797_, _22767_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _44776_ (_13799_, _13797_, _22762_);
  and _44777_ (_26864_[6], _13799_, _13796_);
  and _44778_ (_13800_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  and _44779_ (_13801_, _12941_, _23898_);
  or _44780_ (_27100_, _13801_, _13800_);
  and _44781_ (_13802_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  and _44782_ (_13803_, _12970_, _24050_);
  or _44783_ (_04171_, _13803_, _13802_);
  and _44784_ (_13804_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  and _44785_ (_13805_, _12970_, _23747_);
  or _44786_ (_04174_, _13805_, _13804_);
  and _44787_ (_13806_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and _44788_ (_13807_, _12906_, _23778_);
  or _44789_ (_04193_, _13807_, _13806_);
  and _44790_ (_13808_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and _44791_ (_13809_, _12974_, _23898_);
  or _44792_ (_04195_, _13809_, _13808_);
  and _44793_ (_13810_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and _44794_ (_13811_, _12980_, _24050_);
  or _44795_ (_04199_, _13811_, _13810_);
  and _44796_ (_13812_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and _44797_ (_13813_, _12980_, _23778_);
  or _44798_ (_04203_, _13813_, _13812_);
  and _44799_ (_13814_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and _44800_ (_13815_, _13785_, _23778_);
  or _44801_ (_04209_, _13815_, _13814_);
  and _44802_ (_13816_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and _44803_ (_13817_, _12906_, _23898_);
  or _44804_ (_04212_, _13817_, _13816_);
  and _44805_ (_13818_, _05336_, _23656_);
  not _44806_ (_13819_, _13818_);
  and _44807_ (_13820_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  and _44808_ (_13821_, _13818_, _23747_);
  or _44809_ (_04214_, _13821_, _13820_);
  and _44810_ (_13822_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  and _44811_ (_13823_, _13818_, _23778_);
  or _44812_ (_04217_, _13823_, _13822_);
  and _44813_ (_13824_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and _44814_ (_13825_, _13777_, _23649_);
  or _44815_ (_04225_, _13825_, _13824_);
  and _44816_ (_13826_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and _44817_ (_13827_, _12935_, _23778_);
  or _44818_ (_04238_, _13827_, _13826_);
  and _44819_ (_13828_, _06886_, _24329_);
  not _44820_ (_13829_, _13828_);
  and _44821_ (_13830_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  and _44822_ (_13831_, _13828_, _23707_);
  or _44823_ (_04246_, _13831_, _13830_);
  and _44824_ (_13832_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and _44825_ (_13833_, _12974_, _23946_);
  or _44826_ (_04258_, _13833_, _13832_);
  and _44827_ (_13834_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and _44828_ (_13835_, _13756_, _23778_);
  or _44829_ (_04270_, _13835_, _13834_);
  and _44830_ (_13836_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  and _44831_ (_13837_, _13769_, _23946_);
  or _44832_ (_04275_, _13837_, _13836_);
  and _44833_ (_13838_, _05125_, _23898_);
  and _44834_ (_13839_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  or _44835_ (_04330_, _13839_, _13838_);
  and _44836_ (_13840_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and _44837_ (_13841_, _13785_, _23747_);
  or _44838_ (_04332_, _13841_, _13840_);
  and _44839_ (_13842_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and _44840_ (_13843_, _13785_, _23898_);
  or _44841_ (_04345_, _13843_, _13842_);
  and _44842_ (_13844_, _08043_, _23747_);
  and _44843_ (_13845_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or _44844_ (_27211_, _13845_, _13844_);
  and _44845_ (_13846_, _05288_, _23824_);
  and _44846_ (_13847_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  or _44847_ (_27056_, _13847_, _13846_);
  and _44848_ (_13848_, _05288_, _23778_);
  and _44849_ (_13849_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  or _44850_ (_04352_, _13849_, _13848_);
  and _44851_ (_13850_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and _44852_ (_13851_, _13756_, _23747_);
  or _44853_ (_04355_, _13851_, _13850_);
  and _44854_ (_13852_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and _44855_ (_13853_, _13785_, _23824_);
  or _44856_ (_04359_, _13853_, _13852_);
  and _44857_ (_13854_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  and _44858_ (_13855_, _01967_, _23946_);
  or _44859_ (_04364_, _13855_, _13854_);
  and _44860_ (_13856_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and _44861_ (_13857_, _13756_, _23824_);
  or _44862_ (_04371_, _13857_, _13856_);
  and _44863_ (_13858_, _12733_, _23707_);
  and _44864_ (_13859_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  or _44865_ (_04379_, _13859_, _13858_);
  and _44866_ (_13860_, _05288_, _23747_);
  and _44867_ (_13861_, _05290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  or _44868_ (_04382_, _13861_, _13860_);
  and _44869_ (_13862_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and _44870_ (_13863_, _13785_, _23946_);
  or _44871_ (_04385_, _13863_, _13862_);
  and _44872_ (_13864_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and _44873_ (_13865_, _13756_, _23898_);
  or _44874_ (_27012_, _13865_, _13864_);
  and _44875_ (_13866_, _05125_, _23946_);
  and _44876_ (_13867_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  or _44877_ (_27059_, _13867_, _13866_);
  and _44878_ (_13868_, _05125_, _23747_);
  and _44879_ (_13869_, _05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  or _44880_ (_04400_, _13869_, _13868_);
  and _44881_ (_13870_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and _44882_ (_13871_, _08351_, _23778_);
  or _44883_ (_04409_, _13871_, _13870_);
  and _44884_ (_13872_, _13786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and _44885_ (_13873_, _13785_, _24050_);
  or _44886_ (_04412_, _13873_, _13872_);
  and _44887_ (_13874_, _12733_, _24050_);
  and _44888_ (_13875_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  or _44889_ (_04419_, _13875_, _13874_);
  and _44890_ (_13876_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  and _44891_ (_13877_, _13752_, _23778_);
  or _44892_ (_04422_, _13877_, _13876_);
  and _44893_ (_13878_, _05008_, _23747_);
  and _44894_ (_13879_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or _44895_ (_04446_, _13879_, _13878_);
  and _44896_ (_13880_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  and _44897_ (_13881_, _13828_, _23898_);
  or _44898_ (_04450_, _13881_, _13880_);
  and _44899_ (_13882_, _05008_, _23707_);
  and _44900_ (_13883_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or _44901_ (_27062_, _13883_, _13882_);
  and _44902_ (_13884_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  and _44903_ (_13885_, _13752_, _23898_);
  or _44904_ (_04456_, _13885_, _13884_);
  and _44905_ (_13886_, _05008_, _24050_);
  and _44906_ (_13887_, _05011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or _44907_ (_27061_, _13887_, _13886_);
  and _44908_ (_13888_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  and _44909_ (_13889_, _13828_, _23778_);
  or _44910_ (_27010_, _13889_, _13888_);
  and _44911_ (_13890_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and _44912_ (_13891_, _13777_, _23898_);
  or _44913_ (_04468_, _13891_, _13890_);
  and _44914_ (_13892_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and _44915_ (_13893_, _13777_, _23747_);
  or _44916_ (_04472_, _13893_, _13892_);
  and _44917_ (_13894_, _06886_, _23752_);
  not _44918_ (_13895_, _13894_);
  and _44919_ (_13896_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and _44920_ (_13897_, _13894_, _23707_);
  or _44921_ (_04482_, _13897_, _13896_);
  and _44922_ (_13898_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and _44923_ (_13899_, _13777_, _23946_);
  or _44924_ (_04489_, _13899_, _13898_);
  and _44925_ (_13900_, _02246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  and _44926_ (_13901_, _02245_, _24050_);
  or _44927_ (_04492_, _13901_, _13900_);
  and _44928_ (_13902_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and _44929_ (_13903_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or _44930_ (_13904_, _13903_, _13902_);
  and _44931_ (_13905_, _13904_, _02393_);
  and _44932_ (_13906_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and _44933_ (_13907_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or _44934_ (_13908_, _13907_, _13906_);
  and _44935_ (_13909_, _13908_, _02445_);
  or _44936_ (_13910_, _13909_, _13905_);
  and _44937_ (_13911_, _13910_, _02421_);
  and _44938_ (_13912_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and _44939_ (_13913_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or _44940_ (_13914_, _13913_, _13912_);
  and _44941_ (_13915_, _13914_, _02393_);
  and _44942_ (_13916_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and _44943_ (_13917_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or _44944_ (_13918_, _13917_, _13916_);
  and _44945_ (_13919_, _13918_, _02445_);
  or _44946_ (_13920_, _13919_, _13915_);
  and _44947_ (_13921_, _13920_, _02459_);
  or _44948_ (_13922_, _13921_, _13911_);
  and _44949_ (_13923_, _13922_, _02458_);
  or _44950_ (_13924_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or _44951_ (_13925_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and _44952_ (_13926_, _13925_, _13924_);
  and _44953_ (_13927_, _13926_, _02393_);
  or _44954_ (_13928_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or _44955_ (_13929_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and _44956_ (_13930_, _13929_, _13928_);
  and _44957_ (_13931_, _13930_, _02445_);
  or _44958_ (_13932_, _13931_, _13927_);
  and _44959_ (_13933_, _13932_, _02421_);
  or _44960_ (_13934_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or _44961_ (_13935_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and _44962_ (_13936_, _13935_, _13934_);
  and _44963_ (_13937_, _13936_, _02393_);
  or _44964_ (_13938_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or _44965_ (_13939_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and _44966_ (_13940_, _13939_, _13938_);
  and _44967_ (_13941_, _13940_, _02445_);
  or _44968_ (_13942_, _13941_, _13937_);
  and _44969_ (_13943_, _13942_, _02459_);
  or _44970_ (_13944_, _13943_, _13933_);
  and _44971_ (_13945_, _13944_, _02414_);
  or _44972_ (_13946_, _13945_, _13923_);
  and _44973_ (_13947_, _13946_, _02398_);
  and _44974_ (_13948_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and _44975_ (_13949_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or _44976_ (_13950_, _13949_, _13948_);
  and _44977_ (_13951_, _13950_, _02393_);
  and _44978_ (_13952_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and _44979_ (_13953_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or _44980_ (_13954_, _13953_, _13952_);
  and _44981_ (_13955_, _13954_, _02445_);
  or _44982_ (_13956_, _13955_, _13951_);
  and _44983_ (_13957_, _13956_, _02421_);
  and _44984_ (_13958_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and _44985_ (_13959_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or _44986_ (_13960_, _13959_, _13958_);
  and _44987_ (_13961_, _13960_, _02393_);
  and _44988_ (_13962_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and _44989_ (_13963_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or _44990_ (_13964_, _13963_, _13962_);
  and _44991_ (_13965_, _13964_, _02445_);
  or _44992_ (_13966_, _13965_, _13961_);
  and _44993_ (_13967_, _13966_, _02459_);
  or _44994_ (_13968_, _13967_, _13957_);
  and _44995_ (_13969_, _13968_, _02458_);
  or _44996_ (_13970_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or _44997_ (_13971_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and _44998_ (_13972_, _13971_, _02445_);
  and _44999_ (_13973_, _13972_, _13970_);
  or _45000_ (_13974_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or _45001_ (_13975_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and _45002_ (_13976_, _13975_, _02393_);
  and _45003_ (_13977_, _13976_, _13974_);
  or _45004_ (_13978_, _13977_, _13973_);
  and _45005_ (_13979_, _13978_, _02421_);
  or _45006_ (_13980_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or _45007_ (_13981_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and _45008_ (_13982_, _13981_, _02445_);
  and _45009_ (_13983_, _13982_, _13980_);
  or _45010_ (_13984_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or _45011_ (_13985_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and _45012_ (_13986_, _13985_, _02393_);
  and _45013_ (_13987_, _13986_, _13984_);
  or _45014_ (_13988_, _13987_, _13983_);
  and _45015_ (_13989_, _13988_, _02459_);
  or _45016_ (_13990_, _13989_, _13979_);
  and _45017_ (_13991_, _13990_, _02414_);
  or _45018_ (_13992_, _13991_, _13969_);
  and _45019_ (_13993_, _13992_, _02496_);
  or _45020_ (_13994_, _13993_, _13947_);
  and _45021_ (_13995_, _13994_, _02400_);
  and _45022_ (_13996_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and _45023_ (_13997_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or _45024_ (_13998_, _13997_, _13996_);
  and _45025_ (_13999_, _13998_, _02393_);
  and _45026_ (_14000_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and _45027_ (_14001_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or _45028_ (_14002_, _14001_, _14000_);
  and _45029_ (_14003_, _14002_, _02445_);
  or _45030_ (_14004_, _14003_, _13999_);
  or _45031_ (_14005_, _14004_, _02459_);
  and _45032_ (_14006_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and _45033_ (_14007_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or _45034_ (_14008_, _14007_, _14006_);
  and _45035_ (_14009_, _14008_, _02393_);
  and _45036_ (_14010_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and _45037_ (_14011_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or _45038_ (_14012_, _14011_, _14010_);
  and _45039_ (_14013_, _14012_, _02445_);
  or _45040_ (_14014_, _14013_, _14009_);
  or _45041_ (_14015_, _14014_, _02421_);
  and _45042_ (_14016_, _14015_, _02458_);
  and _45043_ (_14017_, _14016_, _14005_);
  or _45044_ (_14018_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or _45045_ (_14019_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and _45046_ (_14020_, _14019_, _02445_);
  and _45047_ (_14021_, _14020_, _14018_);
  or _45048_ (_14022_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or _45049_ (_14023_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and _45050_ (_14024_, _14023_, _02393_);
  and _45051_ (_14025_, _14024_, _14022_);
  or _45052_ (_14026_, _14025_, _14021_);
  or _45053_ (_14027_, _14026_, _02459_);
  or _45054_ (_14028_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or _45055_ (_14029_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and _45056_ (_14030_, _14029_, _02445_);
  and _45057_ (_14031_, _14030_, _14028_);
  or _45058_ (_14032_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or _45059_ (_14033_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and _45060_ (_14034_, _14033_, _02393_);
  and _45061_ (_14035_, _14034_, _14032_);
  or _45062_ (_14036_, _14035_, _14031_);
  or _45063_ (_14037_, _14036_, _02421_);
  and _45064_ (_14038_, _14037_, _02414_);
  and _45065_ (_14039_, _14038_, _14027_);
  or _45066_ (_14040_, _14039_, _14017_);
  and _45067_ (_14041_, _14040_, _02496_);
  and _45068_ (_14042_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and _45069_ (_14043_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or _45070_ (_14044_, _14043_, _14042_);
  and _45071_ (_14045_, _14044_, _02393_);
  and _45072_ (_14046_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and _45073_ (_14047_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or _45074_ (_14048_, _14047_, _14046_);
  and _45075_ (_14049_, _14048_, _02445_);
  or _45076_ (_14050_, _14049_, _14045_);
  or _45077_ (_14051_, _14050_, _02459_);
  and _45078_ (_14052_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and _45079_ (_14053_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or _45080_ (_14054_, _14053_, _14052_);
  and _45081_ (_14055_, _14054_, _02393_);
  and _45082_ (_14056_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and _45083_ (_14057_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or _45084_ (_14058_, _14057_, _14056_);
  and _45085_ (_14059_, _14058_, _02445_);
  or _45086_ (_14060_, _14059_, _14055_);
  or _45087_ (_14061_, _14060_, _02421_);
  and _45088_ (_14062_, _14061_, _02458_);
  and _45089_ (_14063_, _14062_, _14051_);
  or _45090_ (_14064_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or _45091_ (_14065_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and _45092_ (_14066_, _14065_, _14064_);
  and _45093_ (_14067_, _14066_, _02393_);
  or _45094_ (_14068_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or _45095_ (_14069_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and _45096_ (_14070_, _14069_, _14068_);
  and _45097_ (_14071_, _14070_, _02445_);
  or _45098_ (_14072_, _14071_, _14067_);
  or _45099_ (_14073_, _14072_, _02459_);
  or _45100_ (_14074_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or _45101_ (_14075_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and _45102_ (_14076_, _14075_, _14074_);
  and _45103_ (_14077_, _14076_, _02393_);
  or _45104_ (_14078_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or _45105_ (_14079_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and _45106_ (_14080_, _14079_, _14078_);
  and _45107_ (_14081_, _14080_, _02445_);
  or _45108_ (_14082_, _14081_, _14077_);
  or _45109_ (_14083_, _14082_, _02421_);
  and _45110_ (_14084_, _14083_, _02414_);
  and _45111_ (_14085_, _14084_, _14073_);
  or _45112_ (_14086_, _14085_, _14063_);
  and _45113_ (_14087_, _14086_, _02398_);
  or _45114_ (_14088_, _14087_, _14041_);
  and _45115_ (_14089_, _14088_, _02546_);
  or _45116_ (_14090_, _14089_, _13995_);
  and _45117_ (_14091_, _14090_, _02646_);
  or _45118_ (_14092_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or _45119_ (_14093_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and _45120_ (_14094_, _14093_, _02445_);
  and _45121_ (_14095_, _14094_, _14092_);
  or _45122_ (_14096_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or _45123_ (_14097_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and _45124_ (_14098_, _14097_, _02393_);
  and _45125_ (_14099_, _14098_, _14096_);
  or _45126_ (_14100_, _14099_, _14095_);
  and _45127_ (_14101_, _14100_, _02459_);
  or _45128_ (_14102_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or _45129_ (_14103_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and _45130_ (_14104_, _14103_, _02445_);
  and _45131_ (_14105_, _14104_, _14102_);
  or _45132_ (_14106_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or _45133_ (_14107_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and _45134_ (_14108_, _14107_, _02393_);
  and _45135_ (_14109_, _14108_, _14106_);
  or _45136_ (_14110_, _14109_, _14105_);
  and _45137_ (_14111_, _14110_, _02421_);
  or _45138_ (_14112_, _14111_, _14101_);
  and _45139_ (_14113_, _14112_, _02414_);
  and _45140_ (_14114_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and _45141_ (_14115_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or _45142_ (_14116_, _14115_, _14114_);
  and _45143_ (_14117_, _14116_, _02393_);
  and _45144_ (_14118_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and _45145_ (_14119_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or _45146_ (_14120_, _14119_, _14118_);
  and _45147_ (_14121_, _14120_, _02445_);
  or _45148_ (_14122_, _14121_, _14117_);
  and _45149_ (_14123_, _14122_, _02459_);
  and _45150_ (_14124_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and _45151_ (_14125_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or _45152_ (_14126_, _14125_, _14124_);
  and _45153_ (_14127_, _14126_, _02393_);
  and _45154_ (_14128_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and _45155_ (_14129_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or _45156_ (_14130_, _14129_, _14128_);
  and _45157_ (_14131_, _14130_, _02445_);
  or _45158_ (_14132_, _14131_, _14127_);
  and _45159_ (_14133_, _14132_, _02421_);
  or _45160_ (_14134_, _14133_, _14123_);
  and _45161_ (_14135_, _14134_, _02458_);
  or _45162_ (_14136_, _14135_, _14113_);
  and _45163_ (_14137_, _14136_, _02496_);
  or _45164_ (_14138_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or _45165_ (_14139_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and _45166_ (_14140_, _14139_, _14138_);
  and _45167_ (_14141_, _14140_, _02393_);
  or _45168_ (_14142_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or _45169_ (_14143_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and _45170_ (_14144_, _14143_, _14142_);
  and _45171_ (_14145_, _14144_, _02445_);
  or _45172_ (_14146_, _14145_, _14141_);
  and _45173_ (_14147_, _14146_, _02459_);
  or _45174_ (_14148_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or _45175_ (_14149_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and _45176_ (_14150_, _14149_, _14148_);
  and _45177_ (_14151_, _14150_, _02393_);
  or _45178_ (_14152_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or _45179_ (_14153_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and _45180_ (_14154_, _14153_, _14152_);
  and _45181_ (_14155_, _14154_, _02445_);
  or _45182_ (_14156_, _14155_, _14151_);
  and _45183_ (_14157_, _14156_, _02421_);
  or _45184_ (_14158_, _14157_, _14147_);
  and _45185_ (_14159_, _14158_, _02414_);
  and _45186_ (_14160_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and _45187_ (_14161_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or _45188_ (_14162_, _14161_, _14160_);
  and _45189_ (_14163_, _14162_, _02393_);
  and _45190_ (_14164_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and _45191_ (_14165_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or _45192_ (_14166_, _14165_, _14164_);
  and _45193_ (_14167_, _14166_, _02445_);
  or _45194_ (_14168_, _14167_, _14163_);
  and _45195_ (_14169_, _14168_, _02459_);
  and _45196_ (_14170_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and _45197_ (_14171_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or _45198_ (_14172_, _14171_, _14170_);
  and _45199_ (_14173_, _14172_, _02393_);
  and _45200_ (_14174_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and _45201_ (_14175_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or _45202_ (_14176_, _14175_, _14174_);
  and _45203_ (_14177_, _14176_, _02445_);
  or _45204_ (_14178_, _14177_, _14173_);
  and _45205_ (_14179_, _14178_, _02421_);
  or _45206_ (_14180_, _14179_, _14169_);
  and _45207_ (_14181_, _14180_, _02458_);
  or _45208_ (_14182_, _14181_, _14159_);
  and _45209_ (_14183_, _14182_, _02398_);
  or _45210_ (_14184_, _14183_, _14137_);
  and _45211_ (_14185_, _14184_, _02400_);
  and _45212_ (_14186_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and _45213_ (_14187_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or _45214_ (_14188_, _14187_, _14186_);
  and _45215_ (_14189_, _14188_, _02393_);
  and _45216_ (_14190_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and _45217_ (_14191_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or _45218_ (_14192_, _14191_, _14190_);
  and _45219_ (_14193_, _14192_, _02445_);
  or _45220_ (_14194_, _14193_, _14189_);
  or _45221_ (_14195_, _14194_, _02459_);
  and _45222_ (_14196_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and _45223_ (_14197_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or _45224_ (_14198_, _14197_, _14196_);
  and _45225_ (_14199_, _14198_, _02393_);
  and _45226_ (_14200_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and _45227_ (_14201_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or _45228_ (_14202_, _14201_, _14200_);
  and _45229_ (_14203_, _14202_, _02445_);
  or _45230_ (_14204_, _14203_, _14199_);
  or _45231_ (_14205_, _14204_, _02421_);
  and _45232_ (_14206_, _14205_, _02458_);
  and _45233_ (_14207_, _14206_, _14195_);
  or _45234_ (_14208_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or _45235_ (_14209_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and _45236_ (_14210_, _14209_, _14208_);
  and _45237_ (_14211_, _14210_, _02393_);
  or _45238_ (_14212_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or _45239_ (_14213_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and _45240_ (_14214_, _14213_, _14212_);
  and _45241_ (_14215_, _14214_, _02445_);
  or _45242_ (_14216_, _14215_, _14211_);
  or _45243_ (_14217_, _14216_, _02459_);
  or _45244_ (_14218_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or _45245_ (_14219_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and _45246_ (_14220_, _14219_, _14218_);
  and _45247_ (_14221_, _14220_, _02393_);
  or _45248_ (_14222_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or _45249_ (_14223_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and _45250_ (_14224_, _14223_, _14222_);
  and _45251_ (_14225_, _14224_, _02445_);
  or _45252_ (_14226_, _14225_, _14221_);
  or _45253_ (_14227_, _14226_, _02421_);
  and _45254_ (_14228_, _14227_, _02414_);
  and _45255_ (_14229_, _14228_, _14217_);
  or _45256_ (_14230_, _14229_, _14207_);
  and _45257_ (_14231_, _14230_, _02398_);
  and _45258_ (_14232_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and _45259_ (_14233_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or _45260_ (_14234_, _14233_, _14232_);
  and _45261_ (_14235_, _14234_, _02393_);
  and _45262_ (_14236_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and _45263_ (_14237_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or _45264_ (_14238_, _14237_, _14236_);
  and _45265_ (_14239_, _14238_, _02445_);
  or _45266_ (_14240_, _14239_, _14235_);
  or _45267_ (_14241_, _14240_, _02459_);
  and _45268_ (_14242_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and _45269_ (_14243_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or _45270_ (_14244_, _14243_, _14242_);
  and _45271_ (_14245_, _14244_, _02393_);
  and _45272_ (_14246_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and _45273_ (_14247_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or _45274_ (_14248_, _14247_, _14246_);
  and _45275_ (_14249_, _14248_, _02445_);
  or _45276_ (_14250_, _14249_, _14245_);
  or _45277_ (_14251_, _14250_, _02421_);
  and _45278_ (_14252_, _14251_, _02458_);
  and _45279_ (_14253_, _14252_, _14241_);
  or _45280_ (_14254_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or _45281_ (_14255_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and _45282_ (_14256_, _14255_, _02445_);
  and _45283_ (_14257_, _14256_, _14254_);
  or _45284_ (_14258_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or _45285_ (_14259_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and _45286_ (_14260_, _14259_, _02393_);
  and _45287_ (_14261_, _14260_, _14258_);
  or _45288_ (_14262_, _14261_, _14257_);
  or _45289_ (_14263_, _14262_, _02459_);
  or _45290_ (_14264_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or _45291_ (_14265_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and _45292_ (_14266_, _14265_, _02445_);
  and _45293_ (_14267_, _14266_, _14264_);
  or _45294_ (_14268_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or _45295_ (_14269_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and _45296_ (_14270_, _14269_, _02393_);
  and _45297_ (_14271_, _14270_, _14268_);
  or _45298_ (_14272_, _14271_, _14267_);
  or _45299_ (_14273_, _14272_, _02421_);
  and _45300_ (_14274_, _14273_, _02414_);
  and _45301_ (_14275_, _14274_, _14263_);
  or _45302_ (_14276_, _14275_, _14253_);
  and _45303_ (_14277_, _14276_, _02496_);
  or _45304_ (_14278_, _14277_, _14231_);
  and _45305_ (_14279_, _14278_, _02546_);
  or _45306_ (_14280_, _14279_, _14185_);
  and _45307_ (_14281_, _14280_, _02405_);
  or _45308_ (_14282_, _14281_, _14091_);
  and _45309_ (_14283_, _14282_, _26777_);
  and _45310_ (_14284_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and _45311_ (_14285_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or _45312_ (_14286_, _14285_, _14284_);
  and _45313_ (_14287_, _14286_, _02393_);
  and _45314_ (_14288_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and _45315_ (_14289_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or _45316_ (_14290_, _14289_, _14288_);
  and _45317_ (_14291_, _14290_, _02445_);
  or _45318_ (_14292_, _14291_, _14287_);
  and _45319_ (_14293_, _14292_, _02421_);
  and _45320_ (_14294_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and _45321_ (_14295_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or _45322_ (_14296_, _14295_, _14294_);
  and _45323_ (_14297_, _14296_, _02393_);
  and _45324_ (_14298_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  and _45325_ (_14299_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or _45326_ (_14300_, _14299_, _14298_);
  and _45327_ (_14301_, _14300_, _02445_);
  or _45328_ (_14302_, _14301_, _14297_);
  and _45329_ (_14303_, _14302_, _02459_);
  or _45330_ (_14304_, _14303_, _02414_);
  or _45331_ (_14305_, _14304_, _14293_);
  or _45332_ (_14306_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or _45333_ (_14307_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  and _45334_ (_14308_, _14307_, _14306_);
  and _45335_ (_14309_, _14308_, _02393_);
  or _45336_ (_14310_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or _45337_ (_14311_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and _45338_ (_14312_, _14311_, _14310_);
  and _45339_ (_14313_, _14312_, _02445_);
  or _45340_ (_14314_, _14313_, _14309_);
  and _45341_ (_14315_, _14314_, _02421_);
  or _45342_ (_14316_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or _45343_ (_14317_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and _45344_ (_14318_, _14317_, _14316_);
  and _45345_ (_14319_, _14318_, _02393_);
  or _45346_ (_14320_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or _45347_ (_14321_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and _45348_ (_14322_, _14321_, _14320_);
  and _45349_ (_14323_, _14322_, _02445_);
  or _45350_ (_14324_, _14323_, _14319_);
  and _45351_ (_14325_, _14324_, _02459_);
  or _45352_ (_14326_, _14325_, _02458_);
  or _45353_ (_14327_, _14326_, _14315_);
  and _45354_ (_14328_, _14327_, _14305_);
  or _45355_ (_14329_, _14328_, _02496_);
  and _45356_ (_14330_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and _45357_ (_14331_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or _45358_ (_14332_, _14331_, _14330_);
  and _45359_ (_14333_, _14332_, _02393_);
  and _45360_ (_14334_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and _45361_ (_14335_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or _45362_ (_14336_, _14335_, _14334_);
  and _45363_ (_14337_, _14336_, _02445_);
  or _45364_ (_14338_, _14337_, _14333_);
  and _45365_ (_14339_, _14338_, _02421_);
  and _45366_ (_14340_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and _45367_ (_14341_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _45368_ (_14342_, _14341_, _14340_);
  and _45369_ (_14343_, _14342_, _02393_);
  and _45370_ (_14344_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and _45371_ (_14345_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or _45372_ (_14346_, _14345_, _14344_);
  and _45373_ (_14347_, _14346_, _02445_);
  or _45374_ (_14348_, _14347_, _14343_);
  and _45375_ (_14349_, _14348_, _02459_);
  or _45376_ (_14350_, _14349_, _02414_);
  or _45377_ (_14351_, _14350_, _14339_);
  or _45378_ (_14352_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or _45379_ (_14353_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and _45380_ (_14354_, _14353_, _02445_);
  and _45381_ (_14355_, _14354_, _14352_);
  or _45382_ (_14356_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or _45383_ (_14357_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and _45384_ (_14358_, _14357_, _02393_);
  and _45385_ (_14359_, _14358_, _14356_);
  or _45386_ (_14360_, _14359_, _14355_);
  and _45387_ (_14361_, _14360_, _02421_);
  or _45388_ (_14362_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or _45389_ (_14363_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and _45390_ (_14364_, _14363_, _02445_);
  and _45391_ (_14365_, _14364_, _14362_);
  or _45392_ (_14366_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or _45393_ (_14367_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and _45394_ (_14368_, _14367_, _02393_);
  and _45395_ (_14369_, _14368_, _14366_);
  or _45396_ (_14370_, _14369_, _14365_);
  and _45397_ (_14371_, _14370_, _02459_);
  or _45398_ (_14372_, _14371_, _02458_);
  or _45399_ (_14373_, _14372_, _14361_);
  and _45400_ (_14374_, _14373_, _14351_);
  or _45401_ (_14375_, _14374_, _02398_);
  and _45402_ (_14376_, _14375_, _14329_);
  and _45403_ (_14377_, _14376_, _02400_);
  and _45404_ (_14378_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and _45405_ (_14379_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or _45406_ (_14380_, _14379_, _14378_);
  and _45407_ (_14381_, _14380_, _02393_);
  and _45408_ (_14382_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and _45409_ (_14383_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or _45410_ (_14384_, _14383_, _14382_);
  and _45411_ (_14385_, _14384_, _02445_);
  or _45412_ (_14386_, _14385_, _14381_);
  or _45413_ (_14387_, _14386_, _02459_);
  and _45414_ (_14388_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  and _45415_ (_14389_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or _45416_ (_14390_, _14389_, _14388_);
  and _45417_ (_14391_, _14390_, _02393_);
  and _45418_ (_14392_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and _45419_ (_14393_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or _45420_ (_14394_, _14393_, _14392_);
  and _45421_ (_14395_, _14394_, _02445_);
  or _45422_ (_14396_, _14395_, _14391_);
  or _45423_ (_14397_, _14396_, _02421_);
  and _45424_ (_14398_, _14397_, _02458_);
  and _45425_ (_14399_, _14398_, _14387_);
  or _45426_ (_14400_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or _45427_ (_14401_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and _45428_ (_14402_, _14401_, _02445_);
  and _45429_ (_14403_, _14402_, _14400_);
  or _45430_ (_14404_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or _45431_ (_14405_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and _45432_ (_14406_, _14405_, _02393_);
  and _45433_ (_14407_, _14406_, _14404_);
  or _45434_ (_14408_, _14407_, _14403_);
  or _45435_ (_14409_, _14408_, _02459_);
  or _45436_ (_14410_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or _45437_ (_14411_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  and _45438_ (_14412_, _14411_, _02445_);
  and _45439_ (_14413_, _14412_, _14410_);
  or _45440_ (_14414_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or _45441_ (_14415_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and _45442_ (_14416_, _14415_, _02393_);
  and _45443_ (_14417_, _14416_, _14414_);
  or _45444_ (_14418_, _14417_, _14413_);
  or _45445_ (_14419_, _14418_, _02421_);
  and _45446_ (_14420_, _14419_, _02414_);
  and _45447_ (_14421_, _14420_, _14409_);
  or _45448_ (_14422_, _14421_, _14399_);
  or _45449_ (_14423_, _14422_, _02398_);
  and _45450_ (_14424_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and _45451_ (_14425_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or _45452_ (_14426_, _14425_, _14424_);
  and _45453_ (_14427_, _14426_, _02393_);
  and _45454_ (_14428_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and _45455_ (_14429_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or _45456_ (_14430_, _14429_, _14428_);
  and _45457_ (_14431_, _14430_, _02445_);
  or _45458_ (_14432_, _14431_, _14427_);
  or _45459_ (_14433_, _14432_, _02459_);
  and _45460_ (_14434_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and _45461_ (_14435_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or _45462_ (_14436_, _14435_, _14434_);
  and _45463_ (_14437_, _14436_, _02393_);
  and _45464_ (_14438_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  and _45465_ (_14439_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or _45466_ (_14440_, _14439_, _14438_);
  and _45467_ (_14441_, _14440_, _02445_);
  or _45468_ (_14442_, _14441_, _14437_);
  or _45469_ (_14443_, _14442_, _02421_);
  and _45470_ (_14444_, _14443_, _02458_);
  and _45471_ (_14445_, _14444_, _14433_);
  or _45472_ (_14446_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or _45473_ (_14447_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  and _45474_ (_14448_, _14447_, _14446_);
  and _45475_ (_14449_, _14448_, _02393_);
  or _45476_ (_14451_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or _45477_ (_14452_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and _45478_ (_14453_, _14452_, _14451_);
  and _45479_ (_14454_, _14453_, _02445_);
  or _45480_ (_14455_, _14454_, _14449_);
  or _45481_ (_14456_, _14455_, _02459_);
  or _45482_ (_14457_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or _45483_ (_14458_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and _45484_ (_14459_, _14458_, _14457_);
  and _45485_ (_14460_, _14459_, _02393_);
  or _45486_ (_14461_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or _45487_ (_14462_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and _45488_ (_14463_, _14462_, _14461_);
  and _45489_ (_14464_, _14463_, _02445_);
  or _45490_ (_14465_, _14464_, _14460_);
  or _45491_ (_14466_, _14465_, _02421_);
  and _45492_ (_14467_, _14466_, _02414_);
  and _45493_ (_14468_, _14467_, _14456_);
  or _45494_ (_14469_, _14468_, _14445_);
  or _45495_ (_14470_, _14469_, _02496_);
  and _45496_ (_14471_, _14470_, _14423_);
  and _45497_ (_14472_, _14471_, _02546_);
  or _45498_ (_14473_, _14472_, _14377_);
  and _45499_ (_14474_, _14473_, _02646_);
  and _45500_ (_14475_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  and _45501_ (_14476_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or _45502_ (_14477_, _14476_, _14475_);
  and _45503_ (_14478_, _14477_, _02445_);
  and _45504_ (_14479_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and _45505_ (_14480_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or _45506_ (_14481_, _14480_, _14479_);
  and _45507_ (_14482_, _14481_, _02393_);
  or _45508_ (_14483_, _14482_, _14478_);
  or _45509_ (_14484_, _14483_, _02459_);
  and _45510_ (_14485_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and _45511_ (_14486_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or _45512_ (_14487_, _14486_, _14485_);
  and _45513_ (_14488_, _14487_, _02445_);
  and _45514_ (_14489_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and _45515_ (_14490_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or _45516_ (_14491_, _14490_, _14489_);
  and _45517_ (_14492_, _14491_, _02393_);
  or _45518_ (_14493_, _14492_, _14488_);
  or _45519_ (_14494_, _14493_, _02421_);
  and _45520_ (_14495_, _14494_, _02458_);
  and _45521_ (_14496_, _14495_, _14484_);
  or _45522_ (_14497_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or _45523_ (_14498_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and _45524_ (_14499_, _14498_, _02393_);
  and _45525_ (_14500_, _14499_, _14497_);
  or _45526_ (_14501_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or _45527_ (_14502_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  and _45528_ (_14503_, _14502_, _02445_);
  and _45529_ (_14504_, _14503_, _14501_);
  or _45530_ (_14505_, _14504_, _14500_);
  or _45531_ (_14506_, _14505_, _02459_);
  or _45532_ (_14507_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or _45533_ (_14508_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and _45534_ (_14509_, _14508_, _02393_);
  and _45535_ (_14510_, _14509_, _14507_);
  or _45536_ (_14511_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or _45537_ (_14512_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  and _45538_ (_14513_, _14512_, _02445_);
  and _45539_ (_14514_, _14513_, _14511_);
  or _45540_ (_14515_, _14514_, _14510_);
  or _45541_ (_14516_, _14515_, _02421_);
  and _45542_ (_14517_, _14516_, _02414_);
  and _45543_ (_14518_, _14517_, _14506_);
  or _45544_ (_14519_, _14518_, _14496_);
  or _45545_ (_14520_, _14519_, _02398_);
  and _45546_ (_14521_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and _45547_ (_14522_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or _45548_ (_14523_, _14522_, _02393_);
  or _45549_ (_14524_, _14523_, _14521_);
  and _45550_ (_14525_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and _45551_ (_14526_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or _45552_ (_14527_, _14526_, _02445_);
  or _45553_ (_14528_, _14527_, _14525_);
  and _45554_ (_14529_, _14528_, _14524_);
  or _45555_ (_14530_, _14529_, _02459_);
  and _45556_ (_14531_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and _45557_ (_14532_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or _45558_ (_14533_, _14532_, _02393_);
  or _45559_ (_14534_, _14533_, _14531_);
  and _45560_ (_14535_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and _45561_ (_14536_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or _45562_ (_14537_, _14536_, _02445_);
  or _45563_ (_14538_, _14537_, _14535_);
  and _45564_ (_14539_, _14538_, _14534_);
  or _45565_ (_14540_, _14539_, _02421_);
  and _45566_ (_14541_, _14540_, _02458_);
  and _45567_ (_14542_, _14541_, _14530_);
  or _45568_ (_14543_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or _45569_ (_14544_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and _45570_ (_14545_, _14544_, _14543_);
  or _45571_ (_14546_, _14545_, _02445_);
  or _45572_ (_14547_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or _45573_ (_14548_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and _45574_ (_14549_, _14548_, _14547_);
  or _45575_ (_14550_, _14549_, _02393_);
  and _45576_ (_14551_, _14550_, _14546_);
  or _45577_ (_14552_, _14551_, _02459_);
  or _45578_ (_14553_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or _45579_ (_14554_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and _45580_ (_14555_, _14554_, _14553_);
  or _45581_ (_14556_, _14555_, _02445_);
  or _45582_ (_14557_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or _45583_ (_14558_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and _45584_ (_14559_, _14558_, _14557_);
  or _45585_ (_14560_, _14559_, _02393_);
  and _45586_ (_14561_, _14560_, _14556_);
  or _45587_ (_14562_, _14561_, _02421_);
  and _45588_ (_14563_, _14562_, _02414_);
  and _45589_ (_14564_, _14563_, _14552_);
  or _45590_ (_14565_, _14564_, _14542_);
  or _45591_ (_14566_, _14565_, _02496_);
  and _45592_ (_14567_, _14566_, _02546_);
  and _45593_ (_14568_, _14567_, _14520_);
  and _45594_ (_14569_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and _45595_ (_14570_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or _45596_ (_14571_, _14570_, _14569_);
  and _45597_ (_14572_, _14571_, _02393_);
  and _45598_ (_14573_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and _45599_ (_14574_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or _45600_ (_14575_, _14574_, _14573_);
  and _45601_ (_14576_, _14575_, _02445_);
  or _45602_ (_14577_, _14576_, _14572_);
  and _45603_ (_14578_, _14577_, _02421_);
  and _45604_ (_14579_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  and _45605_ (_14580_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or _45606_ (_14581_, _14580_, _14579_);
  and _45607_ (_14582_, _14581_, _02393_);
  and _45608_ (_14583_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and _45609_ (_14584_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or _45610_ (_14585_, _14584_, _14583_);
  and _45611_ (_14586_, _14585_, _02445_);
  or _45612_ (_14587_, _14586_, _14582_);
  and _45613_ (_14588_, _14587_, _02459_);
  or _45614_ (_14589_, _14588_, _02414_);
  or _45615_ (_14590_, _14589_, _14578_);
  or _45616_ (_14591_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or _45617_ (_14592_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and _45618_ (_14593_, _14592_, _14591_);
  and _45619_ (_14594_, _14593_, _02393_);
  or _45620_ (_14595_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or _45621_ (_14596_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and _45622_ (_14597_, _14596_, _14595_);
  and _45623_ (_14598_, _14597_, _02445_);
  or _45624_ (_14599_, _14598_, _14594_);
  and _45625_ (_14600_, _14599_, _02421_);
  or _45626_ (_14602_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or _45627_ (_14603_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and _45628_ (_14604_, _14603_, _14602_);
  and _45629_ (_14605_, _14604_, _02393_);
  or _45630_ (_14606_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or _45631_ (_14607_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  and _45632_ (_14608_, _14607_, _14606_);
  and _45633_ (_14609_, _14608_, _02445_);
  or _45634_ (_14610_, _14609_, _14605_);
  and _45635_ (_14611_, _14610_, _02459_);
  or _45636_ (_14612_, _14611_, _02458_);
  or _45637_ (_14613_, _14612_, _14600_);
  and _45638_ (_14614_, _14613_, _14590_);
  or _45639_ (_14615_, _14614_, _02496_);
  and _45640_ (_14616_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  and _45641_ (_14617_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or _45642_ (_14618_, _14617_, _14616_);
  and _45643_ (_14619_, _14618_, _02393_);
  and _45644_ (_14620_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  and _45645_ (_14621_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  or _45646_ (_14622_, _14621_, _14620_);
  and _45647_ (_14623_, _14622_, _02445_);
  or _45648_ (_14624_, _14623_, _14619_);
  and _45649_ (_14625_, _14624_, _02421_);
  and _45650_ (_14626_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  and _45651_ (_14627_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or _45652_ (_14628_, _14627_, _14626_);
  and _45653_ (_14629_, _14628_, _02393_);
  and _45654_ (_14630_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  and _45655_ (_14631_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  or _45656_ (_14632_, _14631_, _14630_);
  and _45657_ (_14633_, _14632_, _02445_);
  or _45658_ (_14634_, _14633_, _14629_);
  and _45659_ (_14635_, _14634_, _02459_);
  or _45660_ (_14636_, _14635_, _02414_);
  or _45661_ (_14637_, _14636_, _14625_);
  or _45662_ (_14638_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or _45663_ (_14639_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  and _45664_ (_14640_, _14639_, _14638_);
  and _45665_ (_14641_, _14640_, _02393_);
  or _45666_ (_14642_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  or _45667_ (_14643_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  and _45668_ (_14644_, _14643_, _14642_);
  and _45669_ (_14645_, _14644_, _02445_);
  or _45670_ (_14646_, _14645_, _14641_);
  and _45671_ (_14647_, _14646_, _02421_);
  or _45672_ (_14648_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or _45673_ (_14649_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  and _45674_ (_14650_, _14649_, _14648_);
  and _45675_ (_14651_, _14650_, _02393_);
  or _45676_ (_14652_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or _45677_ (_14653_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  and _45678_ (_14654_, _14653_, _14652_);
  and _45679_ (_14655_, _14654_, _02445_);
  or _45680_ (_14656_, _14655_, _14651_);
  and _45681_ (_14657_, _14656_, _02459_);
  or _45682_ (_14658_, _14657_, _02458_);
  or _45683_ (_14659_, _14658_, _14647_);
  and _45684_ (_14660_, _14659_, _14637_);
  or _45685_ (_14661_, _14660_, _02398_);
  and _45686_ (_14662_, _14661_, _14615_);
  and _45687_ (_14663_, _14662_, _02400_);
  or _45688_ (_14664_, _14663_, _14568_);
  and _45689_ (_14665_, _14664_, _02405_);
  or _45690_ (_14666_, _14665_, _14474_);
  and _45691_ (_14667_, _14666_, _02444_);
  or _45692_ (_14668_, _14667_, _14283_);
  or _45693_ (_14669_, _14668_, _02443_);
  or _45694_ (_14670_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and _45695_ (_14671_, _14670_, _22762_);
  and _45696_ (_04499_, _14671_, _14669_);
  and _45697_ (_14672_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and _45698_ (_14673_, _13777_, _24050_);
  or _45699_ (_04502_, _14673_, _14672_);
  and _45700_ (_14674_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and _45701_ (_14675_, _02204_, _23898_);
  or _45702_ (_04503_, _14675_, _14674_);
  and _45703_ (_14676_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and _45704_ (_14677_, _13763_, _24050_);
  or _45705_ (_27245_, _14677_, _14676_);
  and _45706_ (_14678_, _02205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and _45707_ (_14679_, _02204_, _23707_);
  or _45708_ (_04512_, _14679_, _14678_);
  and _45709_ (_14680_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and _45710_ (_14681_, _13777_, _23707_);
  or _45711_ (_27090_, _14681_, _14680_);
  and _45712_ (_14682_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and _45713_ (_14683_, _25763_, _23747_);
  or _45714_ (_04530_, _14683_, _14682_);
  and _45715_ (_14684_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  and _45716_ (_14685_, _13769_, _23778_);
  or _45717_ (_04534_, _14685_, _14684_);
  and _45718_ (_14686_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  and _45719_ (_14687_, _13828_, _23649_);
  or _45720_ (_04539_, _14687_, _14686_);
  and _45721_ (_14688_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and _45722_ (_14689_, _25763_, _23707_);
  or _45723_ (_04542_, _14689_, _14688_);
  nor _45724_ (_14690_, t2ex_i, rst);
  and _45725_ (_04546_, _14690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  and _45726_ (_14691_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  and _45727_ (_14692_, _13769_, _23824_);
  or _45728_ (_04548_, _14692_, _14691_);
  and _45729_ (_14693_, _25764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and _45730_ (_14694_, _25763_, _24050_);
  or _45731_ (_04550_, _14694_, _14693_);
  and _45732_ (_14695_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  and _45733_ (_14696_, _13769_, _23649_);
  or _45734_ (_04553_, _14696_, _14695_);
  and _45735_ (_14697_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  and _45736_ (_14698_, _13828_, _23747_);
  or _45737_ (_27011_, _14698_, _14697_);
  and _45738_ (_14699_, _25543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  and _45739_ (_14700_, _25542_, _23898_);
  or _45740_ (_04562_, _14700_, _14699_);
  and _45741_ (_14701_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  and _45742_ (_14702_, _13769_, _24050_);
  or _45743_ (_27092_, _14702_, _14701_);
  and _45744_ (_14703_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  and _45745_ (_14704_, _13828_, _23824_);
  or _45746_ (_04566_, _14704_, _14703_);
  and _45747_ (_14705_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  and _45748_ (_14706_, _25252_, _23649_);
  or _45749_ (_27044_, _14706_, _14705_);
  and _45750_ (_14707_, _13770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  and _45751_ (_14708_, _13769_, _23707_);
  or _45752_ (_04573_, _14708_, _14707_);
  and _45753_ (_14709_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not _45754_ (_14710_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _45755_ (_14711_, _22770_, _14710_);
  or _45756_ (_14712_, _14711_, _14709_);
  and _45757_ (_26882_[15], _14712_, _22762_);
  and _45758_ (_14713_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  and _45759_ (_14714_, _25252_, _23824_);
  or _45760_ (_04577_, _14714_, _14713_);
  and _45761_ (_14715_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  and _45762_ (_14716_, _13818_, _23898_);
  or _45763_ (_04580_, _14716_, _14715_);
  and _45764_ (_14717_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and _45765_ (_14718_, _24767_, _23778_);
  or _45766_ (_04583_, _14718_, _14717_);
  not _45767_ (_14719_, _24174_);
  and _45768_ (_14720_, _14719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _45769_ (_14721_, _24145_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _45770_ (_14722_, _14721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _45771_ (_14723_, _14722_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _45772_ (_14724_, _14723_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _45773_ (_14725_, _24173_, _24178_);
  and _45774_ (_14726_, _14725_, _14724_);
  and _45775_ (_14727_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _45776_ (_14728_, _14727_, _14726_);
  nor _45777_ (_14729_, _14728_, _24127_);
  or _45778_ (_14730_, _14729_, _14720_);
  and _45779_ (_14731_, _14730_, _24166_);
  and _45780_ (_14732_, _24121_, _23738_);
  or _45781_ (_04585_, _14732_, _14731_);
  and _45782_ (_14733_, _25253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  and _45783_ (_14734_, _25252_, _23707_);
  or _45784_ (_04587_, _14734_, _14733_);
  and _45785_ (_14735_, _24121_, _24685_);
  nor _45786_ (_14736_, _24145_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _45787_ (_14737_, _14736_, _14721_);
  and _45788_ (_14738_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _45789_ (_14739_, _14738_, _14737_);
  nand _45790_ (_14740_, _14739_, _24174_);
  or _45791_ (_14741_, _24174_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _45792_ (_14742_, _14741_, _14740_);
  and _45793_ (_14743_, _14742_, _24166_);
  or _45794_ (_04590_, _14743_, _14735_);
  and _45795_ (_14744_, _08799_, _24050_);
  and _45796_ (_14745_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  or _45797_ (_04592_, _14745_, _14744_);
  and _45798_ (_14746_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and _45799_ (_14747_, _24767_, _23707_);
  or _45800_ (_04597_, _14747_, _14746_);
  and _45801_ (_14748_, _24852_, _23778_);
  and _45802_ (_14749_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  or _45803_ (_04610_, _14749_, _14748_);
  nor _45804_ (_26897_[1], _00392_, rst);
  and _45805_ (_14750_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  and _45806_ (_14751_, _13818_, _23824_);
  or _45807_ (_04614_, _14751_, _14750_);
  and _45808_ (_14752_, _24768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and _45809_ (_14753_, _24767_, _23649_);
  or _45810_ (_04617_, _14753_, _14752_);
  and _45811_ (_14754_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  and _45812_ (_14755_, _13818_, _23649_);
  or _45813_ (_04620_, _14755_, _14754_);
  or _45814_ (_14756_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _45815_ (_14757_, _14756_, _22762_);
  or _45816_ (_14758_, _02037_, _23642_);
  and _45817_ (_04622_, _14758_, _14757_);
  and _45818_ (_14759_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand _45819_ (_14760_, _24127_, _23772_);
  nor _45820_ (_14761_, _24159_, _24155_);
  and _45821_ (_14762_, _14761_, _24157_);
  nor _45822_ (_14763_, _14761_, _24157_);
  or _45823_ (_14764_, _14763_, _14762_);
  or _45824_ (_14765_, _14764_, _24127_);
  and _45825_ (_14766_, _14765_, _14760_);
  and _45826_ (_14767_, _14766_, _24166_);
  or _45827_ (_04624_, _14767_, _14759_);
  and _45828_ (_14768_, _24226_, _23824_);
  and _45829_ (_14769_, _24229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  or _45830_ (_04626_, _14769_, _14768_);
  and _45831_ (_14770_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  and _45832_ (_14771_, _13818_, _23946_);
  or _45833_ (_27093_, _14771_, _14770_);
  and _45834_ (_14772_, _24194_, _23824_);
  and _45835_ (_14773_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or _45836_ (_27047_, _14773_, _14772_);
  and _45837_ (_14774_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  and _45838_ (_14775_, _13818_, _24050_);
  or _45839_ (_27094_, _14775_, _14774_);
  and _45840_ (_14776_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and _45841_ (_14777_, _13894_, _23824_);
  or _45842_ (_04635_, _14777_, _14776_);
  and _45843_ (_14778_, _02313_, _23824_);
  and _45844_ (_14779_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or _45845_ (_04638_, _14779_, _14778_);
  and _45846_ (_14780_, _08043_, _23649_);
  and _45847_ (_14781_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or _45848_ (_04640_, _14781_, _14780_);
  and _45849_ (_14782_, _26113_, _26110_);
  nor _45850_ (_14783_, _09920_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _45851_ (_14784_, _14783_, _14782_);
  and _45852_ (_14785_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _45853_ (_14786_, _14785_, _04864_);
  nor _45854_ (_14787_, _14786_, _14784_);
  nor _45855_ (_14788_, _14787_, _24299_);
  and _45856_ (_14789_, _24299_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _45857_ (_14790_, _14789_, _14788_);
  and _45858_ (_14791_, _14790_, _24294_);
  and _45859_ (_14792_, _24293_, _23738_);
  or _45860_ (_14793_, _14792_, _14791_);
  and _45861_ (_04642_, _14793_, _22762_);
  and _45862_ (_14794_, _24194_, _23946_);
  and _45863_ (_14795_, _24196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or _45864_ (_04645_, _14795_, _14794_);
  and _45865_ (_14796_, _02313_, _23898_);
  and _45866_ (_14797_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or _45867_ (_04647_, _14797_, _14796_);
  and _45868_ (_14798_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and _45869_ (_14799_, _13894_, _23898_);
  or _45870_ (_04649_, _14799_, _14798_);
  and _45871_ (_14800_, _24081_, _24050_);
  and _45872_ (_14801_, _24083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or _45873_ (_04651_, _14801_, _14800_);
  and _45874_ (_14802_, _02313_, _23778_);
  and _45875_ (_14803_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or _45876_ (_04653_, _14803_, _14802_);
  and _45877_ (_14804_, _13819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  and _45878_ (_14805_, _13818_, _23707_);
  or _45879_ (_04655_, _14805_, _14804_);
  or _45880_ (_14806_, _04891_, _23816_);
  or _45881_ (_14807_, _04880_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _45882_ (_14808_, _14807_, _26097_);
  nor _45883_ (_14809_, _14808_, _04881_);
  and _45884_ (_14810_, _04864_, _24307_);
  or _45885_ (_14811_, _14810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  not _45886_ (_14812_, _04866_);
  and _45887_ (_14813_, _14812_, _04860_);
  and _45888_ (_14814_, _14813_, _14811_);
  and _45889_ (_14815_, _24307_, _24300_);
  and _45890_ (_14816_, _14815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _45891_ (_14817_, _14816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _45892_ (_14818_, _04874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _45893_ (_14819_, _14818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _45894_ (_14820_, _14819_, _14817_);
  or _45895_ (_14821_, _14820_, _14814_);
  or _45896_ (_14822_, _14821_, _14809_);
  or _45897_ (_14823_, _14822_, _24299_);
  and _45898_ (_14824_, _14823_, _24294_);
  and _45899_ (_14825_, _14824_, _14806_);
  and _45900_ (_14826_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _45901_ (_14827_, _14826_, _14825_);
  and _45902_ (_04657_, _14827_, _22762_);
  or _45903_ (_14828_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _45904_ (_14829_, _14828_, _22762_);
  or _45905_ (_14830_, _24079_, _23816_);
  and _45906_ (_04659_, _14830_, _14829_);
  and _45907_ (_14831_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and _45908_ (_14832_, _13894_, _23778_);
  or _45909_ (_04662_, _14832_, _14831_);
  and _45910_ (_14833_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  and _45911_ (_14834_, _13752_, _23747_);
  or _45912_ (_04664_, _14834_, _14833_);
  and _45913_ (_14835_, _23898_, _23755_);
  and _45914_ (_14836_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  or _45915_ (_04670_, _14836_, _14835_);
  and _45916_ (_14837_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  and _45917_ (_14838_, _13752_, _23649_);
  or _45918_ (_04672_, _14838_, _14837_);
  and _45919_ (_14839_, _08799_, _23946_);
  and _45920_ (_14840_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or _45921_ (_04687_, _14840_, _14839_);
  and _45922_ (_14841_, _23833_, _23707_);
  and _45923_ (_14842_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or _45924_ (_04689_, _14842_, _14841_);
  and _45925_ (_14843_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  and _45926_ (_14844_, _13752_, _24050_);
  or _45927_ (_04692_, _14844_, _14843_);
  and _45928_ (_14845_, _02313_, _23707_);
  and _45929_ (_14846_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or _45930_ (_04697_, _14846_, _14845_);
  and _45931_ (_14847_, _02200_, _23747_);
  and _45932_ (_14848_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or _45933_ (_04699_, _14848_, _14847_);
  and _45934_ (_14849_, _02200_, _23946_);
  and _45935_ (_14850_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or _45936_ (_27167_, _14850_, _14849_);
  and _45937_ (_14851_, _24331_, _23747_);
  and _45938_ (_14852_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or _45939_ (_04710_, _14852_, _14851_);
  and _45940_ (_14853_, _13753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  and _45941_ (_14854_, _13752_, _23707_);
  or _45942_ (_04713_, _14854_, _14853_);
  or _45943_ (_14855_, _24464_, _23837_);
  or _45944_ (_14856_, _22767_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _45945_ (_14857_, _14856_, _22762_);
  and _45946_ (_26864_[4], _14857_, _14855_);
  and _45947_ (_14858_, _02313_, _23946_);
  and _45948_ (_14859_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or _45949_ (_04716_, _14859_, _14858_);
  and _45950_ (_14860_, _24331_, _23898_);
  and _45951_ (_14861_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or _45952_ (_04719_, _14861_, _14860_);
  and _45953_ (_14862_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and _45954_ (_14863_, _12980_, _23898_);
  or _45955_ (_04722_, _14863_, _14862_);
  and _45956_ (_14864_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and _45957_ (_14865_, _12980_, _23824_);
  or _45958_ (_04731_, _14865_, _14864_);
  and _45959_ (_14866_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or _45960_ (_04733_, _14866_, _05664_);
  and _45961_ (_14867_, _05350_, _23946_);
  and _45962_ (_14868_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  or _45963_ (_27065_, _14868_, _14867_);
  and _45964_ (_14869_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and _45965_ (_14870_, _13894_, _23946_);
  or _45966_ (_04739_, _14870_, _14869_);
  and _45967_ (_14871_, _02313_, _23747_);
  and _45968_ (_14872_, _02315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or _45969_ (_27156_, _14872_, _14871_);
  and _45970_ (_14873_, _04811_, _24050_);
  and _45971_ (_14874_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  or _45972_ (_04747_, _14874_, _14873_);
  and _45973_ (_14875_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and _45974_ (_14876_, _12980_, _23747_);
  or _45975_ (_04750_, _14876_, _14875_);
  and _45976_ (_14877_, _04811_, _23649_);
  and _45977_ (_14878_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  or _45978_ (_04753_, _14878_, _14877_);
  and _45979_ (_14879_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and _45980_ (_14880_, _12980_, _23946_);
  or _45981_ (_04755_, _14880_, _14879_);
  and _45982_ (_14881_, _05281_, _23649_);
  and _45983_ (_14882_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or _45984_ (_04759_, _14882_, _14881_);
  and _45985_ (_14883_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and _45986_ (_14884_, _13894_, _23649_);
  or _45987_ (_04765_, _14884_, _14883_);
  and _45988_ (_14885_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and _45989_ (_14886_, _13894_, _23747_);
  or _45990_ (_04777_, _14886_, _14885_);
  and _45991_ (_14887_, _12981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and _45992_ (_14888_, _12980_, _23707_);
  or _45993_ (_27095_, _14888_, _14887_);
  and _45994_ (_14889_, _02321_, _23824_);
  and _45995_ (_14890_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  or _45996_ (_04779_, _14890_, _14889_);
  and _45997_ (_14891_, _02321_, _23747_);
  and _45998_ (_14892_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  or _45999_ (_27139_, _14892_, _14891_);
  and _46000_ (_14893_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and _46001_ (_14894_, _12974_, _23778_);
  or _46002_ (_04784_, _14894_, _14893_);
  and _46003_ (_14895_, _02370_, _23707_);
  and _46004_ (_14896_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or _46005_ (_27067_, _14896_, _14895_);
  and _46006_ (_14897_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and _46007_ (_14898_, _12974_, _23824_);
  or _46008_ (_04796_, _14898_, _14897_);
  and _46009_ (_14899_, _04922_, _23824_);
  and _46010_ (_14900_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  or _46011_ (_04798_, _14900_, _14899_);
  and _46012_ (_14901_, _25739_, _23707_);
  and _46013_ (_14902_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or _46014_ (_04803_, _14902_, _14901_);
  and _46015_ (_14903_, _06886_, _23656_);
  not _46016_ (_14904_, _14903_);
  and _46017_ (_14905_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  and _46018_ (_14906_, _14903_, _23747_);
  or _46019_ (_04808_, _14906_, _14905_);
  and _46020_ (_14907_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  and _46021_ (_14908_, _14903_, _23824_);
  or _46022_ (_04815_, _14908_, _14907_);
  and _46023_ (_14909_, _02321_, _23946_);
  and _46024_ (_14910_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  or _46025_ (_04818_, _14910_, _14909_);
  and _46026_ (_14911_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and _46027_ (_14912_, _12974_, _23747_);
  or _46028_ (_04824_, _14912_, _14911_);
  and _46029_ (_14913_, _04922_, _24050_);
  and _46030_ (_14914_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  or _46031_ (_04827_, _14914_, _14913_);
  and _46032_ (_14915_, _02321_, _23707_);
  and _46033_ (_14916_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  or _46034_ (_27140_, _14916_, _14915_);
  and _46035_ (_14917_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and _46036_ (_14918_, _12974_, _24050_);
  or _46037_ (_04837_, _14918_, _14917_);
  and _46038_ (_14919_, _25748_, _23778_);
  and _46039_ (_14920_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or _46040_ (_04841_, _14920_, _14919_);
  and _46041_ (_14921_, _09913_, _24050_);
  and _46042_ (_14922_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or _46043_ (_04844_, _14922_, _14921_);
  and _46044_ (_14923_, _02321_, _24050_);
  and _46045_ (_14924_, _02323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  or _46046_ (_04847_, _14924_, _14923_);
  and _46047_ (_14925_, _24852_, _23946_);
  and _46048_ (_14926_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  or _46049_ (_04849_, _14926_, _14925_);
  and _46050_ (_14927_, _25748_, _23946_);
  and _46051_ (_14928_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or _46052_ (_04865_, _14928_, _14927_);
  and _46053_ (_14929_, _12975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and _46054_ (_14930_, _12974_, _23707_);
  or _46055_ (_04868_, _14930_, _14929_);
  and _46056_ (_14931_, _25748_, _23747_);
  and _46057_ (_14932_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or _46058_ (_04870_, _14932_, _14931_);
  and _46059_ (_14933_, _07743_, _23824_);
  and _46060_ (_14934_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  or _46061_ (_04875_, _14934_, _14933_);
  and _46062_ (_14935_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  and _46063_ (_14936_, _12970_, _23778_);
  or _46064_ (_27097_, _14936_, _14935_);
  and _46065_ (_14937_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  and _46066_ (_14939_, _14903_, _23649_);
  or _46067_ (_04884_, _14939_, _14937_);
  and _46068_ (_14940_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  and _46069_ (_14941_, _12970_, _23824_);
  or _46070_ (_04889_, _14941_, _14940_);
  and _46071_ (_14942_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  and _46072_ (_14943_, _14903_, _24050_);
  or _46073_ (_04893_, _14943_, _14942_);
  and _46074_ (_14944_, _24639_, _23898_);
  and _46075_ (_14945_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or _46076_ (_04899_, _14945_, _14944_);
  and _46077_ (_14946_, _05350_, _23778_);
  and _46078_ (_14947_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  or _46079_ (_04902_, _14947_, _14946_);
  and _46080_ (_14948_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  and _46081_ (_14949_, _14903_, _23946_);
  or _46082_ (_04904_, _14949_, _14948_);
  and _46083_ (_14950_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  and _46084_ (_14951_, _12970_, _23649_);
  or _46085_ (_04906_, _14951_, _14950_);
  and _46086_ (_14952_, _02200_, _24050_);
  and _46087_ (_14953_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or _46088_ (_04910_, _14953_, _14952_);
  and _46089_ (_14954_, _09913_, _23649_);
  and _46090_ (_14955_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or _46091_ (_04912_, _14955_, _14954_);
  and _46092_ (_14956_, _23911_, _23664_);
  and _46093_ (_14957_, _14956_, _23649_);
  not _46094_ (_14958_, _14956_);
  and _46095_ (_14959_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or _46096_ (_04916_, _14959_, _14957_);
  and _46097_ (_14960_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  and _46098_ (_14961_, _12970_, _23946_);
  or _46099_ (_04921_, _14961_, _14960_);
  and _46100_ (_14962_, _12971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  and _46101_ (_14963_, _12970_, _23707_);
  or _46102_ (_04923_, _14963_, _14962_);
  and _46103_ (_14964_, _24639_, _23946_);
  and _46104_ (_14965_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or _46105_ (_27169_, _14965_, _14964_);
  and _46106_ (_14966_, _14956_, _23707_);
  and _46107_ (_14967_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or _46108_ (_04930_, _14967_, _14966_);
  and _46109_ (_14968_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  and _46110_ (_14969_, _12941_, _23778_);
  or _46111_ (_04932_, _14969_, _14968_);
  and _46112_ (_14970_, _24639_, _23824_);
  and _46113_ (_14971_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or _46114_ (_04933_, _14971_, _14970_);
  and _46115_ (_14972_, _12782_, _23946_);
  and _46116_ (_14973_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or _46117_ (_04951_, _14973_, _14972_);
  and _46118_ (_14974_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  and _46119_ (_14975_, _12941_, _23824_);
  or _46120_ (_04954_, _14975_, _14974_);
  and _46121_ (_14976_, _24639_, _23747_);
  and _46122_ (_14977_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or _46123_ (_04960_, _14977_, _14976_);
  and _46124_ (_14978_, _08799_, _23649_);
  and _46125_ (_14979_, _08801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  or _46126_ (_04963_, _14979_, _14978_);
  and _46127_ (_14980_, _23946_, _23665_);
  and _46128_ (_14981_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or _46129_ (_04971_, _14981_, _14980_);
  and _46130_ (_14982_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  and _46131_ (_14983_, _12941_, _23747_);
  or _46132_ (_27101_, _14983_, _14982_);
  and _46133_ (_14984_, _23824_, _23665_);
  and _46134_ (_14985_, _23709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  or _46135_ (_04975_, _14985_, _14984_);
  and _46136_ (_14986_, _02107_, _23747_);
  and _46137_ (_14987_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  or _46138_ (_04986_, _14987_, _14986_);
  and _46139_ (_14988_, _03300_, _23649_);
  and _46140_ (_14989_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or _46141_ (_04988_, _14989_, _14988_);
  and _46142_ (_14990_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  and _46143_ (_14991_, _12941_, _23946_);
  or _46144_ (_04990_, _14991_, _14990_);
  and _46145_ (_14992_, _12942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  and _46146_ (_14993_, _12941_, _23707_);
  or _46147_ (_04997_, _14993_, _14992_);
  and _46148_ (_14994_, _02107_, _23824_);
  and _46149_ (_14995_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  or _46150_ (_04999_, _14995_, _14994_);
  and _46151_ (_14996_, _06886_, _25078_);
  not _46152_ (_14997_, _14996_);
  and _46153_ (_14998_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  and _46154_ (_14999_, _14996_, _23946_);
  or _46155_ (_05002_, _14999_, _14998_);
  and _46156_ (_15000_, _01971_, _23747_);
  and _46157_ (_15001_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  or _46158_ (_05004_, _15001_, _15000_);
  and _46159_ (_15002_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and _46160_ (_15003_, _12935_, _23898_);
  or _46161_ (_05010_, _15003_, _15002_);
  and _46162_ (_15004_, _01808_, _23664_);
  and _46163_ (_15005_, _15004_, _23824_);
  not _46164_ (_15006_, _15004_);
  and _46165_ (_15007_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or _46166_ (_05015_, _15007_, _15005_);
  and _46167_ (_15008_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  and _46168_ (_15009_, _14996_, _23649_);
  or _46169_ (_05021_, _15009_, _15008_);
  and _46170_ (_15010_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  and _46171_ (_15011_, _14996_, _23747_);
  or _46172_ (_05040_, _15011_, _15010_);
  and _46173_ (_15012_, _23664_, _23069_);
  and _46174_ (_15013_, _15012_, _23778_);
  not _46175_ (_15014_, _15012_);
  and _46176_ (_15015_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or _46177_ (_05043_, _15015_, _15013_);
  and _46178_ (_15016_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and _46179_ (_15017_, _12935_, _23824_);
  or _46180_ (_05046_, _15017_, _15016_);
  and _46181_ (_15018_, _02107_, _23707_);
  and _46182_ (_15019_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  or _46183_ (_05048_, _15019_, _15018_);
  and _46184_ (_15020_, _15004_, _24050_);
  and _46185_ (_15021_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or _46186_ (_05051_, _15021_, _15020_);
  and _46187_ (_15022_, _15012_, _23946_);
  and _46188_ (_15023_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or _46189_ (_05056_, _15023_, _15022_);
  and _46190_ (_15024_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and _46191_ (_15025_, _12935_, _23747_);
  or _46192_ (_05059_, _15025_, _15024_);
  and _46193_ (_15026_, _15012_, _23824_);
  and _46194_ (_15027_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or _46195_ (_05062_, _15027_, _15026_);
  and _46196_ (_15028_, _02107_, _24050_);
  and _46197_ (_15029_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  or _46198_ (_05069_, _15029_, _15028_);
  and _46199_ (_15030_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and _46200_ (_15031_, _12935_, _23946_);
  or _46201_ (_05071_, _15031_, _15030_);
  and _46202_ (_15032_, _12733_, _23898_);
  and _46203_ (_15033_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  or _46204_ (_05076_, _15033_, _15032_);
  and _46205_ (_15034_, _12936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and _46206_ (_15035_, _12935_, _23707_);
  or _46207_ (_05078_, _15035_, _15034_);
  and _46208_ (_15036_, _05042_, _23898_);
  and _46209_ (_15037_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or _46210_ (_27134_, _15037_, _15036_);
  and _46211_ (_15038_, _02107_, _23946_);
  and _46212_ (_15039_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  or _46213_ (_05082_, _15039_, _15038_);
  and _46214_ (_15040_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and _46215_ (_15041_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or _46216_ (_15042_, _15041_, _15040_);
  and _46217_ (_15043_, _15042_, _02393_);
  and _46218_ (_15044_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and _46219_ (_15045_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or _46220_ (_15046_, _15045_, _15044_);
  and _46221_ (_15047_, _15046_, _02445_);
  or _46222_ (_15048_, _15047_, _15043_);
  and _46223_ (_15049_, _15048_, _02421_);
  and _46224_ (_15050_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and _46225_ (_15051_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or _46226_ (_15052_, _15051_, _15050_);
  and _46227_ (_15053_, _15052_, _02393_);
  and _46228_ (_15054_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and _46229_ (_15055_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or _46230_ (_15056_, _15055_, _15054_);
  and _46231_ (_15057_, _15056_, _02445_);
  or _46232_ (_15058_, _15057_, _15053_);
  and _46233_ (_15059_, _15058_, _02459_);
  or _46234_ (_15060_, _15059_, _15049_);
  and _46235_ (_15061_, _15060_, _02458_);
  or _46236_ (_15062_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or _46237_ (_15063_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and _46238_ (_15064_, _15063_, _15062_);
  and _46239_ (_15065_, _15064_, _02393_);
  or _46240_ (_15066_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or _46241_ (_15067_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and _46242_ (_15068_, _15067_, _15066_);
  and _46243_ (_15069_, _15068_, _02445_);
  or _46244_ (_15070_, _15069_, _15065_);
  and _46245_ (_15071_, _15070_, _02421_);
  or _46246_ (_15072_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or _46247_ (_15073_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and _46248_ (_15074_, _15073_, _15072_);
  and _46249_ (_15075_, _15074_, _02393_);
  or _46250_ (_15076_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or _46251_ (_15077_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and _46252_ (_15078_, _15077_, _15076_);
  and _46253_ (_15079_, _15078_, _02445_);
  or _46254_ (_15080_, _15079_, _15075_);
  and _46255_ (_15081_, _15080_, _02459_);
  or _46256_ (_15082_, _15081_, _15071_);
  and _46257_ (_15083_, _15082_, _02414_);
  or _46258_ (_15084_, _15083_, _15061_);
  and _46259_ (_15085_, _15084_, _02398_);
  and _46260_ (_15086_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and _46261_ (_15087_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or _46262_ (_15088_, _15087_, _15086_);
  and _46263_ (_15089_, _15088_, _02393_);
  and _46264_ (_15090_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and _46265_ (_15091_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or _46266_ (_15092_, _15091_, _15090_);
  and _46267_ (_15093_, _15092_, _02445_);
  or _46268_ (_15094_, _15093_, _15089_);
  and _46269_ (_15095_, _15094_, _02421_);
  and _46270_ (_15096_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and _46271_ (_15097_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or _46272_ (_15098_, _15097_, _15096_);
  and _46273_ (_15099_, _15098_, _02393_);
  and _46274_ (_15100_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and _46275_ (_15101_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or _46276_ (_15102_, _15101_, _15100_);
  and _46277_ (_15103_, _15102_, _02445_);
  or _46278_ (_15104_, _15103_, _15099_);
  and _46279_ (_15105_, _15104_, _02459_);
  or _46280_ (_15106_, _15105_, _15095_);
  and _46281_ (_15107_, _15106_, _02458_);
  or _46282_ (_15108_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or _46283_ (_15109_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and _46284_ (_15110_, _15109_, _02445_);
  and _46285_ (_15111_, _15110_, _15108_);
  or _46286_ (_15112_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or _46287_ (_15113_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and _46288_ (_15114_, _15113_, _02393_);
  and _46289_ (_15115_, _15114_, _15112_);
  or _46290_ (_15116_, _15115_, _15111_);
  and _46291_ (_15117_, _15116_, _02421_);
  or _46292_ (_15118_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or _46293_ (_15119_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and _46294_ (_15120_, _15119_, _02445_);
  and _46295_ (_15121_, _15120_, _15118_);
  or _46296_ (_15122_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or _46297_ (_15123_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and _46298_ (_15124_, _15123_, _02393_);
  and _46299_ (_15125_, _15124_, _15122_);
  or _46300_ (_15126_, _15125_, _15121_);
  and _46301_ (_15127_, _15126_, _02459_);
  or _46302_ (_15128_, _15127_, _15117_);
  and _46303_ (_15129_, _15128_, _02414_);
  or _46304_ (_15130_, _15129_, _15107_);
  and _46305_ (_15131_, _15130_, _02496_);
  or _46306_ (_15133_, _15131_, _15085_);
  and _46307_ (_15134_, _15133_, _02400_);
  and _46308_ (_15135_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and _46309_ (_15136_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or _46310_ (_15137_, _15136_, _15135_);
  and _46311_ (_15138_, _15137_, _02393_);
  and _46312_ (_15139_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and _46313_ (_15140_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or _46314_ (_15141_, _15140_, _15139_);
  and _46315_ (_15142_, _15141_, _02445_);
  or _46316_ (_15143_, _15142_, _15138_);
  or _46317_ (_15144_, _15143_, _02459_);
  and _46318_ (_15145_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and _46319_ (_15146_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or _46320_ (_15147_, _15146_, _15145_);
  and _46321_ (_15148_, _15147_, _02393_);
  and _46322_ (_15149_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and _46323_ (_15150_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or _46324_ (_15151_, _15150_, _15149_);
  and _46325_ (_15152_, _15151_, _02445_);
  or _46326_ (_15154_, _15152_, _15148_);
  or _46327_ (_15155_, _15154_, _02421_);
  and _46328_ (_15156_, _15155_, _02458_);
  and _46329_ (_15157_, _15156_, _15144_);
  or _46330_ (_15158_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or _46331_ (_15159_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and _46332_ (_15160_, _15159_, _02445_);
  and _46333_ (_15161_, _15160_, _15158_);
  or _46334_ (_15162_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or _46335_ (_15163_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and _46336_ (_15164_, _15163_, _02393_);
  and _46337_ (_15165_, _15164_, _15162_);
  or _46338_ (_15166_, _15165_, _15161_);
  or _46339_ (_15167_, _15166_, _02459_);
  or _46340_ (_15168_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or _46341_ (_15169_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and _46342_ (_15170_, _15169_, _02445_);
  and _46343_ (_15171_, _15170_, _15168_);
  or _46344_ (_15172_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or _46345_ (_15173_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and _46346_ (_15174_, _15173_, _02393_);
  and _46347_ (_15175_, _15174_, _15172_);
  or _46348_ (_15176_, _15175_, _15171_);
  or _46349_ (_15177_, _15176_, _02421_);
  and _46350_ (_15178_, _15177_, _02414_);
  and _46351_ (_15179_, _15178_, _15167_);
  or _46352_ (_15180_, _15179_, _15157_);
  and _46353_ (_15181_, _15180_, _02496_);
  and _46354_ (_15182_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and _46355_ (_15183_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or _46356_ (_15184_, _15183_, _15182_);
  and _46357_ (_15185_, _15184_, _02393_);
  and _46358_ (_15186_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and _46359_ (_15187_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or _46360_ (_15188_, _15187_, _15186_);
  and _46361_ (_15189_, _15188_, _02445_);
  or _46362_ (_15190_, _15189_, _15185_);
  or _46363_ (_15191_, _15190_, _02459_);
  and _46364_ (_15192_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and _46365_ (_15193_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or _46366_ (_15194_, _15193_, _15192_);
  and _46367_ (_15195_, _15194_, _02393_);
  and _46368_ (_15196_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and _46369_ (_15197_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or _46370_ (_15198_, _15197_, _15196_);
  and _46371_ (_15199_, _15198_, _02445_);
  or _46372_ (_15200_, _15199_, _15195_);
  or _46373_ (_15201_, _15200_, _02421_);
  and _46374_ (_15202_, _15201_, _02458_);
  and _46375_ (_15203_, _15202_, _15191_);
  or _46376_ (_15204_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or _46377_ (_15205_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and _46378_ (_15206_, _15205_, _15204_);
  and _46379_ (_15207_, _15206_, _02393_);
  or _46380_ (_15208_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or _46381_ (_15209_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and _46382_ (_15210_, _15209_, _15208_);
  and _46383_ (_15211_, _15210_, _02445_);
  or _46384_ (_15212_, _15211_, _15207_);
  or _46385_ (_15213_, _15212_, _02459_);
  or _46386_ (_15214_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or _46387_ (_15215_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and _46388_ (_15216_, _15215_, _15214_);
  and _46389_ (_15217_, _15216_, _02393_);
  or _46390_ (_15218_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or _46391_ (_15219_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and _46392_ (_15220_, _15219_, _15218_);
  and _46393_ (_15221_, _15220_, _02445_);
  or _46394_ (_15222_, _15221_, _15217_);
  or _46395_ (_15223_, _15222_, _02421_);
  and _46396_ (_15224_, _15223_, _02414_);
  and _46397_ (_15225_, _15224_, _15213_);
  or _46398_ (_15226_, _15225_, _15203_);
  and _46399_ (_15227_, _15226_, _02398_);
  or _46400_ (_15228_, _15227_, _15181_);
  and _46401_ (_15229_, _15228_, _02546_);
  or _46402_ (_15230_, _15229_, _15134_);
  and _46403_ (_15231_, _15230_, _02646_);
  and _46404_ (_15232_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and _46405_ (_15233_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or _46406_ (_15234_, _15233_, _15232_);
  and _46407_ (_15235_, _15234_, _02445_);
  and _46408_ (_15236_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and _46409_ (_15237_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or _46410_ (_15238_, _15237_, _15236_);
  and _46411_ (_15239_, _15238_, _02393_);
  or _46412_ (_15240_, _15239_, _15235_);
  or _46413_ (_15241_, _15240_, _02459_);
  and _46414_ (_15242_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and _46415_ (_15243_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or _46416_ (_15244_, _15243_, _15242_);
  and _46417_ (_15245_, _15244_, _02445_);
  and _46418_ (_15246_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and _46419_ (_15247_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or _46420_ (_15248_, _15247_, _15246_);
  and _46421_ (_15249_, _15248_, _02393_);
  or _46422_ (_15250_, _15249_, _15245_);
  or _46423_ (_15251_, _15250_, _02421_);
  and _46424_ (_15252_, _15251_, _02458_);
  and _46425_ (_15253_, _15252_, _15241_);
  or _46426_ (_15254_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or _46427_ (_15255_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and _46428_ (_15256_, _15255_, _02393_);
  and _46429_ (_15257_, _15256_, _15254_);
  or _46430_ (_15258_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or _46431_ (_15259_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and _46432_ (_15260_, _15259_, _02445_);
  and _46433_ (_15261_, _15260_, _15258_);
  or _46434_ (_15262_, _15261_, _15257_);
  or _46435_ (_15263_, _15262_, _02459_);
  or _46436_ (_15264_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or _46437_ (_15265_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and _46438_ (_15266_, _15265_, _02393_);
  and _46439_ (_15267_, _15266_, _15264_);
  or _46440_ (_15268_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or _46441_ (_15269_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and _46442_ (_15270_, _15269_, _02445_);
  and _46443_ (_15271_, _15270_, _15268_);
  or _46444_ (_15272_, _15271_, _15267_);
  or _46445_ (_15273_, _15272_, _02421_);
  and _46446_ (_15274_, _15273_, _02414_);
  and _46447_ (_15275_, _15274_, _15263_);
  or _46448_ (_15276_, _15275_, _15253_);
  or _46449_ (_15277_, _15276_, _02398_);
  and _46450_ (_15278_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and _46451_ (_15279_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or _46452_ (_15280_, _15279_, _02393_);
  or _46453_ (_15281_, _15280_, _15278_);
  and _46454_ (_15282_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and _46455_ (_15283_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or _46456_ (_15284_, _15283_, _02445_);
  or _46457_ (_15285_, _15284_, _15282_);
  and _46458_ (_15286_, _15285_, _15281_);
  or _46459_ (_15287_, _15286_, _02459_);
  and _46460_ (_15288_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and _46461_ (_15289_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or _46462_ (_15290_, _15289_, _02393_);
  or _46463_ (_15291_, _15290_, _15288_);
  and _46464_ (_15292_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and _46465_ (_15293_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or _46466_ (_15294_, _15293_, _02445_);
  or _46467_ (_15295_, _15294_, _15292_);
  and _46468_ (_15296_, _15295_, _15291_);
  or _46469_ (_15297_, _15296_, _02421_);
  and _46470_ (_15298_, _15297_, _02458_);
  and _46471_ (_15299_, _15298_, _15287_);
  or _46472_ (_15300_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or _46473_ (_15301_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and _46474_ (_15302_, _15301_, _15300_);
  or _46475_ (_15303_, _15302_, _02445_);
  or _46476_ (_15304_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or _46477_ (_15305_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and _46478_ (_15306_, _15305_, _15304_);
  or _46479_ (_15307_, _15306_, _02393_);
  and _46480_ (_15308_, _15307_, _15303_);
  or _46481_ (_15309_, _15308_, _02459_);
  or _46482_ (_15310_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or _46483_ (_15311_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and _46484_ (_15312_, _15311_, _15310_);
  or _46485_ (_15313_, _15312_, _02445_);
  or _46486_ (_15314_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or _46487_ (_15315_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and _46488_ (_15316_, _15315_, _15314_);
  or _46489_ (_15317_, _15316_, _02393_);
  and _46490_ (_15318_, _15317_, _15313_);
  or _46491_ (_15319_, _15318_, _02421_);
  and _46492_ (_15320_, _15319_, _02414_);
  and _46493_ (_15321_, _15320_, _15309_);
  or _46494_ (_15322_, _15321_, _15299_);
  or _46495_ (_15323_, _15322_, _02496_);
  and _46496_ (_15324_, _15323_, _02546_);
  and _46497_ (_15325_, _15324_, _15277_);
  and _46498_ (_15326_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  and _46499_ (_15327_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  or _46500_ (_15328_, _15327_, _15326_);
  and _46501_ (_15329_, _15328_, _02393_);
  and _46502_ (_15330_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  and _46503_ (_15331_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or _46504_ (_15332_, _15331_, _15330_);
  and _46505_ (_15333_, _15332_, _02445_);
  or _46506_ (_15334_, _15333_, _15329_);
  and _46507_ (_15335_, _15334_, _02421_);
  and _46508_ (_15336_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  and _46509_ (_15337_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  or _46510_ (_15338_, _15337_, _15336_);
  and _46511_ (_15339_, _15338_, _02393_);
  and _46512_ (_15340_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  and _46513_ (_15341_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or _46514_ (_15342_, _15341_, _15340_);
  and _46515_ (_15343_, _15342_, _02445_);
  or _46516_ (_15344_, _15343_, _15339_);
  and _46517_ (_15345_, _15344_, _02459_);
  or _46518_ (_15346_, _15345_, _15335_);
  and _46519_ (_15347_, _15346_, _02458_);
  or _46520_ (_15348_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or _46521_ (_15349_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  and _46522_ (_15350_, _15349_, _15348_);
  and _46523_ (_15351_, _15350_, _02393_);
  or _46524_ (_15352_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  or _46525_ (_15353_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  and _46526_ (_15354_, _15353_, _15352_);
  and _46527_ (_15355_, _15354_, _02445_);
  or _46528_ (_15356_, _15355_, _15351_);
  and _46529_ (_15357_, _15356_, _02421_);
  or _46530_ (_15358_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or _46531_ (_15359_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  and _46532_ (_15360_, _15359_, _15358_);
  and _46533_ (_15361_, _15360_, _02393_);
  or _46534_ (_15362_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or _46535_ (_15363_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  and _46536_ (_15364_, _15363_, _15362_);
  and _46537_ (_15365_, _15364_, _02445_);
  or _46538_ (_15366_, _15365_, _15361_);
  and _46539_ (_15367_, _15366_, _02459_);
  or _46540_ (_15368_, _15367_, _15357_);
  and _46541_ (_15369_, _15368_, _02414_);
  or _46542_ (_15370_, _15369_, _15347_);
  and _46543_ (_15371_, _15370_, _02496_);
  and _46544_ (_15372_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and _46545_ (_15373_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or _46546_ (_15374_, _15373_, _15372_);
  and _46547_ (_15375_, _15374_, _02393_);
  and _46548_ (_15376_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and _46549_ (_15377_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or _46550_ (_15378_, _15377_, _15376_);
  and _46551_ (_15379_, _15378_, _02445_);
  or _46552_ (_15380_, _15379_, _15375_);
  and _46553_ (_15381_, _15380_, _02421_);
  and _46554_ (_15382_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and _46555_ (_15383_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or _46556_ (_15384_, _15383_, _15382_);
  and _46557_ (_15385_, _15384_, _02393_);
  and _46558_ (_15386_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and _46559_ (_15387_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or _46560_ (_15388_, _15387_, _15386_);
  and _46561_ (_15389_, _15388_, _02445_);
  or _46562_ (_15390_, _15389_, _15385_);
  and _46563_ (_15391_, _15390_, _02459_);
  or _46564_ (_15392_, _15391_, _15381_);
  and _46565_ (_15393_, _15392_, _02458_);
  or _46566_ (_15394_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or _46567_ (_15395_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and _46568_ (_15396_, _15395_, _15394_);
  and _46569_ (_15397_, _15396_, _02393_);
  or _46570_ (_15398_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or _46571_ (_15399_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and _46572_ (_15400_, _15399_, _15398_);
  and _46573_ (_15401_, _15400_, _02445_);
  or _46574_ (_15402_, _15401_, _15397_);
  and _46575_ (_15403_, _15402_, _02421_);
  or _46576_ (_15404_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or _46577_ (_15405_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and _46578_ (_15406_, _15405_, _15404_);
  and _46579_ (_15407_, _15406_, _02393_);
  or _46580_ (_15408_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or _46581_ (_15409_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and _46582_ (_15410_, _15409_, _15408_);
  and _46583_ (_15411_, _15410_, _02445_);
  or _46584_ (_15412_, _15411_, _15407_);
  and _46585_ (_15413_, _15412_, _02459_);
  or _46586_ (_15414_, _15413_, _15403_);
  and _46587_ (_15415_, _15414_, _02414_);
  or _46588_ (_15416_, _15415_, _15393_);
  and _46589_ (_15417_, _15416_, _02398_);
  or _46590_ (_15418_, _15417_, _15371_);
  and _46591_ (_15419_, _15418_, _02400_);
  or _46592_ (_15420_, _15419_, _15325_);
  and _46593_ (_15421_, _15420_, _02405_);
  or _46594_ (_15422_, _15421_, _15231_);
  and _46595_ (_15423_, _15422_, _26777_);
  and _46596_ (_15424_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  and _46597_ (_15425_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or _46598_ (_15426_, _15425_, _15424_);
  and _46599_ (_15427_, _15426_, _02445_);
  and _46600_ (_15428_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and _46601_ (_15429_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or _46602_ (_15430_, _15429_, _15428_);
  and _46603_ (_15431_, _15430_, _02393_);
  or _46604_ (_15432_, _15431_, _15427_);
  or _46605_ (_15433_, _15432_, _02459_);
  and _46606_ (_15434_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  and _46607_ (_15435_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or _46608_ (_15436_, _15435_, _15434_);
  and _46609_ (_15437_, _15436_, _02445_);
  and _46610_ (_15438_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and _46611_ (_15439_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or _46612_ (_15440_, _15439_, _15438_);
  and _46613_ (_15441_, _15440_, _02393_);
  or _46614_ (_15442_, _15441_, _15437_);
  or _46615_ (_15443_, _15442_, _02421_);
  and _46616_ (_15444_, _15443_, _02458_);
  and _46617_ (_15445_, _15444_, _15433_);
  or _46618_ (_15446_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or _46619_ (_15447_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and _46620_ (_15448_, _15447_, _02393_);
  and _46621_ (_15449_, _15448_, _15446_);
  or _46622_ (_15450_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or _46623_ (_15451_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  and _46624_ (_15452_, _15451_, _02445_);
  and _46625_ (_15453_, _15452_, _15450_);
  or _46626_ (_15454_, _15453_, _15449_);
  or _46627_ (_15455_, _15454_, _02459_);
  or _46628_ (_15456_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or _46629_ (_15457_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and _46630_ (_15458_, _15457_, _02393_);
  and _46631_ (_15459_, _15458_, _15456_);
  or _46632_ (_15460_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or _46633_ (_15461_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and _46634_ (_15462_, _15461_, _02445_);
  and _46635_ (_15463_, _15462_, _15460_);
  or _46636_ (_15464_, _15463_, _15459_);
  or _46637_ (_15465_, _15464_, _02421_);
  and _46638_ (_15466_, _15465_, _02414_);
  and _46639_ (_15467_, _15466_, _15455_);
  or _46640_ (_15468_, _15467_, _15445_);
  and _46641_ (_15469_, _15468_, _02496_);
  and _46642_ (_15470_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  and _46643_ (_15471_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or _46644_ (_15472_, _15471_, _02393_);
  or _46645_ (_15473_, _15472_, _15470_);
  and _46646_ (_15474_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and _46647_ (_15475_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or _46648_ (_15476_, _15475_, _02445_);
  or _46649_ (_15477_, _15476_, _15474_);
  and _46650_ (_15478_, _15477_, _15473_);
  or _46651_ (_15479_, _15478_, _02459_);
  and _46652_ (_15480_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and _46653_ (_15481_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or _46654_ (_15482_, _15481_, _02393_);
  or _46655_ (_15483_, _15482_, _15480_);
  and _46656_ (_15484_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and _46657_ (_15485_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or _46658_ (_15486_, _15485_, _02445_);
  or _46659_ (_15487_, _15486_, _15484_);
  and _46660_ (_15488_, _15487_, _15483_);
  or _46661_ (_15489_, _15488_, _02421_);
  and _46662_ (_15490_, _15489_, _02458_);
  and _46663_ (_15491_, _15490_, _15479_);
  or _46664_ (_15492_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or _46665_ (_15493_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  and _46666_ (_15494_, _15493_, _15492_);
  or _46667_ (_15495_, _15494_, _02445_);
  or _46668_ (_15496_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or _46669_ (_15497_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and _46670_ (_15498_, _15497_, _15496_);
  or _46671_ (_15499_, _15498_, _02393_);
  and _46672_ (_15500_, _15499_, _15495_);
  or _46673_ (_15501_, _15500_, _02459_);
  or _46674_ (_15502_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or _46675_ (_15503_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and _46676_ (_15504_, _15503_, _15502_);
  or _46677_ (_15505_, _15504_, _02445_);
  or _46678_ (_15506_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or _46679_ (_15507_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  and _46680_ (_15508_, _15507_, _15506_);
  or _46681_ (_15509_, _15508_, _02393_);
  and _46682_ (_15510_, _15509_, _15505_);
  or _46683_ (_15511_, _15510_, _02421_);
  and _46684_ (_15512_, _15511_, _02414_);
  and _46685_ (_15513_, _15512_, _15501_);
  or _46686_ (_15514_, _15513_, _15491_);
  and _46687_ (_15515_, _15514_, _02398_);
  or _46688_ (_15516_, _15515_, _15469_);
  and _46689_ (_15517_, _15516_, _02546_);
  and _46690_ (_15518_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and _46691_ (_15519_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or _46692_ (_15520_, _15519_, _15518_);
  and _46693_ (_15521_, _15520_, _02393_);
  and _46694_ (_15522_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  and _46695_ (_15523_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or _46696_ (_15524_, _15523_, _15522_);
  and _46697_ (_15525_, _15524_, _02445_);
  or _46698_ (_15526_, _15525_, _15521_);
  and _46699_ (_15527_, _15526_, _02421_);
  and _46700_ (_15528_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and _46701_ (_15529_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or _46702_ (_15530_, _15529_, _15528_);
  and _46703_ (_15531_, _15530_, _02393_);
  and _46704_ (_15532_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and _46705_ (_15533_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or _46706_ (_15534_, _15533_, _15532_);
  and _46707_ (_15535_, _15534_, _02445_);
  or _46708_ (_15536_, _15535_, _15531_);
  and _46709_ (_15537_, _15536_, _02459_);
  or _46710_ (_15538_, _15537_, _15527_);
  and _46711_ (_15539_, _15538_, _02458_);
  or _46712_ (_15540_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or _46713_ (_15541_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and _46714_ (_15542_, _15541_, _15540_);
  and _46715_ (_15543_, _15542_, _02393_);
  or _46716_ (_15544_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or _46717_ (_15545_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and _46718_ (_15546_, _15545_, _15544_);
  and _46719_ (_15547_, _15546_, _02445_);
  or _46720_ (_15548_, _15547_, _15543_);
  and _46721_ (_15549_, _15548_, _02421_);
  or _46722_ (_15550_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or _46723_ (_15551_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and _46724_ (_15552_, _15551_, _15550_);
  and _46725_ (_15553_, _15552_, _02393_);
  or _46726_ (_15554_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or _46727_ (_15555_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and _46728_ (_15556_, _15555_, _15554_);
  and _46729_ (_15557_, _15556_, _02445_);
  or _46730_ (_15558_, _15557_, _15553_);
  and _46731_ (_15559_, _15558_, _02459_);
  or _46732_ (_15560_, _15559_, _15549_);
  and _46733_ (_15561_, _15560_, _02414_);
  or _46734_ (_15562_, _15561_, _15539_);
  and _46735_ (_15563_, _15562_, _02398_);
  and _46736_ (_15564_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and _46737_ (_15565_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or _46738_ (_15566_, _15565_, _15564_);
  and _46739_ (_15567_, _15566_, _02393_);
  and _46740_ (_15568_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and _46741_ (_15569_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _46742_ (_15570_, _15569_, _15568_);
  and _46743_ (_15571_, _15570_, _02445_);
  or _46744_ (_15572_, _15571_, _15567_);
  and _46745_ (_15573_, _15572_, _02421_);
  and _46746_ (_15574_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and _46747_ (_15575_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or _46748_ (_15576_, _15575_, _15574_);
  and _46749_ (_15577_, _15576_, _02393_);
  and _46750_ (_15578_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and _46751_ (_15579_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _46752_ (_15580_, _15579_, _15578_);
  and _46753_ (_15581_, _15580_, _02445_);
  or _46754_ (_15582_, _15581_, _15577_);
  and _46755_ (_15583_, _15582_, _02459_);
  or _46756_ (_15584_, _15583_, _15573_);
  and _46757_ (_15585_, _15584_, _02458_);
  or _46758_ (_15586_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or _46759_ (_15587_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and _46760_ (_15588_, _15587_, _15586_);
  and _46761_ (_15589_, _15588_, _02393_);
  or _46762_ (_15590_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or _46763_ (_15591_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and _46764_ (_15592_, _15591_, _15590_);
  and _46765_ (_15593_, _15592_, _02445_);
  or _46766_ (_15594_, _15593_, _15589_);
  and _46767_ (_15595_, _15594_, _02421_);
  or _46768_ (_15596_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or _46769_ (_15597_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _46770_ (_15598_, _15597_, _15596_);
  and _46771_ (_15599_, _15598_, _02393_);
  or _46772_ (_15600_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or _46773_ (_15601_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and _46774_ (_15602_, _15601_, _15600_);
  and _46775_ (_15603_, _15602_, _02445_);
  or _46776_ (_15604_, _15603_, _15599_);
  and _46777_ (_15605_, _15604_, _02459_);
  or _46778_ (_15606_, _15605_, _15595_);
  and _46779_ (_15607_, _15606_, _02414_);
  or _46780_ (_15608_, _15607_, _15585_);
  and _46781_ (_15609_, _15608_, _02496_);
  or _46782_ (_15610_, _15609_, _15563_);
  and _46783_ (_15611_, _15610_, _02400_);
  or _46784_ (_15612_, _15611_, _15517_);
  and _46785_ (_15613_, _15612_, _02646_);
  or _46786_ (_15614_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or _46787_ (_15615_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and _46788_ (_15616_, _15615_, _02445_);
  and _46789_ (_15617_, _15616_, _15614_);
  or _46790_ (_15618_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or _46791_ (_15619_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and _46792_ (_15620_, _15619_, _02393_);
  and _46793_ (_15621_, _15620_, _15618_);
  or _46794_ (_15622_, _15621_, _15617_);
  and _46795_ (_15623_, _15622_, _02459_);
  or _46796_ (_15624_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or _46797_ (_15625_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and _46798_ (_15626_, _15625_, _02445_);
  and _46799_ (_15627_, _15626_, _15624_);
  or _46800_ (_15628_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or _46801_ (_15629_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  and _46802_ (_15630_, _15629_, _02393_);
  and _46803_ (_15631_, _15630_, _15628_);
  or _46804_ (_15632_, _15631_, _15627_);
  and _46805_ (_15633_, _15632_, _02421_);
  or _46806_ (_15634_, _15633_, _15623_);
  and _46807_ (_15635_, _15634_, _02414_);
  and _46808_ (_15636_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and _46809_ (_15637_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or _46810_ (_15638_, _15637_, _15636_);
  and _46811_ (_15639_, _15638_, _02393_);
  and _46812_ (_15640_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and _46813_ (_15641_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or _46814_ (_15642_, _15641_, _15640_);
  and _46815_ (_15643_, _15642_, _02445_);
  or _46816_ (_15644_, _15643_, _15639_);
  and _46817_ (_15645_, _15644_, _02459_);
  and _46818_ (_15646_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  and _46819_ (_15647_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or _46820_ (_15648_, _15647_, _15646_);
  and _46821_ (_15649_, _15648_, _02393_);
  and _46822_ (_15650_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and _46823_ (_15651_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or _46824_ (_15652_, _15651_, _15650_);
  and _46825_ (_15653_, _15652_, _02445_);
  or _46826_ (_15654_, _15653_, _15649_);
  and _46827_ (_15655_, _15654_, _02421_);
  or _46828_ (_15656_, _15655_, _15645_);
  and _46829_ (_15657_, _15656_, _02458_);
  or _46830_ (_15658_, _15657_, _15635_);
  and _46831_ (_15659_, _15658_, _02496_);
  or _46832_ (_15660_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or _46833_ (_15661_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and _46834_ (_15662_, _15661_, _15660_);
  and _46835_ (_15663_, _15662_, _02393_);
  or _46836_ (_15664_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or _46837_ (_15665_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and _46838_ (_15666_, _15665_, _15664_);
  and _46839_ (_15667_, _15666_, _02445_);
  or _46840_ (_15668_, _15667_, _15663_);
  and _46841_ (_15669_, _15668_, _02459_);
  or _46842_ (_15670_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or _46843_ (_15671_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and _46844_ (_15672_, _15671_, _15670_);
  and _46845_ (_15673_, _15672_, _02393_);
  or _46846_ (_15674_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or _46847_ (_15675_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and _46848_ (_15676_, _15675_, _15674_);
  and _46849_ (_15677_, _15676_, _02445_);
  or _46850_ (_15678_, _15677_, _15673_);
  and _46851_ (_15679_, _15678_, _02421_);
  or _46852_ (_15680_, _15679_, _15669_);
  and _46853_ (_15681_, _15680_, _02414_);
  and _46854_ (_15682_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and _46855_ (_15683_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or _46856_ (_15684_, _15683_, _15682_);
  and _46857_ (_15685_, _15684_, _02393_);
  and _46858_ (_15686_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and _46859_ (_15687_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or _46860_ (_15688_, _15687_, _15686_);
  and _46861_ (_15689_, _15688_, _02445_);
  or _46862_ (_15690_, _15689_, _15685_);
  and _46863_ (_15691_, _15690_, _02459_);
  and _46864_ (_15692_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and _46865_ (_15693_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or _46866_ (_15694_, _15693_, _15692_);
  and _46867_ (_15695_, _15694_, _02393_);
  and _46868_ (_15696_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and _46869_ (_15697_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or _46870_ (_15698_, _15697_, _15696_);
  and _46871_ (_15699_, _15698_, _02445_);
  or _46872_ (_15700_, _15699_, _15695_);
  and _46873_ (_15701_, _15700_, _02421_);
  or _46874_ (_15702_, _15701_, _15691_);
  and _46875_ (_15703_, _15702_, _02458_);
  or _46876_ (_15704_, _15703_, _15681_);
  and _46877_ (_15705_, _15704_, _02398_);
  or _46878_ (_15706_, _15705_, _15659_);
  and _46879_ (_15707_, _15706_, _02400_);
  and _46880_ (_15708_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and _46881_ (_15709_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or _46882_ (_15710_, _15709_, _15708_);
  and _46883_ (_15711_, _15710_, _02393_);
  and _46884_ (_15712_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and _46885_ (_15713_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or _46886_ (_15714_, _15713_, _15712_);
  and _46887_ (_15715_, _15714_, _02445_);
  or _46888_ (_15716_, _15715_, _15711_);
  or _46889_ (_15717_, _15716_, _02459_);
  and _46890_ (_15718_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and _46891_ (_15719_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or _46892_ (_15720_, _15719_, _15718_);
  and _46893_ (_15721_, _15720_, _02393_);
  and _46894_ (_15722_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and _46895_ (_15723_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or _46896_ (_15724_, _15723_, _15722_);
  and _46897_ (_15725_, _15724_, _02445_);
  or _46898_ (_15726_, _15725_, _15721_);
  or _46899_ (_15727_, _15726_, _02421_);
  and _46900_ (_15728_, _15727_, _02458_);
  and _46901_ (_15729_, _15728_, _15717_);
  or _46902_ (_15730_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or _46903_ (_15731_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and _46904_ (_15732_, _15731_, _15730_);
  and _46905_ (_15733_, _15732_, _02393_);
  or _46906_ (_15734_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or _46907_ (_15735_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and _46908_ (_15736_, _15735_, _15734_);
  and _46909_ (_15737_, _15736_, _02445_);
  or _46910_ (_15738_, _15737_, _15733_);
  or _46911_ (_15739_, _15738_, _02459_);
  or _46912_ (_15740_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or _46913_ (_15741_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and _46914_ (_15742_, _15741_, _15740_);
  and _46915_ (_15743_, _15742_, _02393_);
  or _46916_ (_15744_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or _46917_ (_15745_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and _46918_ (_15746_, _15745_, _15744_);
  and _46919_ (_15747_, _15746_, _02445_);
  or _46920_ (_15748_, _15747_, _15743_);
  or _46921_ (_15749_, _15748_, _02421_);
  and _46922_ (_15750_, _15749_, _02414_);
  and _46923_ (_15751_, _15750_, _15739_);
  or _46924_ (_15752_, _15751_, _15729_);
  and _46925_ (_15753_, _15752_, _02398_);
  and _46926_ (_15754_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and _46927_ (_15755_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or _46928_ (_15756_, _15755_, _15754_);
  and _46929_ (_15757_, _15756_, _02393_);
  and _46930_ (_15758_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and _46931_ (_15759_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or _46932_ (_15760_, _15759_, _15758_);
  and _46933_ (_15761_, _15760_, _02445_);
  or _46934_ (_15762_, _15761_, _15757_);
  or _46935_ (_15763_, _15762_, _02459_);
  and _46936_ (_15764_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and _46937_ (_15765_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or _46938_ (_15766_, _15765_, _15764_);
  and _46939_ (_15767_, _15766_, _02393_);
  and _46940_ (_15768_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and _46941_ (_15769_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or _46942_ (_15770_, _15769_, _15768_);
  and _46943_ (_15771_, _15770_, _02445_);
  or _46944_ (_15772_, _15771_, _15767_);
  or _46945_ (_15773_, _15772_, _02421_);
  and _46946_ (_15774_, _15773_, _02458_);
  and _46947_ (_15775_, _15774_, _15763_);
  or _46948_ (_15776_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or _46949_ (_15777_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  and _46950_ (_15778_, _15777_, _02445_);
  and _46951_ (_15779_, _15778_, _15776_);
  or _46952_ (_15780_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or _46953_ (_15781_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and _46954_ (_15782_, _15781_, _02393_);
  and _46955_ (_15783_, _15782_, _15780_);
  or _46956_ (_15785_, _15783_, _15779_);
  or _46957_ (_15786_, _15785_, _02459_);
  or _46958_ (_15787_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or _46959_ (_15788_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and _46960_ (_15789_, _15788_, _02445_);
  and _46961_ (_15790_, _15789_, _15787_);
  or _46962_ (_15791_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or _46963_ (_15792_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and _46964_ (_15793_, _15792_, _02393_);
  and _46965_ (_15794_, _15793_, _15791_);
  or _46966_ (_15795_, _15794_, _15790_);
  or _46967_ (_15796_, _15795_, _02421_);
  and _46968_ (_15797_, _15796_, _02414_);
  and _46969_ (_15798_, _15797_, _15786_);
  or _46970_ (_15799_, _15798_, _15775_);
  and _46971_ (_15800_, _15799_, _02496_);
  or _46972_ (_15801_, _15800_, _15753_);
  and _46973_ (_15802_, _15801_, _02546_);
  or _46974_ (_15803_, _15802_, _15707_);
  and _46975_ (_15804_, _15803_, _02405_);
  or _46976_ (_15805_, _15804_, _15613_);
  and _46977_ (_15806_, _15805_, _02444_);
  or _46978_ (_15807_, _15806_, _15423_);
  or _46979_ (_15808_, _15807_, _02443_);
  or _46980_ (_15809_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and _46981_ (_15810_, _15809_, _22762_);
  and _46982_ (_05084_, _15810_, _15808_);
  and _46983_ (_15811_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  and _46984_ (_15812_, _14996_, _24050_);
  or _46985_ (_05092_, _15812_, _15811_);
  and _46986_ (_15813_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  and _46987_ (_15814_, _14903_, _23778_);
  or _46988_ (_05094_, _15814_, _15813_);
  and _46989_ (_15815_, _08360_, _23707_);
  and _46990_ (_15816_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  or _46991_ (_05103_, _15816_, _15815_);
  and _46992_ (_15817_, _08360_, _23649_);
  and _46993_ (_15818_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  or _46994_ (_05106_, _15818_, _15817_);
  and _46995_ (_15819_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and _46996_ (_15820_, _12927_, _23898_);
  or _46997_ (_05108_, _15820_, _15819_);
  and _46998_ (_15821_, _08198_, _23824_);
  and _46999_ (_15822_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or _47000_ (_05112_, _15822_, _15821_);
  and _47001_ (_15823_, _05701_, _23824_);
  and _47002_ (_15824_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or _47003_ (_05115_, _15824_, _15823_);
  and _47004_ (_15825_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and _47005_ (_15826_, _12927_, _23824_);
  or _47006_ (_27104_, _15826_, _15825_);
  nand _47007_ (_15827_, _24402_, _22767_);
  or _47008_ (_15828_, _22767_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _47009_ (_15829_, _15828_, _22762_);
  and _47010_ (_26864_[0], _15829_, _15827_);
  and _47011_ (_15830_, _01808_, _24356_);
  and _47012_ (_15831_, _15830_, _23946_);
  not _47013_ (_15832_, _15830_);
  and _47014_ (_15833_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  or _47015_ (_05123_, _15833_, _15831_);
  and _47016_ (_15834_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  and _47017_ (_15835_, _14996_, _23707_);
  or _47018_ (_05124_, _15835_, _15834_);
  and _47019_ (_15836_, _15830_, _23649_);
  and _47020_ (_15837_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  or _47021_ (_05136_, _15837_, _15836_);
  and _47022_ (_15838_, _15830_, _23747_);
  and _47023_ (_15839_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  or _47024_ (_05150_, _15839_, _15838_);
  and _47025_ (_15840_, _15830_, _23824_);
  and _47026_ (_15841_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  or _47027_ (_05155_, _15841_, _15840_);
  and _47028_ (_15842_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and _47029_ (_15843_, _12829_, _23707_);
  or _47030_ (_05179_, _15843_, _15842_);
  and _47031_ (_15844_, _02107_, _23778_);
  and _47032_ (_15845_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  or _47033_ (_27165_, _15845_, _15844_);
  and _47034_ (_15846_, _06886_, _24282_);
  not _47035_ (_15847_, _15846_);
  and _47036_ (_15848_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and _47037_ (_15849_, _15846_, _23649_);
  or _47038_ (_27005_, _15849_, _15848_);
  and _47039_ (_15850_, _23752_, _23076_);
  and _47040_ (_15851_, _15850_, _23824_);
  not _47041_ (_15852_, _15850_);
  and _47042_ (_15853_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  or _47043_ (_05185_, _15853_, _15851_);
  and _47044_ (_15854_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and _47045_ (_15855_, _15846_, _24050_);
  or _47046_ (_27006_, _15855_, _15854_);
  not _47047_ (_15856_, _26110_);
  nor _47048_ (_15857_, _15856_, _24299_);
  or _47049_ (_15858_, _15857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _47050_ (_15859_, _26114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _47051_ (_15860_, _15859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _47052_ (_15861_, _15860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _47053_ (_15862_, _15861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47054_ (_15863_, _15862_, _26100_);
  nand _47055_ (_15864_, _15863_, _12811_);
  or _47056_ (_15865_, _15864_, _24299_);
  and _47057_ (_15866_, _15865_, _15858_);
  or _47058_ (_15867_, _15866_, _24293_);
  nand _47059_ (_15868_, _24293_, _23772_);
  and _47060_ (_15869_, _15868_, _22762_);
  and _47061_ (_05196_, _15869_, _15867_);
  and _47062_ (_15870_, _15830_, _23707_);
  and _47063_ (_15871_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  or _47064_ (_05198_, _15871_, _15870_);
  and _47065_ (_15872_, _15830_, _24050_);
  and _47066_ (_15873_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  or _47067_ (_05202_, _15873_, _15872_);
  nand _47068_ (_15874_, _24508_, _22767_);
  or _47069_ (_15875_, _22767_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _47070_ (_15876_, _15875_, _22762_);
  and _47071_ (_26864_[7], _15876_, _15874_);
  and _47072_ (_15877_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and _47073_ (_15878_, _15846_, _23946_);
  or _47074_ (_05220_, _15878_, _15877_);
  and _47075_ (_15879_, _12733_, _23946_);
  and _47076_ (_15880_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or _47077_ (_05225_, _15880_, _15879_);
  and _47078_ (_15881_, _15830_, _23898_);
  and _47079_ (_15882_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  or _47080_ (_05232_, _15882_, _15881_);
  and _47081_ (_15883_, _15830_, _23778_);
  and _47082_ (_15884_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  or _47083_ (_27164_, _15884_, _15883_);
  and _47084_ (_15885_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  and _47085_ (_15886_, _14996_, _23778_);
  or _47086_ (_27007_, _15886_, _15885_);
  and _47087_ (_15887_, _05187_, _23946_);
  and _47088_ (_15888_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or _47089_ (_05274_, _15888_, _15887_);
  and _47090_ (_15889_, _05187_, _23649_);
  and _47091_ (_15890_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or _47092_ (_05280_, _15890_, _15889_);
  and _47093_ (_15891_, _05187_, _23747_);
  and _47094_ (_15892_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or _47095_ (_05287_, _15892_, _15891_);
  and _47096_ (_15893_, _15850_, _23649_);
  and _47097_ (_15894_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  or _47098_ (_05300_, _15894_, _15893_);
  and _47099_ (_15895_, _24201_, _23784_);
  not _47100_ (_15896_, _15895_);
  and _47101_ (_15897_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  and _47102_ (_15898_, _15895_, _23707_);
  or _47103_ (_05306_, _15898_, _15897_);
  and _47104_ (_15899_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and _47105_ (_15900_, _15846_, _23707_);
  or _47106_ (_05312_, _15900_, _15899_);
  and _47107_ (_15901_, _05114_, _23778_);
  and _47108_ (_15902_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or _47109_ (_05321_, _15902_, _15901_);
  and _47110_ (_15903_, _05187_, _23707_);
  and _47111_ (_15904_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or _47112_ (_05341_, _15904_, _15903_);
  and _47113_ (_15905_, _05187_, _24050_);
  and _47114_ (_15906_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or _47115_ (_27099_, _15906_, _15905_);
  and _47116_ (_15907_, _06886_, _23911_);
  not _47117_ (_15908_, _15907_);
  and _47118_ (_15909_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and _47119_ (_15910_, _15907_, _23707_);
  or _47120_ (_27003_, _15910_, _15909_);
  and _47121_ (_15911_, _24358_, _23707_);
  and _47122_ (_15912_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or _47123_ (_05370_, _15912_, _15911_);
  and _47124_ (_15913_, _24331_, _23946_);
  and _47125_ (_15914_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or _47126_ (_05383_, _15914_, _15913_);
  and _47127_ (_15915_, _24358_, _24050_);
  and _47128_ (_15916_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  or _47129_ (_05386_, _15916_, _15915_);
  and _47130_ (_15917_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  and _47131_ (_15918_, _15895_, _24050_);
  or _47132_ (_05389_, _15918_, _15917_);
  and _47133_ (_15919_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and _47134_ (_15920_, _15846_, _23824_);
  or _47135_ (_05406_, _15920_, _15919_);
  and _47136_ (_15921_, _05187_, _23898_);
  and _47137_ (_15922_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or _47138_ (_05408_, _15922_, _15921_);
  and _47139_ (_15923_, _05187_, _23778_);
  and _47140_ (_15924_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or _47141_ (_05418_, _15924_, _15923_);
  and _47142_ (_15925_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and _47143_ (_15926_, _15846_, _23898_);
  or _47144_ (_05421_, _15926_, _15925_);
  and _47145_ (_15927_, _04811_, _23747_);
  and _47146_ (_15928_, _04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  or _47147_ (_05423_, _15928_, _15927_);
  and _47148_ (_15929_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  and _47149_ (_15930_, _01967_, _23898_);
  or _47150_ (_27233_, _15930_, _15929_);
  and _47151_ (_15931_, _23790_, _23778_);
  and _47152_ (_15932_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  or _47153_ (_27252_, _15932_, _15931_);
  and _47154_ (_15933_, _05114_, _23649_);
  and _47155_ (_15934_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or _47156_ (_05451_, _15934_, _15933_);
  and _47157_ (_15935_, _05114_, _23747_);
  and _47158_ (_15936_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or _47159_ (_05456_, _15936_, _15935_);
  and _47160_ (_15937_, _05114_, _23824_);
  and _47161_ (_15938_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or _47162_ (_05465_, _15938_, _15937_);
  and _47163_ (_15939_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and _47164_ (_15940_, _15907_, _23898_);
  or _47165_ (_05473_, _15940_, _15939_);
  and _47166_ (_15941_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and _47167_ (_15942_, _15907_, _23778_);
  or _47168_ (_05476_, _15942_, _15941_);
  and _47169_ (_15943_, _09913_, _23707_);
  and _47170_ (_15944_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or _47171_ (_05479_, _15944_, _15943_);
  and _47172_ (_15945_, _05114_, _24050_);
  and _47173_ (_15946_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or _47174_ (_05498_, _15946_, _15945_);
  and _47175_ (_15947_, _05114_, _23946_);
  and _47176_ (_15948_, _05117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or _47177_ (_05503_, _15948_, _15947_);
  and _47178_ (_15949_, _08360_, _23898_);
  and _47179_ (_15950_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  or _47180_ (_27086_, _15950_, _15949_);
  and _47181_ (_15951_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and _47182_ (_15952_, _15907_, _23649_);
  or _47183_ (_27001_, _15952_, _15951_);
  and _47184_ (_15953_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and _47185_ (_15954_, _15907_, _23747_);
  or _47186_ (_27000_, _15954_, _15953_);
  and _47187_ (_15955_, _05338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  and _47188_ (_15956_, _05337_, _23898_);
  or _47189_ (_05542_, _15956_, _15955_);
  and _47190_ (_15957_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and _47191_ (_15958_, _12927_, _23707_);
  or _47192_ (_05543_, _15958_, _15957_);
  and _47193_ (_15959_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  and _47194_ (_15960_, _08477_, _23898_);
  or _47195_ (_05546_, _15960_, _15959_);
  and _47196_ (_15961_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and _47197_ (_15962_, _05398_, _24050_);
  or _47198_ (_05549_, _15962_, _15961_);
  and _47199_ (_15963_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  and _47200_ (_15964_, _05358_, _23778_);
  or _47201_ (_05557_, _15964_, _15963_);
  and _47202_ (_15965_, _05371_, _23824_);
  and _47203_ (_15966_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or _47204_ (_05568_, _15966_, _15965_);
  and _47205_ (_15967_, _08360_, _23778_);
  and _47206_ (_15968_, _08362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or _47207_ (_05570_, _15968_, _15967_);
  and _47208_ (_15969_, _05371_, _23649_);
  and _47209_ (_15970_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or _47210_ (_05573_, _15970_, _15969_);
  and _47211_ (_15971_, _13778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and _47212_ (_15972_, _13777_, _23778_);
  or _47213_ (_05577_, _15972_, _15971_);
  and _47214_ (_15973_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  and _47215_ (_15974_, _05358_, _23747_);
  or _47216_ (_05584_, _15974_, _15973_);
  and _47217_ (_15975_, _06886_, _24010_);
  not _47218_ (_15976_, _15975_);
  and _47219_ (_15977_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  and _47220_ (_15978_, _15975_, _23747_);
  or _47221_ (_05589_, _15978_, _15977_);
  and _47222_ (_15979_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  and _47223_ (_15980_, _05354_, _23824_);
  or _47224_ (_05598_, _15980_, _15979_);
  and _47225_ (_15981_, _05706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and _47226_ (_15982_, _05705_, _23898_);
  or _47227_ (_05622_, _15982_, _15981_);
  and _47228_ (_15983_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  and _47229_ (_15984_, _05358_, _23824_);
  or _47230_ (_05625_, _15984_, _15983_);
  and _47231_ (_15985_, _05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  and _47232_ (_15986_, _05354_, _24050_);
  or _47233_ (_05633_, _15986_, _15985_);
  and _47234_ (_15987_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  and _47235_ (_15988_, _12829_, _23824_);
  or _47236_ (_05639_, _15988_, _15987_);
  and _47237_ (_15989_, _05359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  and _47238_ (_15990_, _05358_, _23649_);
  or _47239_ (_05643_, _15990_, _15989_);
  and _47240_ (_15991_, _04760_, _24085_);
  not _47241_ (_15992_, _15991_);
  and _47242_ (_15993_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  and _47243_ (_15994_, _15991_, _24050_);
  or _47244_ (_05659_, _15994_, _15993_);
  and _47245_ (_15995_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  and _47246_ (_15996_, _15991_, _23747_);
  or _47247_ (_05661_, _15996_, _15995_);
  and _47248_ (_15997_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and _47249_ (_15998_, _12829_, _23898_);
  or _47250_ (_27224_, _15998_, _15997_);
  and _47251_ (_15999_, _24699_, _23778_);
  and _47252_ (_16000_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  or _47253_ (_27189_, _16000_, _15999_);
  nand _47254_ (_16001_, _25172_, _23662_);
  or _47255_ (_16002_, _16001_, _00875_);
  not _47256_ (_16003_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _47257_ (_16004_, _16001_, _16003_);
  and _47258_ (_16005_, _16004_, _24069_);
  and _47259_ (_16006_, _16005_, _16002_);
  nor _47260_ (_16007_, _24068_, _16003_);
  and _47261_ (_16008_, _00265_, _25163_);
  and _47262_ (_16009_, _16008_, _24654_);
  nand _47263_ (_16010_, _16009_, _23594_);
  or _47264_ (_16011_, _16009_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _47265_ (_16012_, _16011_, _24645_);
  and _47266_ (_16013_, _16012_, _16010_);
  or _47267_ (_16014_, _16013_, _16007_);
  or _47268_ (_16015_, _16014_, _16006_);
  and _47269_ (_05678_, _16015_, _22762_);
  and _47270_ (_16016_, _15850_, _23747_);
  and _47271_ (_16017_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  or _47272_ (_05689_, _16017_, _16016_);
  and _47273_ (_16018_, _04760_, _23986_);
  not _47274_ (_16019_, _16018_);
  and _47275_ (_16020_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  and _47276_ (_16021_, _16018_, _23898_);
  or _47277_ (_05700_, _16021_, _16020_);
  and _47278_ (_16022_, _24370_, _23903_);
  and _47279_ (_16023_, _16022_, _23649_);
  not _47280_ (_16024_, _16022_);
  and _47281_ (_16025_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or _47282_ (_05707_, _16025_, _16023_);
  and _47283_ (_16026_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and _47284_ (_16027_, _12927_, _24050_);
  or _47285_ (_05754_, _16027_, _16026_);
  and _47286_ (_16028_, _05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and _47287_ (_16029_, _05398_, _23778_);
  or _47288_ (_05769_, _16029_, _16028_);
  and _47289_ (_16030_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  and _47290_ (_16031_, _15991_, _23649_);
  or _47291_ (_05784_, _16031_, _16030_);
  and _47292_ (_16032_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and _47293_ (_16033_, _12927_, _23649_);
  or _47294_ (_05788_, _16033_, _16032_);
  and _47295_ (_16034_, _05701_, _23946_);
  and _47296_ (_16035_, _05703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or _47297_ (_27087_, _16035_, _16034_);
  and _47298_ (_16036_, _06665_, _24050_);
  and _47299_ (_16037_, _06667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  or _47300_ (_27089_, _16037_, _16036_);
  and _47301_ (_16038_, _12928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and _47302_ (_16039_, _12927_, _23946_);
  or _47303_ (_05804_, _16039_, _16038_);
  and _47304_ (_16040_, _24050_, _23833_);
  and _47305_ (_16041_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or _47306_ (_05815_, _16041_, _16040_);
  and _47307_ (_16042_, _05371_, _23946_);
  and _47308_ (_16043_, _05373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or _47309_ (_05842_, _16043_, _16042_);
  and _47310_ (_16044_, _05180_, _23898_);
  and _47311_ (_16045_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or _47312_ (_05849_, _16045_, _16044_);
  and _47313_ (_16046_, _12733_, _23778_);
  and _47314_ (_16047_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  or _47315_ (_05854_, _16047_, _16046_);
  and _47316_ (_16048_, _04760_, _24010_);
  not _47317_ (_16049_, _16048_);
  and _47318_ (_16050_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  and _47319_ (_16051_, _16048_, _23778_);
  or _47320_ (_05862_, _16051_, _16050_);
  and _47321_ (_16052_, _24121_, _23939_);
  nand _47322_ (_16053_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _47323_ (_16054_, _16053_, _24127_);
  nor _47324_ (_16055_, _24151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or _47325_ (_16056_, _16055_, _12951_);
  nand _47326_ (_16057_, _16056_, _12956_);
  or _47327_ (_16058_, _12956_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _47328_ (_16059_, _16058_, _16057_);
  or _47329_ (_16060_, _16059_, _16054_);
  and _47330_ (_16061_, _16060_, _24166_);
  or _47331_ (_05875_, _16061_, _16052_);
  and _47332_ (_16062_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and _47333_ (_16063_, _11746_, _24050_);
  or _47334_ (_27029_, _16063_, _16062_);
  and _47335_ (_16064_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and _47336_ (_16065_, _11746_, _23824_);
  or _47337_ (_27027_, _16065_, _16064_);
  and _47338_ (_16066_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  and _47339_ (_16067_, _15895_, _23778_);
  or _47340_ (_27222_, _16067_, _16066_);
  and _47341_ (_16068_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  and _47342_ (_16069_, _16048_, _23898_);
  or _47343_ (_05899_, _16069_, _16068_);
  and _47344_ (_16070_, _15012_, _23707_);
  and _47345_ (_16071_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or _47346_ (_05905_, _16071_, _16070_);
  and _47347_ (_16072_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  and _47348_ (_16073_, _11729_, _23707_);
  or _47349_ (_05907_, _16073_, _16072_);
  and _47350_ (_16074_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  and _47351_ (_16075_, _11729_, _23898_);
  or _47352_ (_05915_, _16075_, _16074_);
  and _47353_ (_16076_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and _47354_ (_16077_, _11693_, _24050_);
  or _47355_ (_05949_, _16077_, _16076_);
  and _47356_ (_16078_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and _47357_ (_16079_, _11693_, _23824_);
  or _47358_ (_05956_, _16079_, _16078_);
  and _47359_ (_16080_, _12782_, _23649_);
  and _47360_ (_16081_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or _47361_ (_05964_, _16081_, _16080_);
  and _47362_ (_16082_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and _47363_ (_16083_, _11693_, _23778_);
  or _47364_ (_05968_, _16083_, _16082_);
  and _47365_ (_16084_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  and _47366_ (_16085_, _15975_, _23824_);
  or _47367_ (_05971_, _16085_, _16084_);
  and _47368_ (_16086_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and _47369_ (_16087_, _11652_, _23707_);
  or _47370_ (_05974_, _16087_, _16086_);
  and _47371_ (_16088_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and _47372_ (_16089_, _11652_, _23649_);
  or _47373_ (_27025_, _16089_, _16088_);
  and _47374_ (_16090_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  and _47375_ (_16091_, _10494_, _23946_);
  or _47376_ (_05987_, _16091_, _16090_);
  and _47377_ (_16092_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  and _47378_ (_16093_, _15975_, _23898_);
  or _47379_ (_05991_, _16093_, _16092_);
  and _47380_ (_16094_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  and _47381_ (_16095_, _10494_, _23824_);
  or _47382_ (_05995_, _16095_, _16094_);
  and _47383_ (_16096_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  and _47384_ (_16097_, _08375_, _23707_);
  or _47385_ (_06009_, _16097_, _16096_);
  and _47386_ (_16098_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  and _47387_ (_16099_, _08375_, _23824_);
  or _47388_ (_06016_, _16099_, _16098_);
  and _47389_ (_16100_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and _47390_ (_16101_, _06896_, _23747_);
  or _47391_ (_06023_, _16101_, _16100_);
  and _47392_ (_16102_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  and _47393_ (_16103_, _15975_, _24050_);
  or _47394_ (_06031_, _16103_, _16102_);
  and _47395_ (_16104_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  and _47396_ (_16105_, _15975_, _23946_);
  or _47397_ (_06041_, _16105_, _16104_);
  and _47398_ (_16106_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  and _47399_ (_16107_, _07551_, _23747_);
  or _47400_ (_27019_, _16107_, _16106_);
  and _47401_ (_16108_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  and _47402_ (_16109_, _07525_, _24050_);
  or _47403_ (_06051_, _16109_, _16108_);
  and _47404_ (_16110_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  and _47405_ (_16111_, _07525_, _23824_);
  or _47406_ (_27018_, _16111_, _16110_);
  and _47407_ (_16112_, _05180_, _23747_);
  and _47408_ (_16113_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or _47409_ (_27131_, _16113_, _16112_);
  and _47410_ (_16114_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and _47411_ (_16115_, _06927_, _23707_);
  or _47412_ (_06077_, _16115_, _16114_);
  and _47413_ (_16116_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and _47414_ (_16117_, _06927_, _23747_);
  or _47415_ (_06085_, _16117_, _16116_);
  and _47416_ (_16118_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  and _47417_ (_16119_, _16048_, _23824_);
  or _47418_ (_06088_, _16119_, _16118_);
  and _47419_ (_16120_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  and _47420_ (_16121_, _16048_, _23649_);
  or _47421_ (_06093_, _16121_, _16120_);
  and _47422_ (_16122_, _06886_, _24085_);
  not _47423_ (_16123_, _16122_);
  and _47424_ (_16124_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  and _47425_ (_16125_, _16122_, _23946_);
  or _47426_ (_06098_, _16125_, _16124_);
  and _47427_ (_16126_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and _47428_ (_16127_, _06900_, _23707_);
  or _47429_ (_06100_, _16127_, _16126_);
  and _47430_ (_16128_, _24086_, _23778_);
  and _47431_ (_16129_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or _47432_ (_27254_, _16129_, _16128_);
  and _47433_ (_16130_, _02359_, _23649_);
  and _47434_ (_16131_, _02361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  or _47435_ (_06103_, _16131_, _16130_);
  and _47436_ (_16132_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and _47437_ (_16133_, _06900_, _23649_);
  or _47438_ (_27021_, _16133_, _16132_);
  and _47439_ (_16134_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  and _47440_ (_16135_, _16122_, _23649_);
  or _47441_ (_06109_, _16135_, _16134_);
  and _47442_ (_16136_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and _47443_ (_16137_, _06896_, _23898_);
  or _47444_ (_06112_, _16137_, _16136_);
  and _47445_ (_16138_, _04749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  and _47446_ (_16139_, _04748_, _23898_);
  or _47447_ (_06116_, _16139_, _16138_);
  and _47448_ (_16140_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  and _47449_ (_16141_, _16018_, _23824_);
  or _47450_ (_06121_, _16141_, _16140_);
  and _47451_ (_16142_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  and _47452_ (_16143_, _11729_, _23747_);
  or _47453_ (_06123_, _16143_, _16142_);
  and _47454_ (_16144_, _15012_, _24050_);
  and _47455_ (_16145_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or _47456_ (_06131_, _16145_, _16144_);
  and _47457_ (_16146_, _11695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and _47458_ (_16147_, _11693_, _23649_);
  or _47459_ (_06134_, _16147_, _16146_);
  and _47460_ (_16148_, _06639_, _23649_);
  and _47461_ (_16149_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or _47462_ (_06141_, _16149_, _16148_);
  and _47463_ (_16150_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and _47464_ (_16151_, _11652_, _23898_);
  or _47465_ (_06151_, _16151_, _16150_);
  and _47466_ (_16152_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  and _47467_ (_16153_, _08375_, _23649_);
  or _47468_ (_27023_, _16153_, _16152_);
  and _47469_ (_16154_, _06639_, _24050_);
  and _47470_ (_16155_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or _47471_ (_06160_, _16155_, _16154_);
  and _47472_ (_16156_, _08376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  and _47473_ (_16157_, _08375_, _23778_);
  or _47474_ (_06163_, _16157_, _16156_);
  and _47475_ (_16158_, _06897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and _47476_ (_16159_, _06896_, _23946_);
  or _47477_ (_06168_, _16159_, _16158_);
  and _47478_ (_16160_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and _47479_ (_16161_, _06900_, _23778_);
  or _47480_ (_06171_, _16161_, _16160_);
  and _47481_ (_16162_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  and _47482_ (_16163_, _16122_, _23707_);
  or _47483_ (_06176_, _16163_, _16162_);
  and _47484_ (_16164_, _06639_, _23946_);
  and _47485_ (_16165_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or _47486_ (_06178_, _16165_, _16164_);
  and _47487_ (_16166_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  and _47488_ (_16167_, _07551_, _23946_);
  or _47489_ (_06180_, _16167_, _16166_);
  and _47490_ (_16168_, _07552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  and _47491_ (_16169_, _07551_, _23898_);
  or _47492_ (_06184_, _16169_, _16168_);
  and _47493_ (_16170_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and _47494_ (_16171_, _06927_, _23778_);
  or _47495_ (_06205_, _16171_, _16170_);
  or _47496_ (_26862_[0], _05000_, _12899_);
  and _47497_ (_16172_, _24283_, _23747_);
  and _47498_ (_16173_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  or _47499_ (_06233_, _16173_, _16172_);
  and _47500_ (_16174_, _11747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and _47501_ (_16175_, _11746_, _23747_);
  or _47502_ (_27028_, _16175_, _16174_);
  and _47503_ (_16176_, _23992_, _23824_);
  and _47504_ (_16177_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or _47505_ (_26944_, _16177_, _16176_);
  and _47506_ (_16178_, _11653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and _47507_ (_16179_, _11652_, _23946_);
  or _47508_ (_06254_, _16179_, _16178_);
  and _47509_ (_16180_, _10495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  and _47510_ (_16181_, _10494_, _24050_);
  or _47511_ (_06257_, _16181_, _16180_);
  and _47512_ (_16182_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  and _47513_ (_16183_, _16122_, _23778_);
  or _47514_ (_06264_, _16183_, _16182_);
  and _47515_ (_16184_, _25439_, _24118_);
  nand _47516_ (_16185_, _16184_, _23594_);
  or _47517_ (_16186_, _16184_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _47518_ (_16187_, _16186_, _24645_);
  and _47519_ (_16188_, _16187_, _16185_);
  or _47520_ (_16189_, _25447_, _23738_);
  or _47521_ (_16190_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _47522_ (_16191_, _16190_, _24069_);
  and _47523_ (_16192_, _16191_, _16189_);
  and _47524_ (_16193_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _47525_ (_16194_, _16193_, rst);
  or _47526_ (_16195_, _16194_, _16192_);
  or _47527_ (_06267_, _16195_, _16188_);
  and _47528_ (_16196_, _06886_, _23784_);
  not _47529_ (_16197_, _16196_);
  and _47530_ (_16198_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and _47531_ (_16199_, _16196_, _23707_);
  or _47532_ (_06271_, _16199_, _16198_);
  and _47533_ (_16200_, _07526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  and _47534_ (_16201_, _07525_, _23747_);
  or _47535_ (_06273_, _16201_, _16200_);
  and _47536_ (_16202_, _06928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and _47537_ (_16203_, _06927_, _23649_);
  or _47538_ (_06276_, _16203_, _16202_);
  and _47539_ (_16204_, _25350_, _24296_);
  nand _47540_ (_16205_, _16204_, _23594_);
  or _47541_ (_16206_, _16204_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _47542_ (_16207_, _16206_, _24645_);
  and _47543_ (_16208_, _16207_, _16205_);
  or _47544_ (_16209_, _25359_, _23642_);
  or _47545_ (_16210_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _47546_ (_16211_, _16210_, _24069_);
  and _47547_ (_16212_, _16211_, _16209_);
  nor _47548_ (_16213_, _24068_, _06249_);
  or _47549_ (_16214_, _16213_, rst);
  or _47550_ (_16215_, _16214_, _16212_);
  or _47551_ (_06280_, _16215_, _16208_);
  and _47552_ (_16216_, _11730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  and _47553_ (_16217_, _11729_, _23649_);
  or _47554_ (_06289_, _16217_, _16216_);
  and _47555_ (_16218_, _25260_, _24705_);
  nand _47556_ (_16219_, _16218_, _23594_);
  or _47557_ (_16220_, _16218_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _47558_ (_16221_, _16220_, _24645_);
  and _47559_ (_16222_, _16221_, _16219_);
  or _47560_ (_16223_, _25267_, _24043_);
  or _47561_ (_16224_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _47562_ (_16225_, _16224_, _24069_);
  and _47563_ (_16226_, _16225_, _16223_);
  nor _47564_ (_16227_, _24068_, _06185_);
  or _47565_ (_16228_, _16227_, rst);
  or _47566_ (_16229_, _16228_, _16226_);
  or _47567_ (_06293_, _16229_, _16222_);
  and _47568_ (_16230_, _06902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and _47569_ (_16231_, _06900_, _23898_);
  or _47570_ (_27020_, _16231_, _16230_);
  and _47571_ (_16232_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  and _47572_ (_16233_, _16122_, _23824_);
  or _47573_ (_26997_, _16233_, _16232_);
  and _47574_ (_16234_, _25164_, _24296_);
  nand _47575_ (_16235_, _16234_, _23594_);
  or _47576_ (_16237_, _16234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _47577_ (_16238_, _16237_, _24645_);
  and _47578_ (_16239_, _16238_, _16235_);
  or _47579_ (_16240_, _25174_, _23642_);
  or _47580_ (_16241_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _47581_ (_16242_, _16241_, _24069_);
  and _47582_ (_16243_, _16242_, _16240_);
  nor _47583_ (_16244_, _24068_, _06149_);
  or _47584_ (_16245_, _16244_, rst);
  or _47585_ (_16246_, _16245_, _16243_);
  or _47586_ (_06326_, _16246_, _16239_);
  and _47587_ (_16247_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  and _47588_ (_16248_, _12728_, _24050_);
  or _47589_ (_06332_, _16248_, _16247_);
  and _47590_ (_16249_, _12907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and _47591_ (_16250_, _12906_, _23824_);
  or _47592_ (_06338_, _16250_, _16249_);
  and _47593_ (_16251_, _05710_, _23707_);
  and _47594_ (_16252_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  or _47595_ (_06342_, _16252_, _16251_);
  and _47596_ (_16253_, _13757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and _47597_ (_16254_, _13756_, _23649_);
  or _47598_ (_06360_, _16254_, _16253_);
  and _47599_ (_16255_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  and _47600_ (_16256_, _14903_, _23707_);
  or _47601_ (_06364_, _16256_, _16255_);
  and _47602_ (_16257_, _05710_, _24050_);
  and _47603_ (_16258_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  or _47604_ (_06368_, _16258_, _16257_);
  and _47605_ (_16259_, _14904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  and _47606_ (_16260_, _14903_, _23898_);
  or _47607_ (_06370_, _16260_, _16259_);
  and _47608_ (_16261_, _05710_, _23946_);
  and _47609_ (_16262_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  or _47610_ (_27163_, _16262_, _16261_);
  and _47611_ (_16263_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and _47612_ (_16264_, _15907_, _23946_);
  or _47613_ (_27002_, _16264_, _16263_);
  and _47614_ (_16265_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and _47615_ (_16266_, _16196_, _23824_);
  or _47616_ (_06386_, _16266_, _16265_);
  and _47617_ (_16267_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  and _47618_ (_16268_, _15975_, _23778_);
  or _47619_ (_06391_, _16268_, _16267_);
  and _47620_ (_16269_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  and _47621_ (_16270_, _16122_, _23747_);
  or _47622_ (_06395_, _16270_, _16269_);
  and _47623_ (_16271_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and _47624_ (_16272_, _16196_, _23946_);
  or _47625_ (_06398_, _16272_, _16271_);
  and _47626_ (_16273_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and _47627_ (_16274_, _16196_, _23898_);
  or _47628_ (_06401_, _16274_, _16273_);
  and _47629_ (_16275_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and _47630_ (_16276_, _16196_, _23778_);
  or _47631_ (_06403_, _16276_, _16275_);
  and _47632_ (_16277_, _06506_, _23991_);
  not _47633_ (_16278_, _16277_);
  and _47634_ (_16279_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  and _47635_ (_16280_, _16277_, _23824_);
  or _47636_ (_06415_, _16280_, _16279_);
  and _47637_ (_16281_, _06506_, _23903_);
  not _47638_ (_16282_, _16281_);
  and _47639_ (_16283_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  and _47640_ (_16284_, _16281_, _23824_);
  or _47641_ (_26995_, _16284_, _16283_);
  and _47642_ (_16285_, _06506_, _24005_);
  not _47643_ (_16286_, _16285_);
  and _47644_ (_16287_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and _47645_ (_16288_, _16285_, _23649_);
  or _47646_ (_06430_, _16288_, _16287_);
  and _47647_ (_16289_, _06506_, _23986_);
  not _47648_ (_16290_, _16289_);
  and _47649_ (_16291_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and _47650_ (_16292_, _16289_, _23649_);
  or _47651_ (_26991_, _16292_, _16291_);
  and _47652_ (_16293_, _06506_, _23069_);
  not _47653_ (_16294_, _16293_);
  and _47654_ (_16295_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  and _47655_ (_16296_, _16293_, _24050_);
  or _47656_ (_06440_, _16296_, _16295_);
  and _47657_ (_16297_, _06639_, _23778_);
  and _47658_ (_16298_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or _47659_ (_06446_, _16298_, _16297_);
  and _47660_ (_16299_, _06506_, _24329_);
  not _47661_ (_16300_, _16299_);
  and _47662_ (_16301_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and _47663_ (_16302_, _16299_, _23747_);
  or _47664_ (_06450_, _16302_, _16301_);
  and _47665_ (_16303_, _06506_, _23752_);
  not _47666_ (_16304_, _16303_);
  and _47667_ (_16305_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  and _47668_ (_16306_, _16303_, _23778_);
  or _47669_ (_06457_, _16306_, _16305_);
  and _47670_ (_16307_, _06506_, _23656_);
  not _47671_ (_16308_, _16307_);
  and _47672_ (_16309_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and _47673_ (_16310_, _16307_, _23747_);
  or _47674_ (_06461_, _16310_, _16309_);
  and _47675_ (_16311_, _06506_, _24085_);
  not _47676_ (_16312_, _16311_);
  and _47677_ (_16313_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and _47678_ (_16314_, _16311_, _24050_);
  or _47679_ (_06468_, _16314_, _16313_);
  and _47680_ (_16315_, _06639_, _23898_);
  and _47681_ (_16316_, _06643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or _47682_ (_06470_, _16316_, _16315_);
  and _47683_ (_16317_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and _47684_ (_16318_, _16196_, _23649_);
  or _47685_ (_06473_, _16318_, _16317_);
  and _47686_ (_16319_, _04760_, _24275_);
  not _47687_ (_16320_, _16319_);
  and _47688_ (_16321_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  and _47689_ (_16322_, _16319_, _24050_);
  or _47690_ (_06484_, _16322_, _16321_);
  and _47691_ (_16323_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and _47692_ (_16324_, _16196_, _23747_);
  or _47693_ (_06492_, _16324_, _16323_);
  and _47694_ (_16325_, _04760_, _23903_);
  not _47695_ (_16326_, _16325_);
  and _47696_ (_16327_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and _47697_ (_16328_, _16325_, _23946_);
  or _47698_ (_26968_, _16328_, _16327_);
  and _47699_ (_16329_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and _47700_ (_16330_, _16325_, _23898_);
  or _47701_ (_06512_, _16330_, _16329_);
  and _47702_ (_16331_, _04760_, _24005_);
  not _47703_ (_16332_, _16331_);
  and _47704_ (_16333_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  and _47705_ (_16334_, _16331_, _23946_);
  or _47706_ (_06516_, _16334_, _16333_);
  and _47707_ (_16335_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  and _47708_ (_16336_, _16018_, _23707_);
  or _47709_ (_06519_, _16336_, _16335_);
  and _47710_ (_16337_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  and _47711_ (_16338_, _16018_, _23747_);
  or _47712_ (_06521_, _16338_, _16337_);
  and _47713_ (_16339_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and _47714_ (_16340_, _07513_, _24050_);
  or _47715_ (_06523_, _16340_, _16339_);
  and _47716_ (_16341_, _23992_, _23747_);
  and _47717_ (_16342_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or _47718_ (_06526_, _16342_, _16341_);
  and _47719_ (_16343_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and _47720_ (_16344_, _04761_, _23747_);
  or _47721_ (_06528_, _16344_, _16343_);
  and _47722_ (_16345_, _23992_, _23649_);
  and _47723_ (_16346_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or _47724_ (_06535_, _16346_, _16345_);
  and _47725_ (_16347_, _24050_, _23992_);
  and _47726_ (_16348_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or _47727_ (_06537_, _16348_, _16347_);
  and _47728_ (_16349_, _24275_, _23906_);
  and _47729_ (_16350_, _16349_, _23778_);
  not _47730_ (_16351_, _16349_);
  and _47731_ (_16352_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  or _47732_ (_06543_, _16352_, _16350_);
  and _47733_ (_16353_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  and _47734_ (_16354_, _13828_, _24050_);
  or _47735_ (_06546_, _16354_, _16353_);
  and _47736_ (_16355_, _05714_, _23707_);
  and _47737_ (_16356_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  or _47738_ (_27160_, _16356_, _16355_);
  and _47739_ (_16357_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  and _47740_ (_16358_, _14996_, _23824_);
  or _47741_ (_06549_, _16358_, _16357_);
  and _47742_ (_16359_, _06506_, _24275_);
  not _47743_ (_16360_, _16359_);
  and _47744_ (_16361_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and _47745_ (_16362_, _16359_, _23824_);
  or _47746_ (_06556_, _16362_, _16361_);
  and _47747_ (_16363_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and _47748_ (_16364_, _16359_, _23649_);
  or _47749_ (_06560_, _16364_, _16363_);
  and _47750_ (_16365_, _05710_, _23778_);
  and _47751_ (_16366_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  or _47752_ (_06562_, _16366_, _16365_);
  and _47753_ (_16367_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and _47754_ (_16368_, _16359_, _23747_);
  or _47755_ (_06565_, _16368_, _16367_);
  and _47756_ (_16369_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and _47757_ (_16370_, _16359_, _23898_);
  or _47758_ (_06571_, _16370_, _16369_);
  and _47759_ (_16371_, _06506_, _23784_);
  not _47760_ (_16372_, _16371_);
  and _47761_ (_16373_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  and _47762_ (_16374_, _16371_, _23747_);
  or _47763_ (_06591_, _16374_, _16373_);
  and _47764_ (_16375_, _04760_, _23991_);
  not _47765_ (_16376_, _16375_);
  and _47766_ (_16377_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and _47767_ (_16378_, _16375_, _23898_);
  or _47768_ (_06595_, _16378_, _16377_);
  and _47769_ (_16379_, _08167_, _23778_);
  and _47770_ (_16380_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  or _47771_ (_06601_, _16380_, _16379_);
  and _47772_ (_16381_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and _47773_ (_16382_, _04761_, _23707_);
  or _47774_ (_26962_, _16382_, _16381_);
  and _47775_ (_16383_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  and _47776_ (_16384_, _08477_, _23946_);
  or _47777_ (_06611_, _16384_, _16383_);
  and _47778_ (_16385_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and _47779_ (_16386_, _06507_, _24050_);
  or _47780_ (_26979_, _16386_, _16385_);
  and _47781_ (_16387_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and _47782_ (_16388_, _16359_, _24050_);
  or _47783_ (_06617_, _16388_, _16387_);
  and _47784_ (_16389_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and _47785_ (_16390_, _15907_, _24050_);
  or _47786_ (_06631_, _16390_, _16389_);
  and _47787_ (_16391_, _16197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and _47788_ (_16392_, _16196_, _24050_);
  or _47789_ (_06633_, _16392_, _16391_);
  and _47790_ (_16393_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  and _47791_ (_16394_, _16281_, _23747_);
  or _47792_ (_06635_, _16394_, _16393_);
  and _47793_ (_16395_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  and _47794_ (_16396_, _16303_, _23898_);
  or _47795_ (_06638_, _16396_, _16395_);
  and _47796_ (_16397_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and _47797_ (_16398_, _16359_, _23707_);
  or _47798_ (_06640_, _16398_, _16397_);
  and _47799_ (_16399_, _08167_, _23824_);
  and _47800_ (_16400_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  or _47801_ (_06642_, _16400_, _16399_);
  and _47802_ (_16401_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and _47803_ (_16402_, _16311_, _23707_);
  or _47804_ (_06645_, _16402_, _16401_);
  and _47805_ (_16403_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  and _47806_ (_16404_, _16319_, _23824_);
  or _47807_ (_06648_, _16404_, _16403_);
  and _47808_ (_16405_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  and _47809_ (_16406_, _10331_, _23824_);
  or _47810_ (_06660_, _16406_, _16405_);
  and _47811_ (_16407_, _05710_, _23747_);
  and _47812_ (_16408_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  or _47813_ (_27161_, _16408_, _16407_);
  and _47814_ (_16409_, _05710_, _23824_);
  and _47815_ (_16410_, _05712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  or _47816_ (_06664_, _16410_, _16409_);
  and _47817_ (_16411_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  and _47818_ (_16412_, _16277_, _23946_);
  or _47819_ (_26996_, _16412_, _16411_);
  and _47820_ (_16413_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  and _47821_ (_16414_, _10331_, _23898_);
  or _47822_ (_26982_, _16414_, _16413_);
  and _47823_ (_16415_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and _47824_ (_16416_, _06507_, _23824_);
  or _47825_ (_06679_, _16416_, _16415_);
  and _47826_ (_16417_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and _47827_ (_16418_, _06507_, _23778_);
  or _47828_ (_06684_, _16418_, _16417_);
  and _47829_ (_16419_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and _47830_ (_16420_, _06507_, _23946_);
  or _47831_ (_06689_, _16420_, _16419_);
  and _47832_ (_16421_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  and _47833_ (_16422_, _16277_, _23649_);
  or _47834_ (_06695_, _16422_, _16421_);
  and _47835_ (_16423_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and _47836_ (_16424_, _06507_, _23707_);
  or _47837_ (_06702_, _16424_, _16423_);
  and _47838_ (_16425_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  and _47839_ (_16426_, _08477_, _23649_);
  or _47840_ (_06705_, _16426_, _16425_);
  and _47841_ (_16427_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  and _47842_ (_16428_, _16277_, _23747_);
  or _47843_ (_06707_, _16428_, _16427_);
  and _47844_ (_16429_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and _47845_ (_16430_, _04761_, _23824_);
  or _47846_ (_06709_, _16430_, _16429_);
  and _47847_ (_16431_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and _47848_ (_16432_, _04761_, _24050_);
  or _47849_ (_06711_, _16432_, _16431_);
  and _47850_ (_16433_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and _47851_ (_16434_, _04761_, _23946_);
  or _47852_ (_06714_, _16434_, _16433_);
  and _47853_ (_16435_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and _47854_ (_16436_, _07513_, _23824_);
  or _47855_ (_26964_, _16436_, _16435_);
  and _47856_ (_16437_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and _47857_ (_16438_, _07513_, _23778_);
  or _47858_ (_06721_, _16438_, _16437_);
  or _47859_ (_16439_, _16001_, _26565_);
  not _47860_ (_16440_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _47861_ (_16441_, _16001_, _16440_);
  and _47862_ (_16442_, _16441_, _24069_);
  and _47863_ (_16443_, _16442_, _16439_);
  nor _47864_ (_16444_, _24068_, _16440_);
  or _47865_ (_16445_, _16001_, _23711_);
  and _47866_ (_16446_, _16441_, _24645_);
  and _47867_ (_16447_, _16446_, _16445_);
  or _47868_ (_16448_, _16447_, _16444_);
  or _47869_ (_16449_, _16448_, _16443_);
  and _47870_ (_06742_, _16449_, _22762_);
  or _47871_ (_16450_, _16001_, _00451_);
  not _47872_ (_16451_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _47873_ (_16452_, _16001_, _16451_);
  and _47874_ (_16453_, _16452_, _24069_);
  and _47875_ (_16454_, _16453_, _16450_);
  nor _47876_ (_16456_, _24068_, _16451_);
  and _47877_ (_16457_, _16008_, _24291_);
  nand _47878_ (_16458_, _16457_, _23594_);
  or _47879_ (_16459_, _16457_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _47880_ (_16460_, _16459_, _24645_);
  and _47881_ (_16461_, _16460_, _16458_);
  or _47882_ (_16462_, _16461_, _16456_);
  or _47883_ (_16463_, _16462_, _16454_);
  and _47884_ (_06744_, _16463_, _22762_);
  or _47885_ (_16464_, _16001_, _00373_);
  not _47886_ (_16465_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _47887_ (_16466_, _16001_, _16465_);
  and _47888_ (_16467_, _16466_, _24069_);
  and _47889_ (_16468_, _16467_, _16464_);
  nor _47890_ (_16469_, _24068_, _16465_);
  and _47891_ (_16470_, _16008_, _24067_);
  nand _47892_ (_16471_, _16470_, _23594_);
  or _47893_ (_16472_, _16470_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _47894_ (_16473_, _16472_, _24645_);
  and _47895_ (_16474_, _16473_, _16471_);
  or _47896_ (_16475_, _16474_, _16469_);
  or _47897_ (_16476_, _16475_, _16468_);
  and _47898_ (_06745_, _16476_, _22762_);
  and _47899_ (_16477_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and _47900_ (_16478_, _07513_, _23649_);
  or _47901_ (_06748_, _16478_, _16477_);
  or _47902_ (_16479_, _16001_, _00545_);
  not _47903_ (_16480_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _47904_ (_16481_, _16001_, _16480_);
  and _47905_ (_16482_, _16481_, _24069_);
  and _47906_ (_16483_, _16482_, _16479_);
  nor _47907_ (_16484_, _24068_, _16480_);
  and _47908_ (_16485_, _16008_, _24118_);
  nand _47909_ (_16486_, _16485_, _23594_);
  or _47910_ (_16487_, _16485_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _47911_ (_16488_, _16487_, _24645_);
  and _47912_ (_16489_, _16488_, _16486_);
  or _47913_ (_16490_, _16489_, _16484_);
  or _47914_ (_16491_, _16490_, _16483_);
  and _47915_ (_06752_, _16491_, _22762_);
  and _47916_ (_16492_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  and _47917_ (_16493_, _16018_, _23778_);
  or _47918_ (_06754_, _16493_, _16492_);
  and _47919_ (_16494_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  and _47920_ (_16495_, _16277_, _24050_);
  or _47921_ (_06758_, _16495_, _16494_);
  and _47922_ (_16496_, _05714_, _23824_);
  and _47923_ (_16497_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  or _47924_ (_27159_, _16497_, _16496_);
  or _47925_ (_16498_, _16001_, _00708_);
  not _47926_ (_16499_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _47927_ (_16500_, _16001_, _16499_);
  and _47928_ (_16501_, _16500_, _24069_);
  and _47929_ (_16502_, _16501_, _16498_);
  nor _47930_ (_16503_, _24068_, _16499_);
  and _47931_ (_16504_, _16008_, _24125_);
  nand _47932_ (_16505_, _16504_, _23594_);
  or _47933_ (_16506_, _16504_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _47934_ (_16507_, _16506_, _24645_);
  and _47935_ (_16508_, _16507_, _16505_);
  or _47936_ (_16509_, _16508_, _16503_);
  or _47937_ (_16510_, _16509_, _16502_);
  and _47938_ (_06760_, _16510_, _22762_);
  or _47939_ (_16511_, _16001_, _00620_);
  not _47940_ (_16512_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _47941_ (_16513_, _16001_, _16512_);
  and _47942_ (_16514_, _16513_, _24069_);
  and _47943_ (_16515_, _16514_, _16511_);
  nor _47944_ (_16516_, _24068_, _16512_);
  not _47945_ (_16517_, _16008_);
  or _47946_ (_16518_, _16517_, _24751_);
  and _47947_ (_16519_, _16518_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _47948_ (_16520_, _23065_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _47949_ (_16521_, _16520_, _24745_);
  and _47950_ (_16522_, _16521_, _16008_);
  or _47951_ (_16523_, _16522_, _16519_);
  and _47952_ (_16524_, _16523_, _24645_);
  or _47953_ (_16525_, _16524_, _16516_);
  or _47954_ (_16526_, _16525_, _16515_);
  and _47955_ (_06762_, _16526_, _22762_);
  and _47956_ (_16527_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  and _47957_ (_16528_, _16277_, _23707_);
  or _47958_ (_06765_, _16528_, _16527_);
  or _47959_ (_16529_, _16001_, _00794_);
  not _47960_ (_16530_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _47961_ (_16531_, _16001_, _16530_);
  and _47962_ (_16532_, _16531_, _24069_);
  and _47963_ (_16533_, _16532_, _16529_);
  nor _47964_ (_16534_, _24068_, _16530_);
  and _47965_ (_16535_, _16008_, _24705_);
  nand _47966_ (_16536_, _16535_, _23594_);
  or _47967_ (_16537_, _16535_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _47968_ (_16538_, _16537_, _24645_);
  and _47969_ (_16539_, _16538_, _16536_);
  or _47970_ (_16540_, _16539_, _16534_);
  or _47971_ (_16541_, _16540_, _16533_);
  and _47972_ (_06767_, _16541_, _22762_);
  and _47973_ (_16542_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  and _47974_ (_16543_, _16331_, _23824_);
  or _47975_ (_06770_, _16543_, _16542_);
  and _47976_ (_16544_, _24639_, _23778_);
  and _47977_ (_16545_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or _47978_ (_06777_, _16545_, _16544_);
  and _47979_ (_16546_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and _47980_ (_16547_, _16375_, _23778_);
  or _47981_ (_06782_, _16547_, _16546_);
  and _47982_ (_16548_, _05714_, _23898_);
  and _47983_ (_16549_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  or _47984_ (_06784_, _16549_, _16548_);
  and _47985_ (_16550_, _01810_, _23707_);
  and _47986_ (_16551_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or _47987_ (_06787_, _16551_, _16550_);
  and _47988_ (_16552_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and _47989_ (_16553_, _16325_, _23707_);
  or _47990_ (_06790_, _16553_, _16552_);
  and _47991_ (_16554_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and _47992_ (_16555_, _16375_, _23946_);
  or _47993_ (_06793_, _16555_, _16554_);
  and _47994_ (_16556_, _24121_, _26750_);
  nand _47995_ (_16557_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47996_ (_16558_, _16557_, _24127_);
  nor _47997_ (_16559_, _12952_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or _47998_ (_16560_, _16559_, _24154_);
  nand _47999_ (_16561_, _16560_, _12956_);
  or _48000_ (_16562_, _12956_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _48001_ (_16563_, _16562_, _16561_);
  or _48002_ (_16564_, _16563_, _16558_);
  and _48003_ (_16565_, _16564_, _24166_);
  or _48004_ (_06794_, _16565_, _16556_);
  and _48005_ (_16566_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  and _48006_ (_16567_, _16319_, _23898_);
  or _48007_ (_06802_, _16567_, _16566_);
  and _48008_ (_16568_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  and _48009_ (_16569_, _16319_, _23649_);
  or _48010_ (_06812_, _16569_, _16568_);
  and _48011_ (_16570_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  and _48012_ (_16571_, _16371_, _23824_);
  or _48013_ (_26973_, _16571_, _16570_);
  and _48014_ (_16572_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and _48015_ (_16573_, _16311_, _23778_);
  or _48016_ (_06824_, _16573_, _16572_);
  and _48017_ (_16574_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  and _48018_ (_16575_, _16371_, _24050_);
  or _48019_ (_06831_, _16575_, _16574_);
  and _48020_ (_16576_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and _48021_ (_16577_, _16311_, _23747_);
  or _48022_ (_06833_, _16577_, _16576_);
  and _48023_ (_16578_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  and _48024_ (_16579_, _16281_, _24050_);
  or _48025_ (_06837_, _16579_, _16578_);
  and _48026_ (_16580_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  and _48027_ (_16581_, _16281_, _23946_);
  or _48028_ (_06859_, _16581_, _16580_);
  and _48029_ (_16582_, _06506_, _25078_);
  not _48030_ (_16583_, _16582_);
  and _48031_ (_16584_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and _48032_ (_16585_, _16582_, _24050_);
  or _48033_ (_06864_, _16585_, _16584_);
  or _48034_ (_16586_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _48035_ (_16587_, _16586_, _22762_);
  nand _48036_ (_16588_, _24078_, _23702_);
  and _48037_ (_06866_, _16588_, _16587_);
  and _48038_ (_16589_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  and _48039_ (_16590_, _16281_, _23649_);
  or _48040_ (_06869_, _16590_, _16589_);
  and _48041_ (_16591_, _02200_, _23707_);
  and _48042_ (_16592_, _02202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or _48043_ (_27168_, _16592_, _16591_);
  and _48044_ (_16593_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  and _48045_ (_16594_, _16303_, _24050_);
  or _48046_ (_06885_, _16594_, _16593_);
  and _48047_ (_16595_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  and _48048_ (_16596_, _16303_, _23747_);
  or _48049_ (_06887_, _16596_, _16595_);
  and _48050_ (_16597_, _05714_, _23649_);
  and _48051_ (_16598_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  or _48052_ (_06891_, _16598_, _16597_);
  and _48053_ (_16599_, _06506_, _01808_);
  not _48054_ (_16600_, _16599_);
  and _48055_ (_16601_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  and _48056_ (_16602_, _16599_, _23898_);
  or _48057_ (_26987_, _16602_, _16601_);
  and _48058_ (_16603_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and _48059_ (_16604_, _16299_, _23707_);
  or _48060_ (_06901_, _16604_, _16603_);
  and _48061_ (_16605_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  and _48062_ (_16606_, _16277_, _23898_);
  or _48063_ (_06911_, _16606_, _16605_);
  and _48064_ (_16607_, _16349_, _23898_);
  and _48065_ (_16608_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  or _48066_ (_06913_, _16608_, _16607_);
  and _48067_ (_16609_, _05714_, _23747_);
  and _48068_ (_16610_, _05716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  or _48069_ (_06915_, _16610_, _16609_);
  and _48070_ (_16611_, _16278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  and _48071_ (_16612_, _16277_, _23778_);
  or _48072_ (_06917_, _16612_, _16611_);
  and _48073_ (_16613_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and _48074_ (_16614_, _16289_, _23778_);
  or _48075_ (_06923_, _16614_, _16613_);
  and _48076_ (_16615_, _05350_, _23747_);
  and _48077_ (_16616_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  or _48078_ (_06925_, _16616_, _16615_);
  and _48079_ (_16617_, _16349_, _23747_);
  and _48080_ (_16618_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  or _48081_ (_06926_, _16618_, _16617_);
  and _48082_ (_16619_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and _48083_ (_16620_, _16285_, _24050_);
  or _48084_ (_06929_, _16620_, _16619_);
  and _48085_ (_16621_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  and _48086_ (_16622_, _16281_, _23707_);
  or _48087_ (_06932_, _16622_, _16621_);
  and _48088_ (_16623_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and _48089_ (_16624_, _16359_, _23778_);
  or _48090_ (_06938_, _16624_, _16623_);
  and _48091_ (_06939_, _26682_, _22762_);
  and _48092_ (_06960_, _26727_, _22762_);
  and _48093_ (_16625_, _16360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and _48094_ (_16626_, _16359_, _23946_);
  or _48095_ (_06965_, _16626_, _16625_);
  and _48096_ (_16627_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  and _48097_ (_16628_, _16122_, _23898_);
  or _48098_ (_06969_, _16628_, _16627_);
  and _48099_ (_16629_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  and _48100_ (_16630_, _16122_, _24050_);
  or _48101_ (_06972_, _16630_, _16629_);
  and _48102_ (_16631_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  and _48103_ (_16632_, _15975_, _23707_);
  or _48104_ (_06974_, _16632_, _16631_);
  and _48105_ (_16633_, _15976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  and _48106_ (_16634_, _15975_, _23649_);
  or _48107_ (_26998_, _16634_, _16633_);
  and _48108_ (_16635_, _15908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and _48109_ (_16636_, _15907_, _23824_);
  or _48110_ (_26999_, _16636_, _16635_);
  and _48111_ (_16637_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and _48112_ (_16638_, _15846_, _23747_);
  or _48113_ (_27004_, _16638_, _16637_);
  and _48114_ (_16639_, _06646_, _23649_);
  and _48115_ (_16640_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or _48116_ (_06986_, _16640_, _16639_);
  and _48117_ (_16641_, _15847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and _48118_ (_16642_, _15846_, _23778_);
  or _48119_ (_06994_, _16642_, _16641_);
  and _48120_ (_16643_, _14997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  and _48121_ (_16644_, _14996_, _23898_);
  or _48122_ (_06999_, _16644_, _16643_);
  and _48123_ (_16645_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and _48124_ (_16646_, _16285_, _23946_);
  or _48125_ (_07013_, _16646_, _16645_);
  and _48126_ (_16647_, _13895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and _48127_ (_16648_, _13894_, _24050_);
  or _48128_ (_07018_, _16648_, _16647_);
  and _48129_ (_16649_, _13829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  and _48130_ (_16650_, _13828_, _23946_);
  or _48131_ (_07022_, _16650_, _16649_);
  and _48132_ (_16651_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  and _48133_ (_16652_, _16281_, _23898_);
  or _48134_ (_26994_, _16652_, _16651_);
  and _48135_ (_16653_, _12729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  and _48136_ (_16654_, _12728_, _23747_);
  or _48137_ (_07053_, _16654_, _16653_);
  and _48138_ (_16655_, _06889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  and _48139_ (_16656_, _06888_, _23747_);
  or _48140_ (_07055_, _16656_, _16655_);
  and _48141_ (_16657_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and _48142_ (_16658_, _06918_, _23778_);
  or _48143_ (_27015_, _16658_, _16657_);
  and _48144_ (_16659_, _16282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  and _48145_ (_16660_, _16281_, _23778_);
  or _48146_ (_07061_, _16660_, _16659_);
  and _48147_ (_16661_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  and _48148_ (_16662_, _16285_, _23707_);
  or _48149_ (_07081_, _16662_, _16661_);
  and _48150_ (_16663_, _12782_, _23747_);
  and _48151_ (_16664_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or _48152_ (_07086_, _16664_, _16663_);
  and _48153_ (_16665_, _06646_, _23707_);
  and _48154_ (_16666_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or _48155_ (_07089_, _16666_, _16665_);
  and _48156_ (_16667_, _06646_, _24050_);
  and _48157_ (_16668_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or _48158_ (_07092_, _16668_, _16667_);
  and _48159_ (_16669_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and _48160_ (_16670_, _16289_, _23946_);
  or _48161_ (_07098_, _16670_, _16669_);
  and _48162_ (_16671_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and _48163_ (_16672_, _16289_, _23707_);
  or _48164_ (_07106_, _16672_, _16671_);
  and _48165_ (_16673_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and _48166_ (_16674_, _16289_, _24050_);
  or _48167_ (_07110_, _16674_, _16673_);
  and _48168_ (_16675_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and _48169_ (_16676_, _16285_, _23747_);
  or _48170_ (_07150_, _16676_, _16675_);
  and _48171_ (_16677_, _06755_, _23707_);
  and _48172_ (_16678_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or _48173_ (_27158_, _16678_, _16677_);
  and _48174_ (_16679_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and _48175_ (_16680_, _16285_, _23824_);
  or _48176_ (_07173_, _16680_, _16679_);
  and _48177_ (_16681_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and _48178_ (_16682_, _16285_, _23898_);
  or _48179_ (_26993_, _16682_, _16681_);
  and _48180_ (_16683_, _06755_, _24050_);
  and _48181_ (_16684_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or _48182_ (_07191_, _16684_, _16683_);
  and _48183_ (_16685_, _16286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and _48184_ (_16686_, _16285_, _23778_);
  or _48185_ (_07195_, _16686_, _16685_);
  and _48186_ (_16687_, _10347_, _24050_);
  and _48187_ (_16688_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  or _48188_ (_07203_, _16688_, _16687_);
  nand _48189_ (_07218_, _00077_, _22762_);
  nand _48190_ (_07222_, _00112_, _22762_);
  nor _48191_ (_07226_, _00029_, rst);
  nor _48192_ (_07228_, _00046_, rst);
  nand _48193_ (_07231_, _00147_, _22762_);
  nor _48194_ (_07237_, _26788_, rst);
  nor _48195_ (_07241_, _26826_, rst);
  and _48196_ (_16689_, _05350_, _23649_);
  and _48197_ (_16690_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  or _48198_ (_07244_, _16690_, _16689_);
  and _48199_ (_16691_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  and _48200_ (_16692_, _16293_, _23707_);
  or _48201_ (_07246_, _16692_, _16691_);
  and _48202_ (_16693_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and _48203_ (_16694_, _24692_, _23778_);
  or _48204_ (_07250_, _16694_, _16693_);
  and _48205_ (_16695_, _06646_, _23898_);
  and _48206_ (_16696_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or _48207_ (_07253_, _16696_, _16695_);
  and _48208_ (_16697_, _06646_, _23778_);
  and _48209_ (_16698_, _06649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or _48210_ (_07278_, _16698_, _16697_);
  and _48211_ (_16699_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and _48212_ (_16700_, _01967_, _23778_);
  or _48213_ (_07282_, _16700_, _16699_);
  and _48214_ (_16701_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and _48215_ (_16702_, _16289_, _23898_);
  or _48216_ (_07287_, _16702_, _16701_);
  and _48217_ (_16703_, _15850_, _24050_);
  and _48218_ (_16704_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  or _48219_ (_07290_, _16704_, _16703_);
  nand _48220_ (_16705_, _25644_, _24598_);
  or _48221_ (_26862_[2], _16705_, _04996_);
  and _48222_ (_16706_, _25649_, _23898_);
  and _48223_ (_16707_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or _48224_ (_07300_, _16707_, _16706_);
  and _48225_ (_16708_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and _48226_ (_16709_, _16289_, _23747_);
  or _48227_ (_07305_, _16709_, _16708_);
  and _48228_ (_16710_, _16290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and _48229_ (_16711_, _16289_, _23824_);
  or _48230_ (_07310_, _16711_, _16710_);
  nor _48231_ (_26885_[4], _25919_, rst);
  and _48232_ (_26886_[7], _26752_, _22762_);
  and _48233_ (_16712_, _06755_, _23824_);
  and _48234_ (_16713_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or _48235_ (_07338_, _16713_, _16712_);
  and _48236_ (_16714_, _23946_, _23833_);
  and _48237_ (_16715_, _23835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or _48238_ (_07342_, _16715_, _16714_);
  and _48239_ (_26884_, _26777_, _22762_);
  and _48240_ (_16716_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  and _48241_ (_16717_, _16293_, _23747_);
  or _48242_ (_26989_, _16717_, _16716_);
  and _48243_ (_16718_, _06755_, _23898_);
  and _48244_ (_16719_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or _48245_ (_07359_, _16719_, _16718_);
  and _48246_ (_16720_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  and _48247_ (_16721_, _16293_, _23824_);
  or _48248_ (_07363_, _16721_, _16720_);
  and _48249_ (_16722_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  and _48250_ (_16723_, _16293_, _23898_);
  or _48251_ (_07390_, _16723_, _16722_);
  and _48252_ (_16724_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  and _48253_ (_16725_, _16293_, _23778_);
  or _48254_ (_07396_, _16725_, _16724_);
  and _48255_ (_16726_, _24699_, _24050_);
  and _48256_ (_16727_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  or _48257_ (_07402_, _16727_, _16726_);
  and _48258_ (_16728_, _08167_, _23649_);
  and _48259_ (_16729_, _08169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  or _48260_ (_07408_, _16729_, _16728_);
  and _48261_ (_16730_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and _48262_ (_16731_, _06918_, _23946_);
  or _48263_ (_07416_, _16731_, _16730_);
  and _48264_ (_16732_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and _48265_ (_16733_, _06918_, _23747_);
  or _48266_ (_07425_, _16733_, _16732_);
  and _48267_ (_16734_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  and _48268_ (_16735_, _16293_, _23946_);
  or _48269_ (_07428_, _16735_, _16734_);
  and _48270_ (_16736_, _06919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and _48271_ (_16737_, _06918_, _23824_);
  or _48272_ (_27016_, _16737_, _16736_);
  and _48273_ (_16738_, _06755_, _23649_);
  and _48274_ (_16739_, _06757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or _48275_ (_07435_, _16739_, _16738_);
  and _48276_ (_16740_, _16294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  and _48277_ (_16741_, _16293_, _23649_);
  or _48278_ (_26990_, _16741_, _16740_);
  and _48279_ (_16742_, _04760_, _24329_);
  not _48280_ (_16743_, _16742_);
  and _48281_ (_16744_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  and _48282_ (_16745_, _16742_, _23946_);
  or _48283_ (_07441_, _16745_, _16744_);
  and _48284_ (_16746_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  and _48285_ (_16747_, _16742_, _23747_);
  or _48286_ (_07445_, _16747_, _16746_);
  and _48287_ (_16748_, _04760_, _23752_);
  not _48288_ (_16749_, _16748_);
  and _48289_ (_16750_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and _48290_ (_16751_, _16748_, _23649_);
  or _48291_ (_07453_, _16751_, _16750_);
  and _48292_ (_16752_, _04760_, _23656_);
  not _48293_ (_16753_, _16752_);
  and _48294_ (_16754_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  and _48295_ (_16755_, _16752_, _23747_);
  or _48296_ (_07481_, _16755_, _16754_);
  and _48297_ (_16756_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  and _48298_ (_16757_, _16599_, _23649_);
  or _48299_ (_07485_, _16757_, _16756_);
  and _48300_ (_16758_, _04760_, _25078_);
  not _48301_ (_16759_, _16758_);
  and _48302_ (_16760_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  and _48303_ (_16761_, _16758_, _23747_);
  or _48304_ (_07487_, _16761_, _16760_);
  and _48305_ (_16762_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  and _48306_ (_16763_, _16599_, _23747_);
  or _48307_ (_07491_, _16763_, _16762_);
  and _48308_ (_16764_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  and _48309_ (_16765_, _16599_, _23824_);
  or _48310_ (_07495_, _16765_, _16764_);
  and _48311_ (_16766_, _04760_, _24282_);
  not _48312_ (_16767_, _16766_);
  and _48313_ (_16768_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and _48314_ (_16769_, _16766_, _23649_);
  or _48315_ (_07498_, _16769_, _16768_);
  and _48316_ (_16770_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and _48317_ (_16771_, _16766_, _23824_);
  or _48318_ (_26951_, _16771_, _16770_);
  and _48319_ (_16772_, _04760_, _23911_);
  not _48320_ (_16773_, _16772_);
  and _48321_ (_16774_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and _48322_ (_16775_, _16772_, _23649_);
  or _48323_ (_26948_, _16775_, _16774_);
  and _48324_ (_16776_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  and _48325_ (_16777_, _15991_, _23898_);
  or _48326_ (_07507_, _16777_, _16776_);
  and _48327_ (_16778_, _06651_, _23778_);
  and _48328_ (_16779_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  or _48329_ (_27152_, _16779_, _16778_);
  and _48330_ (_16780_, _04760_, _23784_);
  not _48331_ (_16781_, _16780_);
  and _48332_ (_16782_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and _48333_ (_16783_, _16780_, _24050_);
  or _48334_ (_07520_, _16783_, _16782_);
  and _48335_ (_16784_, _06511_, _23707_);
  and _48336_ (_16785_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or _48337_ (_07523_, _16785_, _16784_);
  and _48338_ (_16786_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and _48339_ (_16787_, _16780_, _23778_);
  or _48340_ (_07529_, _16787_, _16786_);
  and _48341_ (_16788_, _16022_, _24050_);
  and _48342_ (_16789_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or _48343_ (_07531_, _16789_, _16788_);
  and _48344_ (_16790_, _16349_, _23946_);
  and _48345_ (_16791_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  or _48346_ (_07532_, _16791_, _16790_);
  and _48347_ (_16792_, _15850_, _23946_);
  and _48348_ (_16793_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  or _48349_ (_07535_, _16793_, _16792_);
  and _48350_ (_16794_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  and _48351_ (_16795_, _16599_, _23707_);
  or _48352_ (_07538_, _16795_, _16794_);
  and _48353_ (_16796_, _23992_, _23946_);
  and _48354_ (_16797_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or _48355_ (_07540_, _16797_, _16796_);
  and _48356_ (_16798_, _08307_, _24067_);
  nand _48357_ (_16799_, _16798_, _23594_);
  or _48358_ (_16800_, _16798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _48359_ (_16801_, _16800_, _12774_);
  and _48360_ (_16802_, _16801_, _16799_);
  and _48361_ (_16803_, _08313_, _23892_);
  or _48362_ (_16804_, _16803_, _16802_);
  and _48363_ (_07546_, _16804_, _22762_);
  and _48364_ (_16805_, _08307_, _24678_);
  nand _48365_ (_16806_, _16805_, _23594_);
  or _48366_ (_16807_, _16805_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _48367_ (_16808_, _16807_, _12774_);
  and _48368_ (_16809_, _16808_, _16806_);
  and _48369_ (_16810_, _08313_, _24685_);
  or _48370_ (_16811_, _16810_, _16809_);
  and _48371_ (_07549_, _16811_, _22762_);
  and _48372_ (_16812_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  and _48373_ (_16813_, _16048_, _23747_);
  or _48374_ (_26946_, _16813_, _16812_);
  and _48375_ (_16814_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  and _48376_ (_16815_, _16599_, _24050_);
  or _48377_ (_07561_, _16815_, _16814_);
  and _48378_ (_16816_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  and _48379_ (_16817_, _16599_, _23946_);
  or _48380_ (_26988_, _16817_, _16816_);
  and _48381_ (_16818_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  and _48382_ (_16819_, _15991_, _23946_);
  or _48383_ (_07564_, _16819_, _16818_);
  and _48384_ (_16820_, _08307_, _24296_);
  nand _48385_ (_16821_, _16820_, _23594_);
  or _48386_ (_16822_, _16820_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _48387_ (_16823_, _16822_, _12774_);
  and _48388_ (_16824_, _16823_, _16821_);
  and _48389_ (_16825_, _08313_, _23642_);
  or _48390_ (_16826_, _16825_, _16824_);
  and _48391_ (_07565_, _16826_, _22762_);
  and _48392_ (_16827_, _16349_, _23649_);
  and _48393_ (_16828_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  or _48394_ (_07567_, _16828_, _16827_);
  and _48395_ (_16829_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  and _48396_ (_16830_, _15991_, _23707_);
  or _48397_ (_07569_, _16830_, _16829_);
  not _48398_ (_16831_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _48399_ (_16832_, _01999_, _16831_);
  or _48400_ (_16833_, _16832_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _48401_ (_16834_, _16833_, _08307_);
  nand _48402_ (_16835_, _05826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _48403_ (_16836_, _16835_, _08307_);
  or _48404_ (_16837_, _16836_, _05827_);
  and _48405_ (_16838_, _16837_, _16834_);
  or _48406_ (_16839_, _16838_, _08313_);
  or _48407_ (_16840_, _12774_, _24043_);
  and _48408_ (_16841_, _16840_, _22762_);
  and _48409_ (_07571_, _16841_, _16839_);
  and _48410_ (_16842_, _08307_, _24125_);
  nand _48411_ (_16843_, _16842_, _23594_);
  or _48412_ (_16844_, _16842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _48413_ (_16845_, _16844_, _12774_);
  and _48414_ (_16846_, _16845_, _16843_);
  and _48415_ (_16847_, _08313_, _23939_);
  or _48416_ (_16848_, _16847_, _16846_);
  and _48417_ (_07573_, _16848_, _22762_);
  and _48418_ (_16849_, _08307_, _24118_);
  nand _48419_ (_16850_, _16849_, _23594_);
  or _48420_ (_16851_, _16849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _48421_ (_16852_, _16851_, _12774_);
  and _48422_ (_16853_, _16852_, _16850_);
  and _48423_ (_16854_, _08313_, _23738_);
  or _48424_ (_16855_, _16854_, _16853_);
  and _48425_ (_07575_, _16855_, _22762_);
  and _48426_ (_16856_, _24050_, _24006_);
  and _48427_ (_16857_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  or _48428_ (_07579_, _16857_, _16856_);
  and _48429_ (_16858_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and _48430_ (_16859_, _16748_, _24050_);
  or _48431_ (_26960_, _16859_, _16858_);
  and _48432_ (_16860_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and _48433_ (_16861_, _16748_, _23778_);
  or _48434_ (_07587_, _16861_, _16860_);
  and _48435_ (_16862_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _48436_ (_16863_, _16862_, _02041_);
  and _48437_ (_16864_, _02009_, _01988_);
  or _48438_ (_16865_, _16864_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _48439_ (_16866_, _16865_, _12758_);
  or _48440_ (_16867_, _16866_, _02001_);
  or _48441_ (_16868_, _16867_, _16863_);
  nor _48442_ (_16869_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _48443_ (_16870_, _16869_, _12764_);
  and _48444_ (_16871_, _16870_, _16868_);
  and _48445_ (_16872_, _01978_, _23892_);
  and _48446_ (_16873_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _48447_ (_16874_, _16873_, _16872_);
  or _48448_ (_16875_, _16874_, _16871_);
  and _48449_ (_07593_, _16875_, _22762_);
  and _48450_ (_16876_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _48451_ (_16877_, _16876_, _02041_);
  and _48452_ (_16878_, _02009_, _01987_);
  nor _48453_ (_16879_, _16878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor _48454_ (_16880_, _16879_, _16864_);
  or _48455_ (_16881_, _16880_, _02001_);
  or _48456_ (_16882_, _16881_, _16877_);
  or _48457_ (_16883_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _48458_ (_16884_, _16883_, _01979_);
  and _48459_ (_16885_, _16884_, _16882_);
  and _48460_ (_16886_, _01978_, _24685_);
  and _48461_ (_16887_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or _48462_ (_16888_, _16887_, _16886_);
  or _48463_ (_16889_, _16888_, _16885_);
  and _48464_ (_07596_, _16889_, _22762_);
  and _48465_ (_16890_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  and _48466_ (_16891_, _16752_, _23946_);
  or _48467_ (_07598_, _16891_, _16890_);
  and _48468_ (_16892_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  and _48469_ (_16893_, _16752_, _23778_);
  or _48470_ (_07602_, _16893_, _16892_);
  and _48471_ (_16894_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  and _48472_ (_16895_, _16758_, _23946_);
  or _48473_ (_07604_, _16895_, _16894_);
  and _48474_ (_16896_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  and _48475_ (_16897_, _16758_, _23898_);
  or _48476_ (_07607_, _16897_, _16896_);
  nor _48477_ (_16898_, _02025_, _12687_);
  nand _48478_ (_16899_, _16898_, _02041_);
  and _48479_ (_16900_, _02009_, _01992_);
  and _48480_ (_16901_, _16900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _48481_ (_16902_, _16900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _48482_ (_16903_, _16902_, _16901_);
  and _48483_ (_16904_, _16903_, _02002_);
  nand _48484_ (_16905_, _16904_, _16899_);
  nand _48485_ (_16906_, _02001_, _12687_);
  and _48486_ (_16907_, _16906_, _01979_);
  and _48487_ (_16908_, _16907_, _16905_);
  and _48488_ (_16909_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _48489_ (_16910_, _16909_, _16908_);
  and _48490_ (_16911_, _01978_, _23642_);
  or _48491_ (_16912_, _16911_, _16910_);
  and _48492_ (_07609_, _16912_, _22762_);
  and _48493_ (_16913_, _06651_, _23747_);
  and _48494_ (_16914_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  or _48495_ (_07611_, _16914_, _16913_);
  and _48496_ (_16915_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and _48497_ (_16916_, _16766_, _24050_);
  or _48498_ (_07614_, _16916_, _16915_);
  and _48499_ (_16917_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and _48500_ (_16918_, _16299_, _24050_);
  or _48501_ (_07617_, _16918_, _16917_);
  nor _48502_ (_16919_, _02018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _48503_ (_16920_, _16919_, _02019_);
  not _48504_ (_16921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor _48505_ (_16922_, _02025_, _16921_);
  nand _48506_ (_16923_, _16922_, _02041_);
  and _48507_ (_16924_, _16923_, _02002_);
  nand _48508_ (_16925_, _16924_, _16920_);
  nand _48509_ (_16926_, _02001_, _16921_);
  and _48510_ (_16927_, _16926_, _01979_);
  and _48511_ (_16928_, _16927_, _16925_);
  and _48512_ (_16929_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _48513_ (_16930_, _16929_, _16928_);
  and _48514_ (_16931_, _01978_, _24043_);
  or _48515_ (_16932_, _16931_, _16930_);
  and _48516_ (_07620_, _16932_, _22762_);
  and _48517_ (_16933_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor _48518_ (_16934_, _16901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor _48519_ (_16935_, _16934_, _02018_);
  and _48520_ (_16936_, _02026_, _02009_);
  and _48521_ (_16937_, _16936_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _48522_ (_16938_, _16937_, _01996_);
  or _48523_ (_16939_, _16938_, _02001_);
  or _48524_ (_16940_, _16939_, _16935_);
  or _48525_ (_16941_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _48526_ (_16942_, _16941_, _01979_);
  and _48527_ (_16943_, _16942_, _16940_);
  or _48528_ (_16944_, _16943_, _16933_);
  and _48529_ (_16945_, _01978_, _23939_);
  or _48530_ (_16946_, _16945_, _16944_);
  and _48531_ (_07622_, _16946_, _22762_);
  and _48532_ (_16947_, _16349_, _23707_);
  and _48533_ (_16948_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  or _48534_ (_07625_, _16948_, _16947_);
  and _48535_ (_16949_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and _48536_ (_16950_, _16772_, _23898_);
  or _48537_ (_07627_, _16950_, _16949_);
  not _48538_ (_16951_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor _48539_ (_16952_, _02025_, _16951_);
  nand _48540_ (_16953_, _16952_, _02041_);
  and _48541_ (_16954_, _02009_, _01990_);
  nor _48542_ (_16955_, _16954_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _48543_ (_16956_, _16955_, _16900_);
  and _48544_ (_16957_, _16956_, _02002_);
  nand _48545_ (_16958_, _16957_, _16953_);
  and _48546_ (_16959_, _02001_, _16951_);
  nor _48547_ (_16960_, _16959_, _12764_);
  and _48548_ (_16961_, _16960_, _16958_);
  and _48549_ (_16962_, _01977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _48550_ (_16963_, _16962_, _16961_);
  and _48551_ (_16964_, _01978_, _23738_);
  or _48552_ (_16965_, _16964_, _16963_);
  and _48553_ (_07630_, _16965_, _22762_);
  and _48554_ (_16966_, _06651_, _23824_);
  and _48555_ (_16967_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  or _48556_ (_07633_, _16967_, _16966_);
  and _48557_ (_16968_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and _48558_ (_16969_, _16780_, _23747_);
  or _48559_ (_07635_, _16969_, _16968_);
  and _48560_ (_16970_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and _48561_ (_16971_, _16299_, _23946_);
  or _48562_ (_07638_, _16971_, _16970_);
  and _48563_ (_16972_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and _48564_ (_16973_, _16299_, _23649_);
  or _48565_ (_07640_, _16973_, _16972_);
  and _48566_ (_16974_, _16349_, _23824_);
  and _48567_ (_16975_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  or _48568_ (_07644_, _16975_, _16974_);
  and _48569_ (_16976_, _01977_, _23738_);
  and _48570_ (_16977_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _48571_ (_16978_, _16977_, _02041_);
  and _48572_ (_16979_, _02009_, _01982_);
  or _48573_ (_16980_, _16979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _48574_ (_16981_, _16980_, _12742_);
  or _48575_ (_16982_, _16981_, _02001_);
  or _48576_ (_16983_, _16982_, _16978_);
  or _48577_ (_16984_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _48578_ (_16985_, _16984_, _01979_);
  and _48579_ (_16986_, _16985_, _16983_);
  and _48580_ (_16987_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _48581_ (_16988_, _16987_, _16986_);
  or _48582_ (_16989_, _16988_, _16976_);
  and _48583_ (_07646_, _16989_, _22762_);
  and _48584_ (_16990_, _01977_, _23816_);
  and _48585_ (_16991_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _48586_ (_16992_, _16991_, _02041_);
  not _48587_ (_16993_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nand _48588_ (_16994_, _02009_, _01981_);
  and _48589_ (_16995_, _16994_, _16993_);
  nor _48590_ (_16996_, _16995_, _16979_);
  or _48591_ (_16997_, _16996_, _02001_);
  or _48592_ (_16998_, _16997_, _16992_);
  or _48593_ (_16999_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _48594_ (_17000_, _16999_, _01979_);
  and _48595_ (_17001_, _17000_, _16998_);
  and _48596_ (_17002_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _48597_ (_17003_, _17002_, _17001_);
  or _48598_ (_17004_, _17003_, _16990_);
  and _48599_ (_07651_, _17004_, _22762_);
  and _48600_ (_17005_, _23992_, _23707_);
  and _48601_ (_17006_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or _48602_ (_07654_, _17006_, _17005_);
  and _48603_ (_17007_, _02001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _48604_ (_17008_, _12708_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _48605_ (_17009_, _16994_, _02002_);
  and _48606_ (_17010_, _17009_, _17008_);
  or _48607_ (_17011_, _17010_, _17007_);
  or _48608_ (_17012_, _17011_, _01977_);
  and _48609_ (_17013_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _48610_ (_17014_, _17013_, _16936_);
  and _48611_ (_17015_, _17014_, _01996_);
  or _48612_ (_17016_, _17015_, _17012_);
  or _48613_ (_17017_, _02017_, _23892_);
  and _48614_ (_17018_, _17017_, _17016_);
  or _48615_ (_17019_, _17018_, _01978_);
  not _48616_ (_17020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand _48617_ (_17021_, _01978_, _17020_);
  and _48618_ (_17022_, _17021_, _22762_);
  and _48619_ (_07656_, _17022_, _17019_);
  and _48620_ (_17023_, _06651_, _23898_);
  and _48621_ (_17024_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  or _48622_ (_07658_, _17024_, _17023_);
  and _48623_ (_17025_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  and _48624_ (_17026_, _16048_, _23946_);
  or _48625_ (_07680_, _17026_, _17025_);
  and _48626_ (_17027_, _12782_, _23707_);
  and _48627_ (_17028_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or _48628_ (_07688_, _17028_, _17027_);
  and _48629_ (_17029_, _24086_, _23649_);
  and _48630_ (_17030_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or _48631_ (_07690_, _17030_, _17029_);
  and _48632_ (_17031_, _16600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  and _48633_ (_17032_, _16599_, _23778_);
  or _48634_ (_07694_, _17032_, _17031_);
  and _48635_ (_17033_, _01977_, _24043_);
  and _48636_ (_17034_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _48637_ (_17035_, _17034_, _02041_);
  and _48638_ (_17036_, _02009_, _01985_);
  nor _48639_ (_17037_, _17036_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _48640_ (_17038_, _17037_, _02043_);
  or _48641_ (_17039_, _17038_, _02001_);
  or _48642_ (_17040_, _17039_, _17035_);
  or _48643_ (_17041_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _48644_ (_17042_, _17041_, _01979_);
  and _48645_ (_17043_, _17042_, _17040_);
  and _48646_ (_17044_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _48647_ (_17045_, _17044_, _17043_);
  or _48648_ (_17046_, _17045_, _17033_);
  and _48649_ (_07697_, _17046_, _22762_);
  and _48650_ (_17047_, _01977_, _23939_);
  and _48651_ (_17048_, _02026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _48652_ (_17049_, _17048_, _02041_);
  and _48653_ (_17050_, _02009_, _01984_);
  nor _48654_ (_17051_, _17050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _48655_ (_17052_, _17051_, _17036_);
  or _48656_ (_17053_, _17052_, _02001_);
  or _48657_ (_17054_, _17053_, _17049_);
  or _48658_ (_17055_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _48659_ (_17056_, _17055_, _01979_);
  and _48660_ (_17057_, _17056_, _17054_);
  and _48661_ (_17058_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _48662_ (_17059_, _17058_, _17057_);
  or _48663_ (_17060_, _17059_, _17047_);
  and _48664_ (_07699_, _17060_, _22762_);
  and _48665_ (_17061_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and _48666_ (_17062_, _16772_, _23946_);
  or _48667_ (_07702_, _17062_, _17061_);
  nor _48668_ (_26861_[2], _24574_, rst);
  and _48669_ (_17063_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  and _48670_ (_17064_, _15991_, _23824_);
  or _48671_ (_07705_, _17064_, _17063_);
  and _48672_ (_17065_, _02345_, _24050_);
  and _48673_ (_17066_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or _48674_ (_07708_, _17066_, _17065_);
  and _48675_ (_17067_, _16349_, _24050_);
  and _48676_ (_17068_, _16351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  or _48677_ (_07712_, _17068_, _17067_);
  or _48678_ (_17069_, _12675_, _24043_);
  nor _48679_ (_17070_, _02078_, _16921_);
  and _48680_ (_17071_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _48681_ (_17072_, _17071_, _17070_);
  or _48682_ (_17073_, _17072_, _02073_);
  and _48683_ (_17074_, _17073_, _22762_);
  and _48684_ (_07716_, _17074_, _17069_);
  and _48685_ (_17075_, _06511_, _23824_);
  and _48686_ (_17076_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or _48687_ (_07719_, _17076_, _17075_);
  and _48688_ (_17077_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  and _48689_ (_17078_, _16752_, _23898_);
  or _48690_ (_07724_, _17078_, _17077_);
  and _48691_ (_17079_, _06511_, _23898_);
  and _48692_ (_17080_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or _48693_ (_07729_, _17080_, _17079_);
  and _48694_ (_17081_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  and _48695_ (_17082_, _16048_, _24050_);
  or _48696_ (_26947_, _17082_, _17081_);
  and _48697_ (_17083_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and _48698_ (_17084_, _16299_, _23778_);
  or _48699_ (_07739_, _17084_, _17083_);
  and _48700_ (_17085_, _05281_, _23898_);
  and _48701_ (_17086_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or _48702_ (_07741_, _17086_, _17085_);
  and _48703_ (_17087_, _01810_, _23824_);
  and _48704_ (_17088_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or _48705_ (_07744_, _17088_, _17087_);
  and _48706_ (_17089_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and _48707_ (_17090_, _13763_, _23946_);
  or _48708_ (_07746_, _17090_, _17089_);
  and _48709_ (_17091_, _24201_, _23986_);
  not _48710_ (_17092_, _17091_);
  and _48711_ (_17093_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  and _48712_ (_17094_, _17091_, _23707_);
  or _48713_ (_07750_, _17094_, _17093_);
  and _48714_ (_17095_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  and _48715_ (_17096_, _17091_, _23898_);
  or _48716_ (_07752_, _17096_, _17095_);
  and _48717_ (_17097_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  and _48718_ (_17098_, _16303_, _23707_);
  or _48719_ (_07765_, _17098_, _17097_);
  nor _48720_ (_17099_, _02078_, _16951_);
  and _48721_ (_17100_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _48722_ (_17101_, _17100_, _17099_);
  and _48723_ (_17102_, _17101_, _12675_);
  and _48724_ (_17103_, _02073_, _23738_);
  or _48725_ (_17104_, _17103_, _17102_);
  and _48726_ (_07767_, _17104_, _22762_);
  or _48727_ (_17105_, _12675_, _23816_);
  nor _48728_ (_17106_, _02078_, _12754_);
  and _48729_ (_17107_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _48730_ (_17108_, _17107_, _17106_);
  or _48731_ (_17109_, _17108_, _02073_);
  and _48732_ (_17110_, _17109_, _22762_);
  and _48733_ (_07769_, _17110_, _17105_);
  and _48734_ (_17111_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  and _48735_ (_17112_, _02306_, _23747_);
  or _48736_ (_07771_, _17112_, _17111_);
  or _48737_ (_17113_, _12675_, _23892_);
  and _48738_ (_17114_, _17113_, _22762_);
  and _48739_ (_17115_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _48740_ (_17116_, _02079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _48741_ (_17117_, _17116_, _17115_);
  or _48742_ (_17118_, _17117_, _02073_);
  and _48743_ (_07773_, _17118_, _17114_);
  and _48744_ (_17119_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and _48745_ (_17120_, _07492_, _23707_);
  or _48746_ (_07775_, _17120_, _17119_);
  and _48747_ (_17121_, _06511_, _23747_);
  and _48748_ (_17122_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or _48749_ (_07777_, _17122_, _17121_);
  or _48750_ (_17123_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or _48751_ (_17124_, _02079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _48752_ (_17125_, _17124_, _17123_);
  or _48753_ (_17126_, _17125_, _02073_);
  nand _48754_ (_17127_, _02073_, _23772_);
  and _48755_ (_17128_, _17127_, _22762_);
  and _48756_ (_07779_, _17128_, _17126_);
  and _48757_ (_17129_, _06511_, _23946_);
  and _48758_ (_17130_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or _48759_ (_07781_, _17130_, _17129_);
  and _48760_ (_17131_, _06511_, _23649_);
  and _48761_ (_17132_, _06514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or _48762_ (_07797_, _17132_, _17131_);
  and _48763_ (_17133_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  and _48764_ (_17134_, _02298_, _23898_);
  or _48765_ (_07800_, _17134_, _17133_);
  or _48766_ (_17135_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _48767_ (_17136_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _48768_ (_17137_, _17136_, _17135_);
  or _48769_ (_17138_, _17137_, _02077_);
  nand _48770_ (_17139_, _02077_, _23772_);
  and _48771_ (_17140_, _17139_, _17138_);
  or _48772_ (_17141_, _17140_, _02073_);
  or _48773_ (_17142_, _12675_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _48774_ (_17143_, _17142_, _22762_);
  and _48775_ (_07802_, _17143_, _17141_);
  and _48776_ (_17144_, _24693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  and _48777_ (_17145_, _24692_, _23824_);
  or _48778_ (_07805_, _17145_, _17144_);
  and _48779_ (_17146_, _05350_, _23824_);
  and _48780_ (_17147_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  or _48781_ (_07818_, _17147_, _17146_);
  and _48782_ (_17148_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  and _48783_ (_17149_, _01967_, _23747_);
  or _48784_ (_07820_, _17149_, _17148_);
  and _48785_ (_17150_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and _48786_ (_17151_, _16299_, _23824_);
  or _48787_ (_07823_, _17151_, _17150_);
  or _48788_ (_17152_, _12671_, _24043_);
  and _48789_ (_17153_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _48790_ (_17154_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _48791_ (_17155_, _17154_, _17153_);
  or _48792_ (_17156_, _17155_, _02077_);
  and _48793_ (_17157_, _17156_, _12675_);
  and _48794_ (_17158_, _17157_, _17152_);
  and _48795_ (_17159_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _48796_ (_17160_, _17159_, _17158_);
  and _48797_ (_07828_, _17160_, _22762_);
  or _48798_ (_17161_, _12671_, _23939_);
  and _48799_ (_17162_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _48800_ (_17163_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _48801_ (_17164_, _17163_, _17162_);
  or _48802_ (_17165_, _17164_, _02077_);
  and _48803_ (_17166_, _17165_, _12675_);
  and _48804_ (_17167_, _17166_, _17161_);
  and _48805_ (_17168_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _48806_ (_17169_, _17168_, _17167_);
  and _48807_ (_07830_, _17169_, _22762_);
  or _48808_ (_17170_, _12671_, _23642_);
  and _48809_ (_17171_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _48810_ (_17172_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _48811_ (_17173_, _17172_, _17171_);
  or _48812_ (_17174_, _17173_, _02077_);
  and _48813_ (_17175_, _17174_, _12675_);
  and _48814_ (_17176_, _17175_, _17170_);
  and _48815_ (_17177_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _48816_ (_17178_, _17177_, _17176_);
  and _48817_ (_07832_, _17178_, _22762_);
  or _48818_ (_17179_, _12671_, _23738_);
  and _48819_ (_17180_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _48820_ (_17181_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _48821_ (_17182_, _17181_, _17180_);
  or _48822_ (_17183_, _17182_, _02077_);
  and _48823_ (_17184_, _17183_, _12675_);
  and _48824_ (_17185_, _17184_, _17179_);
  and _48825_ (_17186_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _48826_ (_17187_, _17186_, _17185_);
  and _48827_ (_07834_, _17187_, _22762_);
  or _48828_ (_17188_, _12671_, _23816_);
  and _48829_ (_17189_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _48830_ (_17190_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _48831_ (_17191_, _17190_, _17189_);
  or _48832_ (_17192_, _17191_, _02077_);
  and _48833_ (_17193_, _17192_, _12675_);
  and _48834_ (_17194_, _17193_, _17188_);
  and _48835_ (_17195_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _48836_ (_17196_, _17195_, _17194_);
  and _48837_ (_07838_, _17196_, _22762_);
  and _48838_ (_17197_, _16300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and _48839_ (_17198_, _16299_, _23898_);
  or _48840_ (_07851_, _17198_, _17197_);
  and _48841_ (_17199_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  and _48842_ (_17200_, _08351_, _23898_);
  or _48843_ (_07854_, _17200_, _17199_);
  and _48844_ (_17201_, _24331_, _23824_);
  and _48845_ (_17202_, _24333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or _48846_ (_08089_, _17202_, _17201_);
  and _48847_ (_17203_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  and _48848_ (_17204_, _15895_, _23747_);
  or _48849_ (_08090_, _17204_, _17203_);
  and _48850_ (_17205_, _06517_, _23649_);
  and _48851_ (_17206_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or _48852_ (_08092_, _17206_, _17205_);
  and _48853_ (_17207_, _24275_, _23076_);
  and _48854_ (_17208_, _17207_, _23824_);
  not _48855_ (_17209_, _17207_);
  and _48856_ (_17210_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or _48857_ (_08094_, _17210_, _17208_);
  and _48858_ (_17211_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  and _48859_ (_17212_, _16303_, _23824_);
  or _48860_ (_08100_, _17212_, _17211_);
  and _48861_ (_17213_, _06517_, _23747_);
  and _48862_ (_17214_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or _48863_ (_08103_, _17214_, _17213_);
  and _48864_ (_17215_, _23903_, _23076_);
  and _48865_ (_17216_, _17215_, _23946_);
  not _48866_ (_17217_, _17215_);
  and _48867_ (_17218_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  or _48868_ (_08107_, _17218_, _17216_);
  and _48869_ (_17219_, _25733_, _23707_);
  and _48870_ (_17220_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or _48871_ (_08110_, _17220_, _17219_);
  and _48872_ (_17221_, _24085_, _23076_);
  and _48873_ (_17222_, _17221_, _23649_);
  not _48874_ (_17223_, _17221_);
  and _48875_ (_17224_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or _48876_ (_08115_, _17224_, _17222_);
  and _48877_ (_17225_, _06517_, _23707_);
  and _48878_ (_17226_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or _48879_ (_08118_, _17226_, _17225_);
  and _48880_ (_17227_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and _48881_ (_17228_, _16780_, _23898_);
  or _48882_ (_08162_, _17228_, _17227_);
  and _48883_ (_17229_, _25078_, _23076_);
  and _48884_ (_17230_, _17229_, _23707_);
  not _48885_ (_17231_, _17229_);
  and _48886_ (_17232_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or _48887_ (_27207_, _17232_, _17230_);
  and _48888_ (_17233_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and _48889_ (_17234_, _16780_, _23824_);
  or _48890_ (_08170_, _17234_, _17233_);
  and _48891_ (_17235_, _16022_, _23707_);
  and _48892_ (_17236_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or _48893_ (_27195_, _17236_, _17235_);
  and _48894_ (_17237_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and _48895_ (_17238_, _16780_, _23649_);
  or _48896_ (_08172_, _17238_, _17237_);
  and _48897_ (_17239_, _05119_, _23898_);
  and _48898_ (_17240_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  or _48899_ (_08175_, _17240_, _17239_);
  and _48900_ (_17241_, _02345_, _23649_);
  and _48901_ (_17242_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or _48902_ (_08179_, _17242_, _17241_);
  and _48903_ (_17243_, _24699_, _23707_);
  and _48904_ (_17244_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  or _48905_ (_08181_, _17244_, _17243_);
  and _48906_ (_17245_, _24283_, _23649_);
  and _48907_ (_17246_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  or _48908_ (_08183_, _17246_, _17245_);
  and _48909_ (_17247_, _25649_, _23824_);
  and _48910_ (_17248_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or _48911_ (_08188_, _17248_, _17247_);
  and _48912_ (_17249_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  and _48913_ (_17250_, _24222_, _23747_);
  or _48914_ (_08190_, _17250_, _17249_);
  and _48915_ (_17251_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  and _48916_ (_17252_, _05193_, _24050_);
  or _48917_ (_08195_, _17252_, _17251_);
  and _48918_ (_17253_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and _48919_ (_17254_, _16780_, _23946_);
  or _48920_ (_26945_, _17254_, _17253_);
  and _48921_ (_17255_, _23784_, _23076_);
  not _48922_ (_17256_, _17255_);
  and _48923_ (_17257_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and _48924_ (_17258_, _17255_, _23778_);
  or _48925_ (_08202_, _17258_, _17257_);
  and _48926_ (_17259_, _24371_, _24050_);
  and _48927_ (_17260_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or _48928_ (_08203_, _17260_, _17259_);
  and _48929_ (_17261_, _16022_, _23747_);
  and _48930_ (_17262_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or _48931_ (_08205_, _17262_, _17261_);
  and _48932_ (_17263_, _24370_, _23986_);
  and _48933_ (_17264_, _17263_, _23824_);
  not _48934_ (_17265_, _17263_);
  and _48935_ (_17266_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  or _48936_ (_08208_, _17266_, _17264_);
  and _48937_ (_17268_, _25656_, _23778_);
  and _48938_ (_17269_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or _48939_ (_08210_, _17269_, _17268_);
  and _48940_ (_17270_, _04922_, _23747_);
  and _48941_ (_17271_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  or _48942_ (_08215_, _17271_, _17270_);
  and _48943_ (_17272_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  and _48944_ (_17273_, _16303_, _23946_);
  or _48945_ (_08421_, _17273_, _17272_);
  and _48946_ (_17274_, _16304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  and _48947_ (_17275_, _16303_, _23649_);
  or _48948_ (_08424_, _17275_, _17274_);
  and _48949_ (_17276_, _02299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  and _48950_ (_17277_, _02298_, _23824_);
  or _48951_ (_08427_, _17277_, _17276_);
  and _48952_ (_17278_, _06517_, _24050_);
  and _48953_ (_17279_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or _48954_ (_08429_, _17279_, _17278_);
  and _48955_ (_17280_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  and _48956_ (_17281_, _15895_, _23649_);
  or _48957_ (_08432_, _17281_, _17280_);
  and _48958_ (_17282_, _17215_, _24050_);
  and _48959_ (_17283_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  or _48960_ (_08435_, _17283_, _17282_);
  and _48961_ (_17284_, _15850_, _23898_);
  and _48962_ (_17285_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  or _48963_ (_08439_, _17285_, _17284_);
  and _48964_ (_17286_, _05119_, _23824_);
  and _48965_ (_17287_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  or _48966_ (_08442_, _17287_, _17286_);
  and _48967_ (_17288_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and _48968_ (_17289_, _16307_, _23946_);
  or _48969_ (_08449_, _17289_, _17288_);
  and _48970_ (_17290_, _24283_, _23946_);
  and _48971_ (_17291_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  or _48972_ (_08451_, _17291_, _17290_);
  and _48973_ (_17292_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and _48974_ (_17293_, _16307_, _23649_);
  or _48975_ (_08454_, _17293_, _17292_);
  and _48976_ (_17295_, _06524_, _23707_);
  and _48977_ (_17296_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  or _48978_ (_08458_, _17296_, _17295_);
  and _48979_ (_17297_, _06524_, _24050_);
  and _48980_ (_17298_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  or _48981_ (_08463_, _17298_, _17297_);
  and _48982_ (_17299_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  and _48983_ (_17300_, _24222_, _23649_);
  or _48984_ (_27246_, _17300_, _17299_);
  and _48985_ (_17301_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  and _48986_ (_17302_, _15895_, _23946_);
  or _48987_ (_08476_, _17302_, _17301_);
  and _48988_ (_17303_, _02374_, _23898_);
  and _48989_ (_17304_, _02376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  or _48990_ (_08487_, _17304_, _17303_);
  or _48991_ (_17305_, _06686_, _03323_);
  or _48992_ (_17306_, _17305_, _06726_);
  or _48993_ (_17307_, _04938_, _24608_);
  or _48994_ (_17308_, _03274_, _26626_);
  or _48995_ (_17309_, _17308_, _17307_);
  or _48996_ (_17310_, _17309_, _04244_);
  or _48997_ (_17311_, _17310_, _17306_);
  or _48998_ (_17312_, _17311_, _03320_);
  and _48999_ (_17313_, _17312_, _22768_);
  and _49000_ (_17314_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or _49001_ (_17315_, _17314_, _03336_);
  or _49002_ (_17316_, _17315_, _17313_);
  and _49003_ (_26873_, _17316_, _22762_);
  and _49004_ (_17317_, _25618_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and _49005_ (_17318_, _24613_, _24606_);
  or _49006_ (_17319_, _17318_, _26635_);
  or _49007_ (_17320_, _17319_, _06719_);
  or _49008_ (_17321_, _05079_, _25633_);
  or _49009_ (_17322_, _05065_, _05088_);
  or _49010_ (_17323_, _17322_, _17321_);
  or _49011_ (_17324_, _17323_, _17320_);
  and _49012_ (_17325_, _17324_, _25644_);
  or _49013_ (_26870_[1], _17325_, _17317_);
  and _49014_ (_17326_, _25618_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or _49015_ (_17327_, _03275_, _26641_);
  or _49016_ (_17328_, _17327_, _12858_);
  or _49017_ (_17329_, _17328_, _26653_);
  or _49018_ (_17330_, _17329_, _02255_);
  or _49019_ (_17331_, _04962_, _02263_);
  or _49020_ (_17332_, _06686_, _06079_);
  or _49021_ (_17333_, _17332_, _17331_);
  or _49022_ (_17334_, _17333_, _06576_);
  or _49023_ (_17335_, _17334_, _17330_);
  or _49024_ (_17336_, _17335_, _06696_);
  and _49025_ (_17337_, _17336_, _25644_);
  or _49026_ (_26871_[3], _17337_, _17326_);
  and _49027_ (_17338_, _02370_, _23747_);
  and _49028_ (_17339_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or _49029_ (_08522_, _17339_, _17338_);
  or _49030_ (_17340_, _03331_, _26572_);
  or _49031_ (_17341_, _03330_, _25636_);
  and _49032_ (_17342_, _17341_, _22766_);
  and _49033_ (_17343_, _17342_, _17340_);
  and _49034_ (_17344_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _49035_ (_17345_, _17344_, _05003_);
  or _49036_ (_17346_, _17345_, _17343_);
  and _49037_ (_26869_[2], _17346_, _22762_);
  or _49038_ (_17347_, _06870_, _04945_);
  and _49039_ (_17348_, _17347_, _22768_);
  and _49040_ (_17349_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _49041_ (_17350_, _17349_, _24570_);
  or _49042_ (_17351_, _17350_, _17348_);
  and _49043_ (_26872_[1], _17351_, _22762_);
  and _49044_ (_17352_, _02370_, _23649_);
  and _49045_ (_17353_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or _49046_ (_08526_, _17353_, _17352_);
  and _49047_ (_17354_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  and _49048_ (_17355_, _07492_, _23898_);
  or _49049_ (_08538_, _17355_, _17354_);
  and _49050_ (_17356_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and _49051_ (_17357_, _07492_, _23824_);
  or _49052_ (_27240_, _17357_, _17356_);
  and _49053_ (_17358_, _17263_, _23778_);
  and _49054_ (_17359_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  or _49055_ (_27193_, _17359_, _17358_);
  and _49056_ (_17360_, _05281_, _23707_);
  and _49057_ (_17361_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or _49058_ (_08740_, _17361_, _17360_);
  and _49059_ (_17362_, _25656_, _24050_);
  and _49060_ (_17363_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or _49061_ (_08749_, _17363_, _17362_);
  and _49062_ (_17364_, _25656_, _23707_);
  and _49063_ (_17365_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or _49064_ (_08765_, _17365_, _17364_);
  and _49065_ (_17366_, _02370_, _23778_);
  and _49066_ (_17367_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or _49067_ (_08771_, _17367_, _17366_);
  and _49068_ (_17368_, _05281_, _24050_);
  and _49069_ (_17369_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or _49070_ (_08773_, _17369_, _17368_);
  and _49071_ (_17370_, _25739_, _23778_);
  and _49072_ (_17371_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  or _49073_ (_27068_, _17371_, _17370_);
  and _49074_ (_17372_, _25739_, _23898_);
  and _49075_ (_17373_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  or _49076_ (_08826_, _17373_, _17372_);
  and _49077_ (_17374_, _25739_, _23824_);
  and _49078_ (_17375_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  or _49079_ (_08828_, _17375_, _17374_);
  and _49080_ (_17376_, _06524_, _23946_);
  and _49081_ (_17377_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  or _49082_ (_08882_, _17377_, _17376_);
  and _49083_ (_17378_, _23991_, _23789_);
  and _49084_ (_17379_, _17378_, _23778_);
  not _49085_ (_17380_, _17378_);
  and _49086_ (_17381_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  or _49087_ (_27289_, _17381_, _17379_);
  and _49088_ (_17382_, _17263_, _23747_);
  and _49089_ (_17383_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  or _49090_ (_08909_, _17383_, _17382_);
  and _49091_ (_17384_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  and _49092_ (_17385_, _07492_, _23747_);
  or _49093_ (_08931_, _17385_, _17384_);
  and _49094_ (_17386_, _12782_, _24050_);
  and _49095_ (_17387_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or _49096_ (_08939_, _17387_, _17386_);
  and _49097_ (_17388_, _23656_, _23076_);
  and _49098_ (_17389_, _17388_, _24050_);
  not _49099_ (_17390_, _17388_);
  and _49100_ (_17391_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or _49101_ (_08943_, _17391_, _17389_);
  and _49102_ (_17392_, _04922_, _23946_);
  and _49103_ (_17393_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  or _49104_ (_08947_, _17393_, _17392_);
  and _49105_ (_17394_, _04922_, _23649_);
  and _49106_ (_17395_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  or _49107_ (_08951_, _17395_, _17394_);
  and _49108_ (_17396_, _23903_, _23789_);
  and _49109_ (_17397_, _17396_, _23649_);
  not _49110_ (_17398_, _17396_);
  and _49111_ (_17399_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  or _49112_ (_08959_, _17399_, _17397_);
  and _49113_ (_17400_, _17396_, _23898_);
  and _49114_ (_17401_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  or _49115_ (_08963_, _17401_, _17400_);
  and _49116_ (_17402_, _16781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and _49117_ (_17403_, _16780_, _23707_);
  or _49118_ (_08965_, _17403_, _17402_);
  and _49119_ (_17404_, _24005_, _23789_);
  and _49120_ (_17405_, _17404_, _23649_);
  not _49121_ (_17406_, _17404_);
  and _49122_ (_17407_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or _49123_ (_08969_, _17407_, _17405_);
  and _49124_ (_17408_, _17404_, _23824_);
  and _49125_ (_17409_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or _49126_ (_08971_, _17409_, _17408_);
  and _49127_ (_17410_, _23986_, _23789_);
  and _49128_ (_17411_, _17410_, _23946_);
  not _49129_ (_17412_, _17410_);
  and _49130_ (_17413_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or _49131_ (_08975_, _17413_, _17411_);
  and _49132_ (_17414_, _17410_, _23747_);
  and _49133_ (_17415_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or _49134_ (_08977_, _17415_, _17414_);
  and _49135_ (_17416_, _23789_, _23069_);
  and _49136_ (_17418_, _17416_, _23946_);
  not _49137_ (_17419_, _17416_);
  and _49138_ (_17420_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  or _49139_ (_08981_, _17420_, _17418_);
  and _49140_ (_17421_, _17416_, _23747_);
  and _49141_ (_17422_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  or _49142_ (_08983_, _17422_, _17421_);
  and _49143_ (_17423_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and _49144_ (_17424_, _16307_, _23707_);
  or _49145_ (_26986_, _17424_, _17423_);
  and _49146_ (_17425_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and _49147_ (_17426_, _16307_, _24050_);
  or _49148_ (_08988_, _17426_, _17425_);
  and _49149_ (_17427_, _17388_, _23946_);
  and _49150_ (_17428_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or _49151_ (_08995_, _17428_, _17427_);
  and _49152_ (_17429_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  and _49153_ (_17430_, _15895_, _23898_);
  or _49154_ (_09002_, _17430_, _17429_);
  and _49155_ (_17431_, _01808_, _23789_);
  and _49156_ (_17432_, _17431_, _24050_);
  not _49157_ (_17433_, _17431_);
  and _49158_ (_17434_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  or _49159_ (_09010_, _17434_, _17432_);
  and _49160_ (_17435_, _17431_, _23649_);
  and _49161_ (_17436_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  or _49162_ (_09011_, _17436_, _17435_);
  and _49163_ (_17437_, _17431_, _23898_);
  and _49164_ (_17438_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  or _49165_ (_09014_, _17438_, _17437_);
  and _49166_ (_17439_, _24329_, _23789_);
  and _49167_ (_17440_, _17439_, _23707_);
  not _49168_ (_17441_, _17439_);
  and _49169_ (_17442_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or _49170_ (_09018_, _17442_, _17440_);
  and _49171_ (_17443_, _15992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  and _49172_ (_17444_, _15991_, _23778_);
  or _49173_ (_09022_, _17444_, _17443_);
  and _49174_ (_17445_, _17439_, _23747_);
  and _49175_ (_17446_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or _49176_ (_09025_, _17446_, _17445_);
  and _49177_ (_17447_, _25078_, _23789_);
  and _49178_ (_17448_, _17447_, _23707_);
  not _49179_ (_17449_, _17447_);
  and _49180_ (_17450_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or _49181_ (_09035_, _17450_, _17448_);
  and _49182_ (_17451_, _06517_, _23778_);
  and _49183_ (_17452_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or _49184_ (_09038_, _17452_, _17451_);
  and _49185_ (_17453_, _06517_, _23898_);
  and _49186_ (_17454_, _06520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or _49187_ (_27150_, _17454_, _17453_);
  and _49188_ (_17455_, _14956_, _24050_);
  and _49189_ (_17456_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or _49190_ (_09047_, _17456_, _17455_);
  and _49191_ (_17457_, _14956_, _23946_);
  and _49192_ (_17458_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or _49193_ (_09049_, _17458_, _17457_);
  and _49194_ (_17459_, _15850_, _23778_);
  and _49195_ (_17460_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  or _49196_ (_27209_, _17460_, _17459_);
  and _49197_ (_17461_, _15896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  and _49198_ (_17462_, _15895_, _23824_);
  or _49199_ (_09059_, _17462_, _17461_);
  and _49200_ (_17463_, _12733_, _23747_);
  and _49201_ (_17464_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  or _49202_ (_09061_, _17464_, _17463_);
  and _49203_ (_17465_, _17447_, _23778_);
  and _49204_ (_17466_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or _49205_ (_09071_, _17466_, _17465_);
  and _49206_ (_17467_, _24282_, _23789_);
  and _49207_ (_17468_, _17467_, _23707_);
  not _49208_ (_17469_, _17467_);
  and _49209_ (_17470_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  or _49210_ (_09074_, _17470_, _17468_);
  and _49211_ (_17471_, _17467_, _23946_);
  and _49212_ (_17472_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or _49213_ (_09075_, _17472_, _17471_);
  and _49214_ (_17473_, _17467_, _23898_);
  and _49215_ (_17474_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  or _49216_ (_09079_, _17474_, _17473_);
  and _49217_ (_17475_, _23789_, _23752_);
  and _49218_ (_17476_, _17475_, _23946_);
  not _49219_ (_17477_, _17475_);
  and _49220_ (_17478_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or _49221_ (_09086_, _17478_, _17476_);
  and _49222_ (_17479_, _23789_, _23656_);
  and _49223_ (_17480_, _17479_, _24050_);
  not _49224_ (_17481_, _17479_);
  and _49225_ (_17482_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or _49226_ (_27273_, _17482_, _17480_);
  and _49227_ (_17483_, _17378_, _23824_);
  and _49228_ (_17484_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  or _49229_ (_09094_, _17484_, _17483_);
  and _49230_ (_17485_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and _49231_ (_17486_, _16307_, _23778_);
  or _49232_ (_26985_, _17486_, _17485_);
  and _49233_ (_17487_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and _49234_ (_17488_, _16582_, _23707_);
  or _49235_ (_09101_, _17488_, _17487_);
  and _49236_ (_17489_, _17404_, _24050_);
  and _49237_ (_17490_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or _49238_ (_09110_, _17490_, _17489_);
  and _49239_ (_17491_, _16049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  and _49240_ (_17492_, _16048_, _23707_);
  or _49241_ (_09112_, _17492_, _17491_);
  and _49242_ (_17493_, _17410_, _23707_);
  and _49243_ (_17494_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or _49244_ (_09114_, _17494_, _17493_);
  and _49245_ (_17495_, _17416_, _23707_);
  and _49246_ (_17496_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  or _49247_ (_09118_, _17496_, _17495_);
  and _49248_ (_17497_, _02370_, _24050_);
  and _49249_ (_17498_, _02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or _49250_ (_09140_, _17498_, _17497_);
  and _49251_ (_17499_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and _49252_ (_17500_, _16772_, _23778_);
  or _49253_ (_09167_, _17500_, _17499_);
  and _49254_ (_17501_, _17479_, _23824_);
  and _49255_ (_17502_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or _49256_ (_09172_, _17502_, _17501_);
  and _49257_ (_17503_, _17447_, _23649_);
  and _49258_ (_17504_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or _49259_ (_09174_, _17504_, _17503_);
  and _49260_ (_17505_, _17475_, _23707_);
  and _49261_ (_17506_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  or _49262_ (_09179_, _17506_, _17505_);
  and _49263_ (_17507_, _17221_, _24050_);
  and _49264_ (_17508_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or _49265_ (_09184_, _17508_, _17507_);
  and _49266_ (_17509_, _06524_, _23778_);
  and _49267_ (_17510_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  or _49268_ (_09191_, _17510_, _17509_);
  and _49269_ (_17511_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and _49270_ (_17512_, _16307_, _23824_);
  or _49271_ (_09194_, _17512_, _17511_);
  and _49272_ (_17513_, _10347_, _23898_);
  and _49273_ (_17514_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  or _49274_ (_27125_, _17514_, _17513_);
  and _49275_ (_17515_, _17396_, _23946_);
  and _49276_ (_17516_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or _49277_ (_09202_, _17516_, _17515_);
  and _49278_ (_17517_, _17416_, _23778_);
  and _49279_ (_17518_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  or _49280_ (_09206_, _17518_, _17517_);
  and _49281_ (_17519_, _17447_, _23898_);
  and _49282_ (_17520_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or _49283_ (_09215_, _17520_, _17519_);
  and _49284_ (_17521_, _17475_, _23898_);
  and _49285_ (_17522_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  or _49286_ (_09219_, _17522_, _17521_);
  and _49287_ (_17523_, _06530_, _23707_);
  and _49288_ (_17524_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  or _49289_ (_09225_, _17524_, _17523_);
  and _49290_ (_17525_, _16308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and _49291_ (_17526_, _16307_, _23898_);
  or _49292_ (_09228_, _17526_, _17525_);
  and _49293_ (_17527_, _17388_, _23778_);
  and _49294_ (_17528_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or _49295_ (_09254_, _17528_, _17527_);
  and _49296_ (_17529_, _12782_, _23898_);
  and _49297_ (_17530_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or _49298_ (_27076_, _17530_, _17529_);
  and _49299_ (_17531_, _12782_, _23778_);
  and _49300_ (_17532_, _12784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or _49301_ (_09258_, _17532_, _17531_);
  and _49302_ (_17533_, _17410_, _23778_);
  and _49303_ (_17534_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or _49304_ (_09270_, _17534_, _17533_);
  and _49305_ (_17535_, _23906_, _23069_);
  and _49306_ (_17536_, _17535_, _23946_);
  not _49307_ (_17537_, _17535_);
  and _49308_ (_17538_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or _49309_ (_09274_, _17538_, _17536_);
  and _49310_ (_17539_, _01808_, _23906_);
  and _49311_ (_17540_, _17539_, _23707_);
  not _49312_ (_17541_, _17539_);
  and _49313_ (_17542_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or _49314_ (_26933_, _17542_, _17540_);
  and _49315_ (_17543_, _17539_, _23824_);
  and _49316_ (_17544_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or _49317_ (_09282_, _17544_, _17543_);
  and _49318_ (_17545_, _06530_, _24050_);
  and _49319_ (_17546_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  or _49320_ (_27148_, _17546_, _17545_);
  and _49321_ (_17547_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and _49322_ (_17548_, _16772_, _23824_);
  or _49323_ (_09291_, _17548_, _17547_);
  and _49324_ (_17549_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and _49325_ (_17550_, _16582_, _23824_);
  or _49326_ (_09296_, _17550_, _17549_);
  and _49327_ (_17551_, _23906_, _23752_);
  and _49328_ (_17552_, _17551_, _23707_);
  not _49329_ (_17553_, _17551_);
  and _49330_ (_17554_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or _49331_ (_09299_, _17554_, _17552_);
  and _49332_ (_17555_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _49333_ (_17556_, _17555_, _26154_);
  and _49334_ (_17557_, _17555_, _26154_);
  or _49335_ (_17558_, _17557_, _17556_);
  and _49336_ (_09302_, _17558_, _22762_);
  and _49337_ (_17559_, _17551_, _23649_);
  and _49338_ (_17560_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or _49339_ (_09305_, _17560_, _17559_);
  and _49340_ (_17561_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and _49341_ (_17562_, _16582_, _23898_);
  or _49342_ (_09309_, _17562_, _17561_);
  and _49343_ (_09312_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _22762_);
  and _49344_ (_09315_, _00845_, _22762_);
  and _49345_ (_09317_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _22762_);
  or _49346_ (_17563_, _23599_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _49347_ (_17564_, _17555_, rst);
  and _49348_ (_09321_, _17564_, _17563_);
  and _49349_ (_17565_, _05042_, _23946_);
  and _49350_ (_17566_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or _49351_ (_09327_, _17566_, _17565_);
  and _49352_ (_17567_, _12733_, _23824_);
  and _49353_ (_17568_, _12735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  or _49354_ (_09331_, _17568_, _17567_);
  and _49355_ (_17569_, _23906_, _23656_);
  and _49356_ (_17570_, _17569_, _23946_);
  not _49357_ (_17571_, _17569_);
  and _49358_ (_17572_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  or _49359_ (_09334_, _17572_, _17570_);
  and _49360_ (_17573_, _17569_, _23778_);
  and _49361_ (_17574_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  or _49362_ (_09340_, _17574_, _17573_);
  and _49363_ (_17575_, _25078_, _23906_);
  and _49364_ (_17576_, _17575_, _24050_);
  not _49365_ (_17577_, _17575_);
  and _49366_ (_17578_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  or _49367_ (_09343_, _17578_, _17576_);
  and _49368_ (_17579_, _17575_, _23898_);
  and _49369_ (_17580_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  or _49370_ (_09347_, _17580_, _17579_);
  and _49371_ (_17581_, _24282_, _23906_);
  and _49372_ (_17582_, _17581_, _23707_);
  not _49373_ (_17583_, _17581_);
  and _49374_ (_17584_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or _49375_ (_09350_, _17584_, _17582_);
  and _49376_ (_17585_, _17581_, _23824_);
  and _49377_ (_17586_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or _49378_ (_09354_, _17586_, _17585_);
  and _49379_ (_17587_, _24010_, _23906_);
  and _49380_ (_17588_, _17587_, _23946_);
  not _49381_ (_17589_, _17587_);
  and _49382_ (_17590_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  or _49383_ (_09357_, _17590_, _17588_);
  and _49384_ (_17591_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  and _49385_ (_17592_, _08477_, _23747_);
  or _49386_ (_09359_, _17592_, _17591_);
  and _49387_ (_17593_, _24085_, _23906_);
  and _49388_ (_17594_, _17593_, _23946_);
  not _49389_ (_17595_, _17593_);
  and _49390_ (_17596_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  or _49391_ (_09366_, _17596_, _17594_);
  and _49392_ (_17597_, _17593_, _23824_);
  and _49393_ (_17598_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  or _49394_ (_09368_, _17598_, _17597_);
  and _49395_ (_17599_, _23906_, _23784_);
  and _49396_ (_17601_, _17599_, _23707_);
  not _49397_ (_17602_, _17599_);
  and _49398_ (_17603_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or _49399_ (_09370_, _17603_, _17601_);
  and _49400_ (_17604_, _17599_, _23649_);
  and _49401_ (_17605_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or _49402_ (_09373_, _17605_, _17604_);
  and _49403_ (_17606_, _17599_, _23778_);
  and _49404_ (_17607_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or _49405_ (_09375_, _17607_, _17606_);
  and _49406_ (_17608_, _23911_, _23906_);
  and _49407_ (_17609_, _17608_, _24050_);
  not _49408_ (_17610_, _17608_);
  and _49409_ (_17611_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or _49410_ (_09379_, _17611_, _17609_);
  and _49411_ (_17612_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and _49412_ (_17613_, _16582_, _23778_);
  or _49413_ (_09382_, _17613_, _17612_);
  and _49414_ (_17614_, _17608_, _23649_);
  and _49415_ (_17615_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or _49416_ (_09384_, _17615_, _17614_);
  and _49417_ (_17616_, _06524_, _23747_);
  and _49418_ (_17617_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  or _49419_ (_09387_, _17617_, _17616_);
  and _49420_ (_17618_, _05350_, _24050_);
  and _49421_ (_17619_, _05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  or _49422_ (_09421_, _17619_, _17618_);
  and _49423_ (_17620_, _05119_, _23707_);
  and _49424_ (_17621_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or _49425_ (_09523_, _17621_, _17620_);
  and _49426_ (_17622_, _25618_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or _49427_ (_17623_, _02256_, _02273_);
  or _49428_ (_17624_, _17623_, _06686_);
  or _49429_ (_17625_, _06697_, _03273_);
  or _49430_ (_17626_, _17625_, _17624_);
  or _49431_ (_17627_, _17626_, _06696_);
  and _49432_ (_17628_, _17627_, _25644_);
  or _49433_ (_26867_[1], _17628_, _17622_);
  and _49434_ (_17629_, _17388_, _23747_);
  and _49435_ (_17630_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or _49436_ (_09600_, _17630_, _17629_);
  and _49437_ (_17631_, _17388_, _23824_);
  and _49438_ (_17632_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or _49439_ (_09612_, _17632_, _17631_);
  and _49440_ (_17633_, _14956_, _23898_);
  and _49441_ (_17634_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or _49442_ (_09626_, _17634_, _17633_);
  and _49443_ (_17635_, _07536_, _23824_);
  and _49444_ (_17636_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  or _49445_ (_09638_, _17636_, _17635_);
  and _49446_ (_17637_, _14956_, _23778_);
  and _49447_ (_17638_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or _49448_ (_09652_, _17638_, _17637_);
  and _49449_ (_17639_, _17229_, _23747_);
  and _49450_ (_17640_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or _49451_ (_09668_, _17640_, _17639_);
  and _49452_ (_17641_, _05281_, _23778_);
  and _49453_ (_17642_, _05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or _49454_ (_09681_, _17642_, _17641_);
  and _49455_ (_17643_, _17229_, _23824_);
  and _49456_ (_17644_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or _49457_ (_27206_, _17644_, _17643_);
  and _49458_ (_17645_, _14956_, _23747_);
  and _49459_ (_17646_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or _49460_ (_09731_, _17646_, _17645_);
  and _49461_ (_17647_, _17229_, _24050_);
  and _49462_ (_17648_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or _49463_ (_09733_, _17648_, _17647_);
  and _49464_ (_17649_, _14956_, _23824_);
  and _49465_ (_17650_, _14958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or _49466_ (_09737_, _17650_, _17649_);
  and _49467_ (_17651_, _17229_, _23946_);
  and _49468_ (_17652_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or _49469_ (_09753_, _17652_, _17651_);
  or _49470_ (_17653_, _04891_, _24043_);
  or _49471_ (_17654_, _05165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _49472_ (_17655_, _05166_, _26098_);
  and _49473_ (_17656_, _17655_, _17654_);
  and _49474_ (_17657_, _07418_, _24310_);
  or _49475_ (_17658_, _17657_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _49476_ (_17659_, _05144_, _04860_);
  and _49477_ (_17660_, _17659_, _17658_);
  or _49478_ (_17661_, _05151_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _49479_ (_17662_, _05152_);
  and _49480_ (_17663_, _17662_, _24302_);
  and _49481_ (_17664_, _17663_, _17661_);
  and _49482_ (_17665_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _49483_ (_17666_, _17665_, _17664_);
  or _49484_ (_17667_, _17666_, _17660_);
  or _49485_ (_17668_, _17667_, _17656_);
  or _49486_ (_17669_, _17668_, _24299_);
  and _49487_ (_17670_, _17669_, _24294_);
  and _49488_ (_17671_, _17670_, _17653_);
  and _49489_ (_17672_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _49490_ (_17673_, _17672_, _17671_);
  and _49491_ (_09769_, _17673_, _22762_);
  and _49492_ (_17674_, _12786_, _23747_);
  and _49493_ (_17675_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  or _49494_ (_09818_, _17675_, _17674_);
  and _49495_ (_17676_, _24283_, _23707_);
  and _49496_ (_17677_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or _49497_ (_09821_, _17677_, _17676_);
  and _49498_ (_17678_, _09913_, _23778_);
  and _49499_ (_17679_, _09915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or _49500_ (_09823_, _17679_, _17678_);
  and _49501_ (_17680_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  and _49502_ (_17681_, _08477_, _23824_);
  or _49503_ (_09837_, _17681_, _17680_);
  and _49504_ (_17682_, _12786_, _23824_);
  and _49505_ (_17683_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  or _49506_ (_09839_, _17683_, _17682_);
  and _49507_ (_17684_, _24283_, _24050_);
  and _49508_ (_17685_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  or _49509_ (_09854_, _17685_, _17684_);
  and _49510_ (_17686_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and _49511_ (_17687_, _01967_, _23824_);
  or _49512_ (_09860_, _17687_, _17686_);
  and _49513_ (_17688_, _12786_, _23898_);
  and _49514_ (_17689_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  or _49515_ (_27075_, _17689_, _17688_);
  and _49516_ (_17690_, _25649_, _24050_);
  and _49517_ (_17691_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or _49518_ (_09887_, _17691_, _17690_);
  and _49519_ (_17692_, _17207_, _23946_);
  and _49520_ (_17693_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or _49521_ (_09900_, _17693_, _17692_);
  and _49522_ (_17694_, _17207_, _23649_);
  and _49523_ (_17695_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or _49524_ (_09906_, _17695_, _17694_);
  and _49525_ (_17696_, _17207_, _23747_);
  and _49526_ (_17697_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or _49527_ (_09919_, _17697_, _17696_);
  and _49528_ (_17698_, _24652_, _24064_);
  nand _49529_ (_17699_, _17698_, _24118_);
  and _49530_ (_17700_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _49531_ (_17701_, _25170_, _24117_);
  and _49532_ (_17702_, _17701_, _24064_);
  and _49533_ (_17703_, _17702_, _24068_);
  and _49534_ (_17704_, _17703_, _22948_);
  and _49535_ (_17705_, _17704_, _00708_);
  or _49536_ (_17706_, _17705_, _17700_);
  or _49537_ (_17707_, _17706_, _06343_);
  not _49538_ (_17708_, _06343_);
  or _49539_ (_17709_, _17708_, _01255_);
  and _49540_ (_17710_, _17709_, _22762_);
  and _49541_ (_09940_, _17710_, _17707_);
  and _49542_ (_17711_, _17535_, _23824_);
  and _49543_ (_17712_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or _49544_ (_09945_, _17712_, _17711_);
  and _49545_ (_17713_, _17539_, _23649_);
  and _49546_ (_17714_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or _49547_ (_09950_, _17714_, _17713_);
  and _49548_ (_17715_, _06524_, _23824_);
  and _49549_ (_17716_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  or _49550_ (_09952_, _17716_, _17715_);
  and _49551_ (_17717_, _17539_, _23778_);
  and _49552_ (_17718_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or _49553_ (_09954_, _17718_, _17717_);
  and _49554_ (_17719_, _24329_, _23906_);
  and _49555_ (_17720_, _17719_, _23747_);
  not _49556_ (_17721_, _17719_);
  and _49557_ (_17722_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  or _49558_ (_09956_, _17722_, _17720_);
  and _49559_ (_17723_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _49560_ (_17724_, _17704_, _00875_);
  or _49561_ (_17725_, _17724_, _17723_);
  or _49562_ (_17726_, _17725_, _06343_);
  or _49563_ (_17727_, _17708_, _04299_);
  and _49564_ (_17728_, _17727_, _22762_);
  and _49565_ (_09964_, _17728_, _17726_);
  and _49566_ (_17729_, _17719_, _23778_);
  and _49567_ (_17730_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  or _49568_ (_09966_, _17730_, _17729_);
  and _49569_ (_17731_, _06524_, _23898_);
  and _49570_ (_17732_, _06527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  or _49571_ (_27149_, _17732_, _17731_);
  and _49572_ (_17733_, _17551_, _23898_);
  and _49573_ (_17734_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or _49574_ (_09974_, _17734_, _17733_);
  and _49575_ (_17735_, _17698_, _24291_);
  nor _49576_ (_17736_, _17735_, _06343_);
  or _49577_ (_17737_, _17736_, _26565_);
  not _49578_ (_17738_, _17736_);
  or _49579_ (_17739_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _49580_ (_17740_, _17739_, _22762_);
  and _49581_ (_09976_, _17740_, _17737_);
  and _49582_ (_17741_, _17569_, _23824_);
  and _49583_ (_17742_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  or _49584_ (_09988_, _17742_, _17741_);
  and _49585_ (_17743_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and _49586_ (_17744_, _16582_, _23946_);
  or _49587_ (_09991_, _17744_, _17743_);
  and _49588_ (_17745_, _17575_, _23747_);
  and _49589_ (_17746_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  or _49590_ (_26918_, _17746_, _17745_);
  or _49591_ (_17747_, _17736_, _00545_);
  or _49592_ (_17748_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _49593_ (_17749_, _17748_, _22762_);
  and _49594_ (_10005_, _17749_, _17747_);
  and _49595_ (_17750_, _17581_, _23649_);
  and _49596_ (_17751_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or _49597_ (_10007_, _17751_, _17750_);
  and _49598_ (_17752_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  and _49599_ (_17753_, _05199_, _23707_);
  or _49600_ (_10013_, _17753_, _17752_);
  and _49601_ (_17754_, _15012_, _23898_);
  and _49602_ (_17755_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or _49603_ (_10021_, _17755_, _17754_);
  and _49604_ (_17756_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and _49605_ (_17757_, _16582_, _23649_);
  or _49606_ (_10036_, _17757_, _17756_);
  and _49607_ (_17758_, _05838_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _49608_ (_17759_, _17758_, _05839_);
  and _49609_ (_17760_, _17759_, _00276_);
  or _49610_ (_17761_, _00277_, _00276_);
  nor _49611_ (_17762_, _17761_, _23594_);
  and _49612_ (_17763_, _00280_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _49613_ (_17764_, _17763_, _25773_);
  or _49614_ (_17765_, _17764_, _17762_);
  or _49615_ (_17766_, _17765_, _17760_);
  nand _49616_ (_17767_, _25777_, _23702_);
  and _49617_ (_17768_, _17767_, _22762_);
  and _49618_ (_10039_, _17768_, _17766_);
  nand _49619_ (_17769_, _17738_, _00793_);
  or _49620_ (_17770_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _49621_ (_17771_, _17770_, _22762_);
  and _49622_ (_10048_, _17771_, _17769_);
  or _49623_ (_17772_, _17736_, _00451_);
  or _49624_ (_17773_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _49625_ (_17774_, _17773_, _22762_);
  and _49626_ (_10050_, _17774_, _17772_);
  and _49627_ (_17775_, _01808_, _24201_);
  not _49628_ (_17776_, _17775_);
  and _49629_ (_17777_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  and _49630_ (_17778_, _17775_, _23778_);
  or _49631_ (_10055_, _17778_, _17777_);
  and _49632_ (_17779_, _17535_, _24050_);
  and _49633_ (_17780_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or _49634_ (_26934_, _17780_, _17779_);
  and _49635_ (_17781_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _49636_ (_17782_, _17704_, _00620_);
  or _49637_ (_17783_, _17782_, _17781_);
  or _49638_ (_17784_, _17783_, _06343_);
  or _49639_ (_17785_, _17708_, _01192_);
  and _49640_ (_17786_, _17785_, _22762_);
  and _49641_ (_10074_, _17786_, _17784_);
  and _49642_ (_17787_, _17551_, _23946_);
  and _49643_ (_17788_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or _49644_ (_10083_, _17788_, _17787_);
  and _49645_ (_17789_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _49646_ (_17790_, _17704_, _00545_);
  or _49647_ (_17791_, _17790_, _17789_);
  or _49648_ (_17792_, _17791_, _06343_);
  nand _49649_ (_17793_, _06343_, _01129_);
  and _49650_ (_17794_, _17793_, _22762_);
  and _49651_ (_10085_, _17794_, _17792_);
  and _49652_ (_17795_, _17569_, _24050_);
  and _49653_ (_17796_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  or _49654_ (_26921_, _17796_, _17795_);
  and _49655_ (_17797_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and _49656_ (_17798_, _16772_, _23747_);
  or _49657_ (_10089_, _17798_, _17797_);
  and _49658_ (_17799_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _49659_ (_17800_, _17704_, _00451_);
  or _49660_ (_17801_, _17800_, _17799_);
  or _49661_ (_17802_, _17801_, _06343_);
  nand _49662_ (_17803_, _06343_, _01061_);
  and _49663_ (_17804_, _17803_, _22762_);
  and _49664_ (_10097_, _17804_, _17802_);
  and _49665_ (_17805_, _17593_, _23747_);
  and _49666_ (_17806_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  or _49667_ (_10100_, _17806_, _17805_);
  and _49668_ (_17807_, _16583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and _49669_ (_17808_, _16582_, _23747_);
  or _49670_ (_10104_, _17808_, _17807_);
  and _49671_ (_17809_, _17581_, _23778_);
  and _49672_ (_17810_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or _49673_ (_10108_, _17810_, _17809_);
  and _49674_ (_17811_, _17608_, _23898_);
  and _49675_ (_17812_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or _49676_ (_10110_, _17812_, _17811_);
  and _49677_ (_17813_, _17575_, _23707_);
  and _49678_ (_17814_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or _49679_ (_10114_, _17814_, _17813_);
  and _49680_ (_17815_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and _49681_ (_17816_, _16772_, _24050_);
  or _49682_ (_26949_, _17816_, _17815_);
  nand _49683_ (_17817_, _17738_, _00372_);
  or _49684_ (_17818_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _49685_ (_17819_, _17818_, _22762_);
  and _49686_ (_10125_, _17819_, _17817_);
  or _49687_ (_17820_, _17736_, _00708_);
  or _49688_ (_17821_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _49689_ (_17822_, _17821_, _22762_);
  and _49690_ (_10128_, _17822_, _17820_);
  or _49691_ (_17823_, _17736_, _00620_);
  or _49692_ (_17824_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _49693_ (_17825_, _17824_, _22762_);
  and _49694_ (_10130_, _17825_, _17823_);
  nor _49695_ (_17826_, _17699_, _00372_);
  and _49696_ (_17827_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _49697_ (_17828_, _17827_, _06343_);
  or _49698_ (_17829_, _17828_, _17826_);
  nand _49699_ (_17830_, _06343_, _00993_);
  and _49700_ (_17831_, _17830_, _22762_);
  and _49701_ (_10132_, _17831_, _17829_);
  and _49702_ (_17832_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _49703_ (_17833_, _17704_, _26565_);
  or _49704_ (_17834_, _17833_, _17832_);
  or _49705_ (_17835_, _17834_, _06343_);
  or _49706_ (_17836_, _17708_, _00930_);
  and _49707_ (_17837_, _17836_, _22762_);
  and _49708_ (_10133_, _17837_, _17835_);
  or _49709_ (_17838_, _17736_, _00875_);
  or _49710_ (_17839_, _17738_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _49711_ (_17840_, _17839_, _22762_);
  and _49712_ (_10143_, _17840_, _17838_);
  and _49713_ (_17841_, _06530_, _23824_);
  and _49714_ (_17842_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  or _49715_ (_10147_, _17842_, _17841_);
  and _49716_ (_17843_, _17608_, _23778_);
  and _49717_ (_17844_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or _49718_ (_27300_, _17844_, _17843_);
  and _49719_ (_17845_, _17475_, _23778_);
  and _49720_ (_17846_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  or _49721_ (_10157_, _17846_, _17845_);
  and _49722_ (_17847_, _25649_, _23707_);
  and _49723_ (_17848_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or _49724_ (_10163_, _17848_, _17847_);
  and _49725_ (_17849_, _25649_, _23946_);
  and _49726_ (_17850_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or _49727_ (_10165_, _17850_, _17849_);
  nor _49728_ (_17851_, _17699_, _00793_);
  and _49729_ (_17852_, _17699_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _49730_ (_17853_, _17852_, _06343_);
  or _49731_ (_17854_, _17853_, _17851_);
  nand _49732_ (_17855_, _06343_, _01318_);
  and _49733_ (_17856_, _17855_, _22762_);
  and _49734_ (_10169_, _17856_, _17854_);
  and _49735_ (_17857_, _17587_, _24050_);
  and _49736_ (_17858_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  or _49737_ (_10172_, _17858_, _17857_);
  and _49738_ (_26861_[1], _26676_, _22762_);
  and _49739_ (_17859_, _17221_, _23707_);
  and _49740_ (_17860_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or _49741_ (_27202_, _17860_, _17859_);
  and _49742_ (_17861_, _06530_, _23747_);
  and _49743_ (_17862_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  or _49744_ (_27146_, _17862_, _17861_);
  and _49745_ (_17863_, _17479_, _23946_);
  and _49746_ (_17864_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or _49747_ (_10179_, _17864_, _17863_);
  and _49748_ (_17865_, _17221_, _23946_);
  and _49749_ (_17866_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or _49750_ (_10182_, _17866_, _17865_);
  and _49751_ (_17867_, _17587_, _23707_);
  and _49752_ (_17868_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  or _49753_ (_27299_, _17868_, _17867_);
  and _49754_ (_17869_, _17479_, _23707_);
  and _49755_ (_17870_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or _49756_ (_27274_, _17870_, _17869_);
  and _49757_ (_17871_, _16773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and _49758_ (_17872_, _16772_, _23707_);
  or _49759_ (_10188_, _17872_, _17871_);
  and _49760_ (_17873_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and _49761_ (_17874_, _16766_, _23778_);
  or _49762_ (_10192_, _17874_, _17873_);
  and _49763_ (_17875_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  and _49764_ (_17876_, _10331_, _23649_);
  or _49765_ (_10194_, _17876_, _17875_);
  and _49766_ (_17877_, _25649_, _23778_);
  and _49767_ (_17878_, _25651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or _49768_ (_10196_, _17878_, _17877_);
  and _49769_ (_17879_, _17608_, _23824_);
  and _49770_ (_17880_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or _49771_ (_10197_, _17880_, _17879_);
  and _49772_ (_17881_, _17475_, _23824_);
  and _49773_ (_17882_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  or _49774_ (_10201_, _17882_, _17881_);
  and _49775_ (_17883_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  and _49776_ (_17884_, _10331_, _23747_);
  or _49777_ (_26983_, _17884_, _17883_);
  and _49778_ (_17885_, _04922_, _23707_);
  and _49779_ (_17886_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  or _49780_ (_10206_, _17886_, _17885_);
  and _49781_ (_17887_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and _49782_ (_17888_, _16766_, _23898_);
  or _49783_ (_26950_, _17888_, _17887_);
  and _49784_ (_17889_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and _49785_ (_17890_, _16766_, _23747_);
  or _49786_ (_10221_, _17890_, _17889_);
  and _49787_ (_17891_, _17475_, _23747_);
  and _49788_ (_17892_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  or _49789_ (_10225_, _17892_, _17891_);
  and _49790_ (_17893_, _24852_, _24050_);
  and _49791_ (_17894_, _24854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  or _49792_ (_10227_, _17894_, _17893_);
  and _49793_ (_17895_, _17608_, _23747_);
  and _49794_ (_17896_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or _49795_ (_10231_, _17896_, _17895_);
  and _49796_ (_17897_, _24283_, _23778_);
  and _49797_ (_17898_, _24285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  or _49798_ (_10239_, _17898_, _17897_);
  and _49799_ (_17899_, _17608_, _23946_);
  and _49800_ (_17900_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or _49801_ (_10240_, _17900_, _17899_);
  and _49802_ (_17901_, _17475_, _23649_);
  and _49803_ (_17902_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  or _49804_ (_10253_, _17902_, _17901_);
  and _49805_ (_17903_, _17608_, _23707_);
  and _49806_ (_17904_, _17610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or _49807_ (_10258_, _17904_, _17903_);
  and _49808_ (_17905_, _17475_, _24050_);
  and _49809_ (_17906_, _17477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  or _49810_ (_10260_, _17906_, _17905_);
  and _49811_ (_17907_, _24050_, _23912_);
  and _49812_ (_17908_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  or _49813_ (_27268_, _17908_, _17907_);
  and _49814_ (_17909_, _24699_, _23747_);
  and _49815_ (_17910_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  or _49816_ (_27190_, _17910_, _17909_);
  and _49817_ (_17911_, _24699_, _23898_);
  and _49818_ (_17912_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  or _49819_ (_10280_, _17912_, _17911_);
  and _49820_ (_17913_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  and _49821_ (_17914_, _10331_, _23946_);
  or _49822_ (_26984_, _17914_, _17913_);
  and _49823_ (_17915_, _17599_, _23898_);
  and _49824_ (_17916_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or _49825_ (_10287_, _17916_, _17915_);
  and _49826_ (_17917_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  and _49827_ (_17918_, _10331_, _23707_);
  or _49828_ (_10289_, _17918_, _17917_);
  and _49829_ (_17919_, _23912_, _23707_);
  and _49830_ (_17920_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or _49831_ (_10293_, _17920_, _17919_);
  and _49832_ (_17921_, _24699_, _23946_);
  and _49833_ (_17922_, _24701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  or _49834_ (_10297_, _17922_, _17921_);
  and _49835_ (_17923_, _17599_, _23824_);
  and _49836_ (_17924_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or _49837_ (_10301_, _17924_, _17923_);
  and _49838_ (_17925_, _10332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  and _49839_ (_17926_, _10331_, _24050_);
  or _49840_ (_10304_, _17926_, _17925_);
  and _49841_ (_17927_, _17467_, _23778_);
  and _49842_ (_17928_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  or _49843_ (_10308_, _17928_, _17927_);
  and _49844_ (_17929_, _02345_, _23898_);
  and _49845_ (_17930_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or _49846_ (_10310_, _17930_, _17929_);
  and _49847_ (_17931_, _17467_, _23824_);
  and _49848_ (_17932_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  or _49849_ (_10314_, _17932_, _17931_);
  and _49850_ (_17933_, _00276_, _24296_);
  nand _49851_ (_17934_, _17933_, _23594_);
  not _49852_ (_17935_, _25777_);
  or _49853_ (_17936_, _17933_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _49854_ (_17937_, _17936_, _17935_);
  and _49855_ (_17938_, _17937_, _17934_);
  or _49856_ (_17939_, _17938_, _25918_);
  and _49857_ (_10317_, _17939_, _22762_);
  and _49858_ (_17940_, _17599_, _23747_);
  and _49859_ (_17941_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or _49860_ (_27295_, _17941_, _17940_);
  and _49861_ (_17942_, _06530_, _23649_);
  and _49862_ (_17943_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  or _49863_ (_27147_, _17943_, _17942_);
  and _49864_ (_17944_, _00276_, _24118_);
  or _49865_ (_17945_, _17944_, _25775_);
  nand _49866_ (_17946_, _17944_, _23594_);
  and _49867_ (_17947_, _17946_, _17945_);
  or _49868_ (_17948_, _17947_, _25779_);
  and _49869_ (_10329_, _17948_, _22762_);
  and _49870_ (_17949_, _00276_, _24125_);
  nand _49871_ (_17950_, _17949_, _23594_);
  or _49872_ (_17951_, _17949_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _49873_ (_17952_, _17951_, _17935_);
  and _49874_ (_17953_, _17952_, _17950_);
  and _49875_ (_17954_, _25777_, _23939_);
  or _49876_ (_17955_, _17954_, _17953_);
  and _49877_ (_10330_, _17955_, _22762_);
  and _49878_ (_17956_, _17599_, _23946_);
  and _49879_ (_17957_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or _49880_ (_27296_, _17957_, _17956_);
  and _49881_ (_17958_, _17467_, _23747_);
  and _49882_ (_17959_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  or _49883_ (_27269_, _17959_, _17958_);
  and _49884_ (_17960_, _25656_, _23747_);
  and _49885_ (_17961_, _25659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or _49886_ (_10336_, _17961_, _17960_);
  or _49887_ (_17962_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _49888_ (_17963_, _00334_, _26541_);
  or _49889_ (_17964_, _17963_, _00428_);
  or _49890_ (_17965_, _17964_, _00511_);
  or _49891_ (_17966_, _17965_, _00600_);
  or _49892_ (_17967_, _17966_, _00679_);
  and _49893_ (_17968_, _17967_, _23596_);
  and _49894_ (_17969_, _23471_, _23143_);
  not _49895_ (_17970_, _23471_);
  and _49896_ (_17971_, _23473_, _17970_);
  or _49897_ (_17972_, _17971_, _17969_);
  and _49898_ (_17973_, _17972_, _23087_);
  nand _49899_ (_17974_, _23516_, _23482_);
  or _49900_ (_17975_, _23516_, _23145_);
  and _49901_ (_17976_, _17975_, _23480_);
  and _49902_ (_17977_, _17976_, _17974_);
  and _49903_ (_17978_, _23599_, _23214_);
  and _49904_ (_17979_, _17978_, _23418_);
  and _49905_ (_17980_, _01112_, _26152_);
  and _49906_ (_17982_, _17980_, _01233_);
  nand _49907_ (_17983_, _17982_, _17979_);
  nand _49908_ (_17984_, _17983_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _49909_ (_17985_, _17984_, _17977_);
  nor _49910_ (_17986_, _17985_, _17973_);
  nand _49911_ (_17987_, _17986_, _00767_);
  or _49912_ (_17988_, _17987_, _17968_);
  or _49913_ (_17989_, _17988_, _00852_);
  and _49914_ (_17990_, _17989_, _17962_);
  or _49915_ (_17991_, _17990_, _00276_);
  and _49916_ (_17992_, _04388_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _49917_ (_17993_, _17992_, _04389_);
  nand _49918_ (_17994_, _17993_, _00276_);
  and _49919_ (_17995_, _17994_, _17991_);
  or _49920_ (_17996_, _17995_, _25777_);
  or _49921_ (_17997_, _17935_, _23816_);
  and _49922_ (_17998_, _17997_, _22762_);
  and _49923_ (_10338_, _17998_, _17996_);
  and _49924_ (_17999_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  and _49925_ (_18000_, _23501_, _23480_);
  and _49926_ (_18001_, _23467_, _23087_);
  or _49927_ (_18002_, _18001_, _18000_);
  and _49928_ (_18003_, _18002_, _17999_);
  not _49929_ (_18004_, _17999_);
  or _49930_ (_18005_, _18004_, _23579_);
  and _49931_ (_18006_, _18005_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _49932_ (_18007_, _18006_, _00276_);
  or _49933_ (_18008_, _18007_, _18003_);
  or _49934_ (_18009_, _24705_, _00527_);
  nand _49935_ (_18010_, _18009_, _00276_);
  or _49936_ (_18011_, _18010_, _05827_);
  and _49937_ (_18012_, _18011_, _18008_);
  or _49938_ (_18013_, _18012_, _25777_);
  or _49939_ (_18014_, _17935_, _24043_);
  and _49940_ (_18015_, _18014_, _22762_);
  and _49941_ (_10341_, _18015_, _18013_);
  and _49942_ (_18016_, _17263_, _23898_);
  and _49943_ (_18017_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  or _49944_ (_10342_, _18017_, _18016_);
  and _49945_ (_18018_, _17599_, _24050_);
  and _49946_ (_18019_, _17602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or _49947_ (_10345_, _18019_, _18018_);
  and _49948_ (_18020_, _17467_, _23649_);
  and _49949_ (_18021_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  or _49950_ (_10346_, _18021_, _18020_);
  and _49951_ (_18022_, _17593_, _23778_);
  and _49952_ (_18023_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  or _49953_ (_10349_, _18023_, _18022_);
  and _49954_ (_10353_, _05850_, _22762_);
  and _49955_ (_18024_, _17263_, _23946_);
  and _49956_ (_18025_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or _49957_ (_10355_, _18025_, _18024_);
  and _49958_ (_26861_[0], _24632_, _22762_);
  and _49959_ (_18026_, _17467_, _24050_);
  and _49960_ (_18027_, _17469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  or _49961_ (_27270_, _18027_, _18026_);
  and _49962_ (_18028_, _17207_, _24050_);
  and _49963_ (_18029_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or _49964_ (_10360_, _18029_, _18028_);
  and _49965_ (_18030_, _00276_, _24067_);
  nand _49966_ (_18031_, _18030_, _23594_);
  or _49967_ (_18032_, _18030_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _49968_ (_18033_, _18032_, _17935_);
  and _49969_ (_18034_, _18033_, _18031_);
  and _49970_ (_18035_, _25777_, _23892_);
  or _49971_ (_18036_, _18035_, _18034_);
  and _49972_ (_10364_, _18036_, _22762_);
  and _49973_ (_18037_, _17263_, _23649_);
  and _49974_ (_18038_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  or _49975_ (_27194_, _18038_, _18037_);
  and _49976_ (_18039_, _17593_, _23898_);
  and _49977_ (_18040_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  or _49978_ (_10368_, _18040_, _18039_);
  and _49979_ (_18041_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and _49980_ (_18042_, _16311_, _23824_);
  or _49981_ (_10370_, _18042_, _18041_);
  and _49982_ (_18043_, _17447_, _23824_);
  and _49983_ (_18044_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or _49984_ (_10375_, _18044_, _18043_);
  and _49985_ (_18045_, _05119_, _24050_);
  and _49986_ (_18046_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  or _49987_ (_10377_, _18046_, _18045_);
  and _49988_ (_18047_, _17593_, _23649_);
  and _49989_ (_18048_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  or _49990_ (_10379_, _18048_, _18047_);
  and _49991_ (_18049_, _15856_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  or _49992_ (_18050_, _24315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _49993_ (_18051_, _18050_, _26118_);
  nor _49994_ (_18052_, _18051_, _26097_);
  nor _49995_ (_18053_, _18052_, _05168_);
  or _49996_ (_18054_, _18053_, _18049_);
  and _49997_ (_18055_, _18054_, _22762_);
  nor _49998_ (_18056_, _24299_, _24293_);
  and _49999_ (_10382_, _18056_, _18055_);
  or _50000_ (_18057_, _12675_, _23939_);
  and _50001_ (_18058_, _02079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _50002_ (_18059_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _50003_ (_18060_, _18059_, _18058_);
  or _50004_ (_18061_, _18060_, _02073_);
  and _50005_ (_18062_, _18061_, _22762_);
  and _50006_ (_10384_, _18062_, _18057_);
  and _50007_ (_18063_, _17593_, _24050_);
  and _50008_ (_18064_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  or _50009_ (_27297_, _18064_, _18063_);
  and _50010_ (_18065_, _16022_, _23824_);
  and _50011_ (_18066_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or _50012_ (_10390_, _18066_, _18065_);
  and _50013_ (_18067_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and _50014_ (_18068_, _16311_, _23898_);
  or _50015_ (_26976_, _18068_, _18067_);
  and _50016_ (_18069_, _17447_, _23747_);
  and _50017_ (_18070_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or _50018_ (_10395_, _18070_, _18069_);
  and _50019_ (_18071_, _06544_, _24050_);
  and _50020_ (_18072_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or _50021_ (_10397_, _18072_, _18071_);
  and _50022_ (_18073_, _16022_, _23778_);
  and _50023_ (_18074_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or _50024_ (_10399_, _18074_, _18073_);
  and _50025_ (_18075_, _17447_, _23946_);
  and _50026_ (_18076_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or _50027_ (_10401_, _18076_, _18075_);
  and _50028_ (_18077_, _17593_, _23707_);
  and _50029_ (_18078_, _17595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or _50030_ (_10403_, _18078_, _18077_);
  and _50031_ (_18079_, _16022_, _23946_);
  and _50032_ (_18080_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or _50033_ (_10406_, _18080_, _18079_);
  and _50034_ (_18081_, _24371_, _23946_);
  and _50035_ (_18082_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or _50036_ (_27198_, _18082_, _18081_);
  and _50037_ (_18083_, _17587_, _23778_);
  and _50038_ (_18084_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  or _50039_ (_27298_, _18084_, _18083_);
  and _50040_ (_18085_, _17447_, _24050_);
  and _50041_ (_18086_, _17449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or _50042_ (_10413_, _18086_, _18085_);
  and _50043_ (_18087_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and _50044_ (_18088_, _16311_, _23946_);
  or _50045_ (_26977_, _18088_, _18087_);
  and _50046_ (_18089_, _24371_, _23824_);
  and _50047_ (_18090_, _24373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or _50048_ (_10416_, _18090_, _18089_);
  nor _50049_ (_10431_, _05836_, rst);
  and _50050_ (_18091_, _17479_, _23778_);
  and _50051_ (_18092_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or _50052_ (_10436_, _18092_, _18091_);
  and _50053_ (_18093_, _25142_, _23747_);
  and _50054_ (_18094_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  or _50055_ (_10452_, _18094_, _18093_);
  and _50056_ (_18095_, _17587_, _23898_);
  and _50057_ (_18096_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  or _50058_ (_10454_, _18096_, _18095_);
  and _50059_ (_10471_, _05752_, _22762_);
  and _50060_ (_10500_, _05764_, _22762_);
  and _50061_ (_18097_, _17587_, _23824_);
  and _50062_ (_18098_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  or _50063_ (_10511_, _18098_, _18097_);
  and _50064_ (_10516_, _05820_, _22762_);
  and _50065_ (_18099_, _17479_, _23898_);
  and _50066_ (_18100_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or _50067_ (_27271_, _18100_, _18099_);
  and _50068_ (_10550_, _05808_, _22762_);
  and _50069_ (_18101_, _17479_, _23747_);
  and _50070_ (_18102_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or _50071_ (_10559_, _18102_, _18101_);
  and _50072_ (_18103_, _17587_, _23747_);
  and _50073_ (_18104_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  or _50074_ (_10569_, _18104_, _18103_);
  and _50075_ (_18105_, _04797_, _23707_);
  and _50076_ (_18106_, _04800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or _50077_ (_10574_, _18106_, _18105_);
  and _50078_ (_18107_, _16312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and _50079_ (_18108_, _16311_, _23649_);
  or _50080_ (_10599_, _18108_, _18107_);
  and _50081_ (_18109_, _17479_, _23649_);
  and _50082_ (_18110_, _17481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or _50083_ (_27272_, _18110_, _18109_);
  and _50084_ (_18111_, _15012_, _23747_);
  and _50085_ (_18112_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or _50086_ (_10606_, _18112_, _18111_);
  and _50087_ (_18113_, _06530_, _23778_);
  and _50088_ (_18114_, _06532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  or _50089_ (_10623_, _18114_, _18113_);
  and _50090_ (_18115_, _17587_, _23649_);
  and _50091_ (_18116_, _17589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  or _50092_ (_10625_, _18116_, _18115_);
  nor _50093_ (_10641_, _05791_, rst);
  and _50094_ (_18117_, _17221_, _23778_);
  and _50095_ (_18118_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or _50096_ (_10646_, _18118_, _18117_);
  and _50097_ (_18119_, _17439_, _23778_);
  and _50098_ (_18120_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or _50099_ (_27275_, _18120_, _18119_);
  and _50100_ (_18121_, _17229_, _23898_);
  and _50101_ (_18122_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or _50102_ (_10650_, _18122_, _18121_);
  and _50103_ (_10657_, _05778_, _22762_);
  and _50104_ (_18123_, _17581_, _23898_);
  and _50105_ (_18124_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or _50106_ (_10660_, _18124_, _18123_);
  and _50107_ (_18125_, _17581_, _23747_);
  and _50108_ (_18126_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or _50109_ (_10677_, _18126_, _18125_);
  and _50110_ (_18127_, _17439_, _23898_);
  and _50111_ (_18128_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or _50112_ (_10679_, _18128_, _18127_);
  and _50113_ (_18129_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  and _50114_ (_18130_, _16371_, _23649_);
  or _50115_ (_10701_, _18130_, _18129_);
  and _50116_ (_18131_, _17229_, _23649_);
  and _50117_ (_18132_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or _50118_ (_10706_, _18132_, _18131_);
  and _50119_ (_18133_, _17581_, _23946_);
  and _50120_ (_18134_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or _50121_ (_26916_, _18134_, _18133_);
  and _50122_ (_18135_, _12786_, _24050_);
  and _50123_ (_18136_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  or _50124_ (_10710_, _18136_, _18135_);
  and _50125_ (_18137_, _17388_, _23649_);
  and _50126_ (_18138_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or _50127_ (_27208_, _18138_, _18137_);
  and _50128_ (_18139_, _17439_, _23824_);
  and _50129_ (_18140_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or _50130_ (_27276_, _18140_, _18139_);
  and _50131_ (_18141_, _17388_, _23898_);
  and _50132_ (_18142_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or _50133_ (_10731_, _18142_, _18141_);
  and _50134_ (_18143_, _17439_, _23649_);
  and _50135_ (_18144_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or _50136_ (_10735_, _18144_, _18143_);
  and _50137_ (_18145_, _16022_, _23898_);
  and _50138_ (_18146_, _16024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or _50139_ (_10737_, _18146_, _18145_);
  and _50140_ (_18147_, _17581_, _24050_);
  and _50141_ (_18148_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or _50142_ (_10742_, _18148_, _18147_);
  and _50143_ (_18149_, _17388_, _23707_);
  and _50144_ (_18150_, _17390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or _50145_ (_10745_, _18150_, _18149_);
  and _50146_ (_18151_, _17229_, _23778_);
  and _50147_ (_18152_, _17231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or _50148_ (_10748_, _18152_, _18151_);
  and _50149_ (_18153_, _17439_, _23946_);
  and _50150_ (_18154_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or _50151_ (_10750_, _18154_, _18153_);
  and _50152_ (_18155_, _15850_, _23707_);
  and _50153_ (_18156_, _15852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  or _50154_ (_10755_, _18156_, _18155_);
  and _50155_ (_18157_, _17575_, _23778_);
  and _50156_ (_18158_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  or _50157_ (_26917_, _18158_, _18157_);
  and _50158_ (_18159_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  and _50159_ (_18160_, _16371_, _23946_);
  or _50160_ (_26974_, _18160_, _18159_);
  and _50161_ (_18161_, _02345_, _23747_);
  and _50162_ (_18162_, _02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or _50163_ (_10770_, _18162_, _18161_);
  and _50164_ (_18163_, _17575_, _23824_);
  and _50165_ (_18164_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  or _50166_ (_10775_, _18164_, _18163_);
  and _50167_ (_18165_, _08043_, _23946_);
  and _50168_ (_18166_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or _50169_ (_10780_, _18166_, _18165_);
  and _50170_ (_18167_, _23991_, _23076_);
  and _50171_ (_18168_, _18167_, _24050_);
  not _50172_ (_18169_, _18167_);
  and _50173_ (_18170_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  or _50174_ (_10784_, _18170_, _18168_);
  nor _50175_ (_18171_, _14782_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _50176_ (_18172_, _18171_, _26115_);
  and _50177_ (_18173_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _50178_ (_18174_, _18173_, _26118_);
  nor _50179_ (_18175_, _18174_, _18172_);
  nor _50180_ (_18176_, _18175_, _24299_);
  and _50181_ (_18177_, _24299_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _50182_ (_18178_, _18177_, _18176_);
  and _50183_ (_18179_, _18178_, _24294_);
  and _50184_ (_18180_, _24293_, _23642_);
  or _50185_ (_18181_, _18180_, _18179_);
  and _50186_ (_10788_, _18181_, _22762_);
  and _50187_ (_18182_, _17439_, _24050_);
  and _50188_ (_18183_, _17441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or _50189_ (_10791_, _18183_, _18182_);
  and _50190_ (_18184_, _08043_, _23824_);
  and _50191_ (_18185_, _08045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or _50192_ (_10797_, _18185_, _18184_);
  and _50193_ (_18186_, _18167_, _23707_);
  and _50194_ (_18187_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  or _50195_ (_10799_, _18187_, _18186_);
  and _50196_ (_18189_, _15012_, _23649_);
  and _50197_ (_18190_, _15014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or _50198_ (_27084_, _18190_, _18189_);
  and _50199_ (_18191_, _17575_, _23649_);
  and _50200_ (_18192_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  or _50201_ (_26919_, _18192_, _18191_);
  and _50202_ (_18193_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and _50203_ (_18194_, _16766_, _23946_);
  or _50204_ (_10806_, _18194_, _18193_);
  and _50205_ (_18195_, _12786_, _23946_);
  and _50206_ (_18196_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or _50207_ (_10810_, _18196_, _18195_);
  and _50208_ (_18197_, _23778_, _23077_);
  and _50209_ (_18198_, _23652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  or _50210_ (_10813_, _18198_, _18197_);
  and _50211_ (_18199_, _17575_, _23946_);
  and _50212_ (_18200_, _17577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  or _50213_ (_10826_, _18200_, _18199_);
  and _50214_ (_18201_, _17431_, _23778_);
  and _50215_ (_18202_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  or _50216_ (_10830_, _18202_, _18201_);
  and _50217_ (_18203_, _05410_, _23946_);
  and _50218_ (_18204_, _05412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  or _50219_ (_10832_, _18204_, _18203_);
  and _50220_ (_18205_, _17431_, _23824_);
  and _50221_ (_18206_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  or _50222_ (_10834_, _18206_, _18205_);
  and _50223_ (_18207_, _25733_, _23778_);
  and _50224_ (_18208_, _25735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or _50225_ (_10838_, _18208_, _18207_);
  and _50226_ (_18209_, _17569_, _23898_);
  and _50227_ (_18210_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  or _50228_ (_10844_, _18210_, _18209_);
  and _50229_ (_18211_, _02326_, _23824_);
  and _50230_ (_18212_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or _50231_ (_10856_, _18212_, _18211_);
  and _50232_ (_18213_, _17431_, _23747_);
  and _50233_ (_18214_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  or _50234_ (_10864_, _18214_, _18213_);
  and _50235_ (_18215_, _17569_, _23747_);
  and _50236_ (_18216_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  or _50237_ (_26920_, _18216_, _18215_);
  and _50238_ (_18217_, _24005_, _23076_);
  and _50239_ (_18218_, _18217_, _24050_);
  not _50240_ (_18219_, _18217_);
  and _50241_ (_18220_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or _50242_ (_27216_, _18220_, _18218_);
  and _50243_ (_18221_, _17431_, _23946_);
  and _50244_ (_18222_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  or _50245_ (_27277_, _18222_, _18221_);
  or _50246_ (_18223_, _24294_, _24043_);
  and _50247_ (_18224_, _26115_, _26098_);
  nand _50248_ (_18225_, _18224_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _50249_ (_18226_, _18225_, _24299_);
  and _50250_ (_18227_, _18226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand _50251_ (_18228_, _17665_, _26118_);
  or _50252_ (_18229_, _18225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _50253_ (_18230_, _18229_, _18228_);
  nor _50254_ (_18231_, _18230_, _24299_);
  or _50255_ (_18232_, _18231_, _24293_);
  or _50256_ (_18233_, _18232_, _18227_);
  and _50257_ (_18234_, _18233_, _22762_);
  and _50258_ (_10873_, _18234_, _18223_);
  and _50259_ (_18235_, _17431_, _23707_);
  and _50260_ (_18236_, _17433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  or _50261_ (_10876_, _18236_, _18235_);
  and _50262_ (_18237_, _17569_, _23649_);
  and _50263_ (_18238_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  or _50264_ (_10880_, _18238_, _18237_);
  and _50265_ (_18239_, _17569_, _23707_);
  and _50266_ (_18240_, _17571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  or _50267_ (_10886_, _18240_, _18239_);
  and _50268_ (_18241_, _24050_, _23755_);
  and _50269_ (_18242_, _23780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  or _50270_ (_10888_, _18242_, _18241_);
  and _50271_ (_18243_, _17416_, _23898_);
  and _50272_ (_18244_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  or _50273_ (_10892_, _18244_, _18243_);
  and _50274_ (_18245_, _17207_, _23898_);
  and _50275_ (_18246_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or _50276_ (_10895_, _18246_, _18245_);
  and _50277_ (_18247_, _18167_, _23946_);
  and _50278_ (_18248_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  or _50279_ (_10897_, _18248_, _18247_);
  and _50280_ (_18249_, _16767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and _50281_ (_18250_, _16766_, _23707_);
  or _50282_ (_10902_, _18250_, _18249_);
  and _50283_ (_18251_, _17551_, _23778_);
  and _50284_ (_18252_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or _50285_ (_26922_, _18252_, _18251_);
  and _50286_ (_18253_, _17416_, _23824_);
  and _50287_ (_18254_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  or _50288_ (_10915_, _18254_, _18253_);
  and _50289_ (_18255_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  and _50290_ (_18256_, _16758_, _23778_);
  or _50291_ (_26952_, _18256_, _18255_);
  and _50292_ (_18257_, _17207_, _23778_);
  and _50293_ (_18258_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or _50294_ (_10920_, _18258_, _18257_);
  and _50295_ (_18259_, _17551_, _23824_);
  and _50296_ (_18260_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or _50297_ (_10928_, _18260_, _18259_);
  and _50298_ (_18261_, _15004_, _23946_);
  and _50299_ (_18262_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or _50300_ (_10930_, _18262_, _18261_);
  and _50301_ (_18263_, _17207_, _23707_);
  and _50302_ (_18264_, _17209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or _50303_ (_10938_, _18264_, _18263_);
  and _50304_ (_18265_, _25260_, _24654_);
  nand _50305_ (_18266_, _18265_, _23594_);
  or _50306_ (_18267_, _18265_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _50307_ (_18268_, _18267_, _24645_);
  and _50308_ (_18269_, _18268_, _18266_);
  nand _50309_ (_18270_, _25266_, _23702_);
  or _50310_ (_18271_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _50311_ (_18272_, _18271_, _24069_);
  and _50312_ (_18273_, _18272_, _18270_);
  and _50313_ (_18274_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _50314_ (_18275_, _18274_, rst);
  or _50315_ (_18276_, _18275_, _18273_);
  or _50316_ (_10940_, _18276_, _18269_);
  and _50317_ (_18277_, _17416_, _23649_);
  and _50318_ (_18278_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  or _50319_ (_10945_, _18278_, _18277_);
  and _50320_ (_18279_, _12786_, _23649_);
  and _50321_ (_18280_, _12788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  or _50322_ (_10947_, _18280_, _18279_);
  and _50323_ (_18281_, _06544_, _23824_);
  and _50324_ (_18282_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or _50325_ (_10952_, _18282_, _18281_);
  and _50326_ (_18283_, _17416_, _24050_);
  and _50327_ (_18284_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  or _50328_ (_10955_, _18284_, _18283_);
  and _50329_ (_18285_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  and _50330_ (_18286_, _16758_, _23824_);
  or _50331_ (_10958_, _18286_, _18285_);
  and _50332_ (_18287_, _17551_, _23747_);
  and _50333_ (_18288_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or _50334_ (_10960_, _18288_, _18287_);
  and _50335_ (_18289_, _15004_, _23649_);
  and _50336_ (_18290_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or _50337_ (_27083_, _18290_, _18289_);
  and _50338_ (_18291_, _07536_, _23649_);
  and _50339_ (_18292_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  or _50340_ (_10966_, _18292_, _18291_);
  and _50341_ (_18293_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  and _50342_ (_18294_, _16758_, _23649_);
  or _50343_ (_10968_, _18294_, _18293_);
  and _50344_ (_18295_, _17410_, _23898_);
  and _50345_ (_18296_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or _50346_ (_10973_, _18296_, _18295_);
  and _50347_ (_18297_, _15004_, _23747_);
  and _50348_ (_18298_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or _50349_ (_10975_, _18298_, _18297_);
  and _50350_ (_18299_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  and _50351_ (_18300_, _12829_, _23747_);
  or _50352_ (_10980_, _18300_, _18299_);
  and _50353_ (_18301_, _06544_, _23898_);
  and _50354_ (_18302_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or _50355_ (_10982_, _18302_, _18301_);
  and _50356_ (_18304_, _17551_, _24050_);
  and _50357_ (_18305_, _17553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or _50358_ (_26923_, _18305_, _18304_);
  and _50359_ (_18306_, _12830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  and _50360_ (_18307_, _12829_, _23778_);
  or _50361_ (_27223_, _18307_, _18306_);
  and _50362_ (_18308_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  and _50363_ (_18309_, _16758_, _24050_);
  or _50364_ (_26953_, _18309_, _18308_);
  and _50365_ (_18310_, _17410_, _23824_);
  and _50366_ (_18311_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or _50367_ (_27279_, _18311_, _18310_);
  and _50368_ (_18312_, _17719_, _23898_);
  and _50369_ (_18313_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  or _50370_ (_26924_, _18313_, _18312_);
  and _50371_ (_18314_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and _50372_ (_18315_, _08351_, _23707_);
  or _50373_ (_27226_, _18315_, _18314_);
  and _50374_ (_18316_, _16759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  and _50375_ (_18317_, _16758_, _23707_);
  or _50376_ (_26954_, _18317_, _18316_);
  and _50377_ (_18318_, _17410_, _23649_);
  and _50378_ (_18319_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or _50379_ (_27280_, _18319_, _18318_);
  and _50380_ (_18320_, _08352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and _50381_ (_18321_, _08351_, _23649_);
  or _50382_ (_27225_, _18321_, _18320_);
  and _50383_ (_18322_, _17410_, _24050_);
  and _50384_ (_18323_, _17412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or _50385_ (_27281_, _18323_, _18322_);
  and _50386_ (_18324_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  and _50387_ (_18325_, _05193_, _23946_);
  or _50388_ (_27229_, _18325_, _18324_);
  and _50389_ (_18326_, _17719_, _23824_);
  and _50390_ (_18327_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  or _50391_ (_26925_, _18327_, _18326_);
  and _50392_ (_18328_, _17215_, _23707_);
  and _50393_ (_18329_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  or _50394_ (_27218_, _18329_, _18328_);
  and _50395_ (_18330_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  and _50396_ (_18331_, _05193_, _23824_);
  or _50397_ (_27227_, _18331_, _18330_);
  and _50398_ (_18332_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  and _50399_ (_18333_, _16371_, _23707_);
  or _50400_ (_26975_, _18333_, _18332_);
  and _50401_ (_18334_, _17719_, _23649_);
  and _50402_ (_18335_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  or _50403_ (_26926_, _18335_, _18334_);
  and _50404_ (_18336_, _17404_, _23778_);
  and _50405_ (_18337_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or _50406_ (_27282_, _18337_, _18336_);
  and _50407_ (_18338_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  and _50408_ (_18339_, _05199_, _23946_);
  or _50409_ (_27231_, _18339_, _18338_);
  and _50410_ (_18340_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  and _50411_ (_18341_, _16752_, _23824_);
  or _50412_ (_26955_, _18341_, _18340_);
  and _50413_ (_18342_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  and _50414_ (_18343_, _16752_, _23649_);
  or _50415_ (_26956_, _18343_, _18342_);
  and _50416_ (_18344_, _18167_, _23898_);
  and _50417_ (_18345_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  or _50418_ (_27220_, _18345_, _18344_);
  and _50419_ (_18346_, _17719_, _23946_);
  and _50420_ (_18347_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  or _50421_ (_26927_, _18347_, _18346_);
  and _50422_ (_18348_, _17404_, _23898_);
  and _50423_ (_18349_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or _50424_ (_27283_, _18349_, _18348_);
  and _50425_ (_18350_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  and _50426_ (_18351_, _16752_, _24050_);
  or _50427_ (_26957_, _18351_, _18350_);
  and _50428_ (_18352_, _17719_, _24050_);
  and _50429_ (_18353_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  or _50430_ (_26928_, _18353_, _18352_);
  and _50431_ (_18354_, _17404_, _23747_);
  and _50432_ (_18355_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or _50433_ (_27284_, _18355_, _18354_);
  and _50434_ (_18356_, _17404_, _23946_);
  and _50435_ (_18357_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or _50436_ (_27285_, _18357_, _18356_);
  and _50437_ (_18358_, _17719_, _23707_);
  and _50438_ (_18359_, _17721_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or _50439_ (_26929_, _18359_, _18358_);
  and _50440_ (_18360_, _16753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  and _50441_ (_18361_, _16752_, _23707_);
  or _50442_ (_26958_, _18361_, _18360_);
  and _50443_ (_18362_, _18167_, _23778_);
  and _50444_ (_18363_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  or _50445_ (_27219_, _18363_, _18362_);
  and _50446_ (_18364_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  and _50447_ (_18365_, _07492_, _23778_);
  or _50448_ (_27239_, _18365_, _18364_);
  and _50449_ (_18366_, _06544_, _23649_);
  and _50450_ (_18367_, _06547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or _50451_ (_27145_, _18367_, _18366_);
  and _50452_ (_18368_, _17539_, _23898_);
  and _50453_ (_18369_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or _50454_ (_26930_, _18369_, _18368_);
  and _50455_ (_18370_, _17404_, _23707_);
  and _50456_ (_18371_, _17406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or _50457_ (_27286_, _18371_, _18370_);
  and _50458_ (_18372_, _25164_, _24654_);
  nand _50459_ (_18373_, _18372_, _23594_);
  or _50460_ (_18374_, _18372_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _50461_ (_18375_, _18374_, _24645_);
  and _50462_ (_18376_, _18375_, _18373_);
  nand _50463_ (_18377_, _25173_, _23702_);
  or _50464_ (_18378_, _25173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _50465_ (_18379_, _18378_, _24069_);
  and _50466_ (_18380_, _18379_, _18377_);
  and _50467_ (_18381_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _50468_ (_18382_, _18381_, rst);
  or _50469_ (_18383_, _18382_, _18380_);
  or _50470_ (_11053_, _18383_, _18376_);
  and _50471_ (_18384_, _17539_, _23747_);
  and _50472_ (_18385_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or _50473_ (_11057_, _18385_, _18384_);
  and _50474_ (_18386_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and _50475_ (_18387_, _16748_, _23898_);
  or _50476_ (_11062_, _18387_, _18386_);
  and _50477_ (_18388_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and _50478_ (_18389_, _16748_, _23824_);
  or _50479_ (_26959_, _18389_, _18388_);
  and _50480_ (_18390_, _17396_, _23778_);
  and _50481_ (_18391_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  or _50482_ (_11071_, _18391_, _18390_);
  and _50483_ (_18392_, _07493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  and _50484_ (_18393_, _07492_, _23649_);
  or _50485_ (_11074_, _18393_, _18392_);
  and _50486_ (_18394_, _17539_, _23946_);
  and _50487_ (_18395_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or _50488_ (_26931_, _18395_, _18394_);
  and _50489_ (_18396_, _17396_, _23824_);
  and _50490_ (_18397_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  or _50491_ (_11077_, _18397_, _18396_);
  and _50492_ (_18398_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  and _50493_ (_18399_, _17775_, _23649_);
  or _50494_ (_11080_, _18399_, _18398_);
  and _50495_ (_18400_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and _50496_ (_18401_, _16748_, _23747_);
  or _50497_ (_11083_, _18401_, _18400_);
  or _50498_ (_18402_, _24294_, _23939_);
  and _50499_ (_18403_, _26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _50500_ (_18404_, _18403_, _26118_);
  nand _50501_ (_18405_, _18225_, _18224_);
  and _50502_ (_18406_, _18405_, _18404_);
  nor _50503_ (_18407_, _18406_, _24299_);
  and _50504_ (_18408_, _18226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _50505_ (_18409_, _18408_, _18407_);
  or _50506_ (_18410_, _18409_, _24293_);
  and _50507_ (_18411_, _18410_, _22762_);
  and _50508_ (_11085_, _18411_, _18402_);
  and _50509_ (_18412_, _25350_, _24654_);
  nand _50510_ (_18413_, _18412_, _23594_);
  or _50511_ (_18414_, _18412_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _50512_ (_18415_, _18414_, _24645_);
  and _50513_ (_18416_, _18415_, _18413_);
  nand _50514_ (_18417_, _25358_, _23702_);
  or _50515_ (_18418_, _25358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _50516_ (_18419_, _18418_, _24069_);
  and _50517_ (_18420_, _18419_, _18417_);
  and _50518_ (_18421_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _50519_ (_18422_, _18421_, rst);
  or _50520_ (_18423_, _18422_, _18420_);
  or _50521_ (_11086_, _18423_, _18416_);
  and _50522_ (_18424_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  and _50523_ (_18425_, _17775_, _23898_);
  or _50524_ (_11092_, _18425_, _18424_);
  and _50525_ (_18426_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and _50526_ (_18427_, _16748_, _23946_);
  or _50527_ (_11094_, _18427_, _18426_);
  and _50528_ (_18428_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  and _50529_ (_18429_, _16319_, _23707_);
  or _50530_ (_26971_, _18429_, _18428_);
  and _50531_ (_18430_, _17539_, _24050_);
  and _50532_ (_18431_, _17541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or _50533_ (_26932_, _18431_, _18430_);
  and _50534_ (_18432_, _17396_, _23747_);
  and _50535_ (_18433_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  or _50536_ (_27287_, _18433_, _18432_);
  and _50537_ (_18434_, _15004_, _23707_);
  and _50538_ (_18435_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or _50539_ (_11100_, _18435_, _18434_);
  and _50540_ (_18436_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  and _50541_ (_18437_, _02306_, _23778_);
  or _50542_ (_11102_, _18437_, _18436_);
  and _50543_ (_18438_, _17535_, _23778_);
  and _50544_ (_18439_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or _50545_ (_11104_, _18439_, _18438_);
  and _50546_ (_18440_, _17396_, _24050_);
  and _50547_ (_18441_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  or _50548_ (_11106_, _18441_, _18440_);
  and _50549_ (_18442_, _16749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and _50550_ (_18443_, _16748_, _23707_);
  or _50551_ (_11109_, _18443_, _18442_);
  and _50552_ (_18444_, _25439_, _24654_);
  nand _50553_ (_18445_, _18444_, _23594_);
  or _50554_ (_18446_, _18444_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _50555_ (_18447_, _18446_, _24645_);
  and _50556_ (_18448_, _18447_, _18445_);
  nand _50557_ (_18449_, _25446_, _23702_);
  or _50558_ (_18450_, _25446_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _50559_ (_18451_, _18450_, _24069_);
  and _50560_ (_18452_, _18451_, _18449_);
  and _50561_ (_18453_, _25181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _50562_ (_18454_, _18453_, rst);
  or _50563_ (_18455_, _18454_, _18452_);
  or _50564_ (_11111_, _18455_, _18448_);
  and _50565_ (_18456_, _06602_, _23946_);
  and _50566_ (_18457_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  or _50567_ (_11117_, _18457_, _18456_);
  and _50568_ (_18458_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  and _50569_ (_18459_, _16742_, _23778_);
  or _50570_ (_11119_, _18459_, _18458_);
  and _50571_ (_18460_, _17396_, _23707_);
  and _50572_ (_18461_, _17398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  or _50573_ (_27288_, _18461_, _18460_);
  and _50574_ (_18462_, _17535_, _23898_);
  and _50575_ (_18463_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or _50576_ (_11124_, _18463_, _18462_);
  and _50577_ (_18464_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  and _50578_ (_18465_, _16742_, _23898_);
  or _50579_ (_26961_, _18465_, _18464_);
  and _50580_ (_18466_, _17535_, _23747_);
  and _50581_ (_18467_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or _50582_ (_11127_, _18467_, _18466_);
  and _50583_ (_18468_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and _50584_ (_18469_, _13763_, _23824_);
  or _50585_ (_11132_, _18469_, _18468_);
  and _50586_ (_18470_, _17378_, _23898_);
  and _50587_ (_18471_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  or _50588_ (_11134_, _18471_, _18470_);
  and _50589_ (_18472_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  and _50590_ (_18473_, _24222_, _23824_);
  or _50591_ (_11136_, _18473_, _18472_);
  and _50592_ (_18474_, _17535_, _23649_);
  and _50593_ (_18475_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or _50594_ (_11139_, _18475_, _18474_);
  and _50595_ (_18476_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  and _50596_ (_18477_, _16742_, _23824_);
  or _50597_ (_11141_, _18477_, _18476_);
  and _50598_ (_18478_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  and _50599_ (_18479_, _16742_, _23649_);
  or _50600_ (_11147_, _18479_, _18478_);
  and _50601_ (_18480_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  and _50602_ (_18481_, _16742_, _24050_);
  or _50603_ (_11149_, _18481_, _18480_);
  and _50604_ (_18482_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and _50605_ (_18483_, _17255_, _23707_);
  or _50606_ (_11153_, _18483_, _18482_);
  and _50607_ (_18484_, _08198_, _23707_);
  and _50608_ (_18485_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or _50609_ (_11156_, _18485_, _18484_);
  and _50610_ (_18486_, _16743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  and _50611_ (_18487_, _16742_, _23707_);
  or _50612_ (_11159_, _18487_, _18486_);
  and _50613_ (_18488_, _04762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and _50614_ (_18489_, _04761_, _23778_);
  or _50615_ (_11161_, _18489_, _18488_);
  and _50616_ (_18490_, _08478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  and _50617_ (_18491_, _08477_, _23778_);
  or _50618_ (_11164_, _18491_, _18490_);
  and _50619_ (_18492_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and _50620_ (_18493_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or _50621_ (_18494_, _18493_, _18492_);
  and _50622_ (_18495_, _18494_, _02393_);
  and _50623_ (_18496_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and _50624_ (_18497_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or _50625_ (_18498_, _18497_, _18496_);
  and _50626_ (_18499_, _18498_, _02445_);
  or _50627_ (_18500_, _18499_, _18495_);
  and _50628_ (_18501_, _18500_, _02421_);
  and _50629_ (_18502_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and _50630_ (_18503_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or _50631_ (_18504_, _18503_, _18502_);
  and _50632_ (_18505_, _18504_, _02393_);
  and _50633_ (_18506_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and _50634_ (_18507_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or _50635_ (_18508_, _18507_, _18506_);
  and _50636_ (_18509_, _18508_, _02445_);
  or _50637_ (_18510_, _18509_, _18505_);
  and _50638_ (_18511_, _18510_, _02459_);
  or _50639_ (_18512_, _18511_, _18501_);
  and _50640_ (_18513_, _18512_, _02458_);
  or _50641_ (_18514_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or _50642_ (_18515_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and _50643_ (_18516_, _18515_, _18514_);
  and _50644_ (_18517_, _18516_, _02393_);
  or _50645_ (_18518_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or _50646_ (_18520_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and _50647_ (_18521_, _18520_, _18518_);
  and _50648_ (_18522_, _18521_, _02445_);
  or _50649_ (_18523_, _18522_, _18517_);
  and _50650_ (_18524_, _18523_, _02421_);
  or _50651_ (_18525_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or _50652_ (_18526_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and _50653_ (_18527_, _18526_, _18525_);
  and _50654_ (_18528_, _18527_, _02393_);
  or _50655_ (_18529_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or _50656_ (_18530_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and _50657_ (_18531_, _18530_, _18529_);
  and _50658_ (_18532_, _18531_, _02445_);
  or _50659_ (_18533_, _18532_, _18528_);
  and _50660_ (_18534_, _18533_, _02459_);
  or _50661_ (_18535_, _18534_, _18524_);
  and _50662_ (_18536_, _18535_, _02414_);
  or _50663_ (_18537_, _18536_, _18513_);
  and _50664_ (_18538_, _18537_, _02398_);
  and _50665_ (_18539_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and _50666_ (_18540_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or _50667_ (_18541_, _18540_, _18539_);
  and _50668_ (_18542_, _18541_, _02393_);
  and _50669_ (_18543_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and _50670_ (_18544_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or _50671_ (_18545_, _18544_, _18543_);
  and _50672_ (_18546_, _18545_, _02445_);
  or _50673_ (_18547_, _18546_, _18542_);
  and _50674_ (_18548_, _18547_, _02421_);
  and _50675_ (_18549_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and _50676_ (_18550_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or _50677_ (_18551_, _18550_, _18549_);
  and _50678_ (_18552_, _18551_, _02393_);
  and _50679_ (_18553_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and _50680_ (_18554_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or _50681_ (_18555_, _18554_, _18553_);
  and _50682_ (_18556_, _18555_, _02445_);
  or _50683_ (_18557_, _18556_, _18552_);
  and _50684_ (_18558_, _18557_, _02459_);
  or _50685_ (_18559_, _18558_, _18548_);
  and _50686_ (_18560_, _18559_, _02458_);
  or _50687_ (_18561_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or _50688_ (_18562_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and _50689_ (_18563_, _18562_, _02445_);
  and _50690_ (_18564_, _18563_, _18561_);
  or _50691_ (_18565_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or _50692_ (_18566_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and _50693_ (_18567_, _18566_, _02393_);
  and _50694_ (_18568_, _18567_, _18565_);
  or _50695_ (_18569_, _18568_, _18564_);
  and _50696_ (_18570_, _18569_, _02421_);
  or _50697_ (_18571_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or _50698_ (_18572_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and _50699_ (_18573_, _18572_, _02445_);
  and _50700_ (_18574_, _18573_, _18571_);
  or _50701_ (_18575_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or _50702_ (_18576_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  and _50703_ (_18577_, _18576_, _02393_);
  and _50704_ (_18578_, _18577_, _18575_);
  or _50705_ (_18579_, _18578_, _18574_);
  and _50706_ (_18580_, _18579_, _02459_);
  or _50707_ (_18581_, _18580_, _18570_);
  and _50708_ (_18582_, _18581_, _02414_);
  or _50709_ (_18583_, _18582_, _18560_);
  and _50710_ (_18584_, _18583_, _02496_);
  or _50711_ (_18585_, _18584_, _18538_);
  and _50712_ (_18586_, _18585_, _02400_);
  and _50713_ (_18587_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and _50714_ (_18588_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or _50715_ (_18589_, _18588_, _18587_);
  and _50716_ (_18590_, _18589_, _02393_);
  and _50717_ (_18591_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and _50718_ (_18592_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or _50719_ (_18593_, _18592_, _18591_);
  and _50720_ (_18594_, _18593_, _02445_);
  or _50721_ (_18595_, _18594_, _18590_);
  or _50722_ (_18596_, _18595_, _02459_);
  and _50723_ (_18597_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and _50724_ (_18598_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or _50725_ (_18599_, _18598_, _18597_);
  and _50726_ (_18601_, _18599_, _02393_);
  and _50727_ (_18602_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and _50728_ (_18603_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or _50729_ (_18604_, _18603_, _18602_);
  and _50730_ (_18605_, _18604_, _02445_);
  or _50731_ (_18606_, _18605_, _18601_);
  or _50732_ (_18607_, _18606_, _02421_);
  and _50733_ (_18608_, _18607_, _02458_);
  and _50734_ (_18609_, _18608_, _18596_);
  or _50735_ (_18610_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or _50736_ (_18611_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and _50737_ (_18612_, _18611_, _02445_);
  and _50738_ (_18613_, _18612_, _18610_);
  or _50739_ (_18614_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or _50740_ (_18615_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and _50741_ (_18616_, _18615_, _02393_);
  and _50742_ (_18617_, _18616_, _18614_);
  or _50743_ (_18618_, _18617_, _18613_);
  or _50744_ (_18619_, _18618_, _02459_);
  or _50745_ (_18620_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or _50746_ (_18621_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and _50747_ (_18622_, _18621_, _02445_);
  and _50748_ (_18623_, _18622_, _18620_);
  or _50749_ (_18624_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or _50750_ (_18625_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and _50751_ (_18626_, _18625_, _02393_);
  and _50752_ (_18627_, _18626_, _18624_);
  or _50753_ (_18628_, _18627_, _18623_);
  or _50754_ (_18629_, _18628_, _02421_);
  and _50755_ (_18630_, _18629_, _02414_);
  and _50756_ (_18631_, _18630_, _18619_);
  or _50757_ (_18632_, _18631_, _18609_);
  and _50758_ (_18633_, _18632_, _02496_);
  and _50759_ (_18634_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and _50760_ (_18635_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or _50761_ (_18636_, _18635_, _18634_);
  and _50762_ (_18637_, _18636_, _02393_);
  and _50763_ (_18638_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and _50764_ (_18639_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or _50765_ (_18640_, _18639_, _18638_);
  and _50766_ (_18641_, _18640_, _02445_);
  or _50767_ (_18642_, _18641_, _18637_);
  or _50768_ (_18643_, _18642_, _02459_);
  and _50769_ (_18644_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and _50770_ (_18645_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or _50771_ (_18646_, _18645_, _18644_);
  and _50772_ (_18647_, _18646_, _02393_);
  and _50773_ (_18648_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and _50774_ (_18649_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or _50775_ (_18650_, _18649_, _18648_);
  and _50776_ (_18651_, _18650_, _02445_);
  or _50777_ (_18652_, _18651_, _18647_);
  or _50778_ (_18653_, _18652_, _02421_);
  and _50779_ (_18654_, _18653_, _02458_);
  and _50780_ (_18655_, _18654_, _18643_);
  or _50781_ (_18656_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or _50782_ (_18657_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and _50783_ (_18658_, _18657_, _18656_);
  and _50784_ (_18659_, _18658_, _02393_);
  or _50785_ (_18660_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or _50786_ (_18661_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and _50787_ (_18662_, _18661_, _18660_);
  and _50788_ (_18663_, _18662_, _02445_);
  or _50789_ (_18664_, _18663_, _18659_);
  or _50790_ (_18665_, _18664_, _02459_);
  or _50791_ (_18666_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or _50792_ (_18667_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and _50793_ (_18668_, _18667_, _18666_);
  and _50794_ (_18669_, _18668_, _02393_);
  or _50795_ (_18670_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or _50796_ (_18671_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and _50797_ (_18672_, _18671_, _18670_);
  and _50798_ (_18673_, _18672_, _02445_);
  or _50799_ (_18674_, _18673_, _18669_);
  or _50800_ (_18675_, _18674_, _02421_);
  and _50801_ (_18676_, _18675_, _02414_);
  and _50802_ (_18677_, _18676_, _18665_);
  or _50803_ (_18678_, _18677_, _18655_);
  and _50804_ (_18679_, _18678_, _02398_);
  or _50805_ (_18680_, _18679_, _18633_);
  and _50806_ (_18681_, _18680_, _02546_);
  or _50807_ (_18682_, _18681_, _18586_);
  and _50808_ (_18683_, _18682_, _02646_);
  or _50809_ (_18684_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or _50810_ (_18685_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  and _50811_ (_18686_, _18685_, _02445_);
  and _50812_ (_18687_, _18686_, _18684_);
  or _50813_ (_18688_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or _50814_ (_18689_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and _50815_ (_18690_, _18689_, _02393_);
  and _50816_ (_18691_, _18690_, _18688_);
  or _50817_ (_18692_, _18691_, _18687_);
  and _50818_ (_18693_, _18692_, _02459_);
  or _50819_ (_18694_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or _50820_ (_18695_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and _50821_ (_18696_, _18695_, _02445_);
  and _50822_ (_18697_, _18696_, _18694_);
  or _50823_ (_18698_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or _50824_ (_18699_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  and _50825_ (_18700_, _18699_, _02393_);
  and _50826_ (_18701_, _18700_, _18698_);
  or _50827_ (_18702_, _18701_, _18697_);
  and _50828_ (_18703_, _18702_, _02421_);
  or _50829_ (_18704_, _18703_, _18693_);
  and _50830_ (_18705_, _18704_, _02414_);
  and _50831_ (_18706_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and _50832_ (_18707_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or _50833_ (_18708_, _18707_, _18706_);
  and _50834_ (_18709_, _18708_, _02393_);
  and _50835_ (_18710_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and _50836_ (_18711_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or _50837_ (_18712_, _18711_, _18710_);
  and _50838_ (_18713_, _18712_, _02445_);
  or _50839_ (_18714_, _18713_, _18709_);
  and _50840_ (_18715_, _18714_, _02459_);
  and _50841_ (_18716_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and _50842_ (_18717_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or _50843_ (_18718_, _18717_, _18716_);
  and _50844_ (_18719_, _18718_, _02393_);
  and _50845_ (_18720_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and _50846_ (_18721_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or _50847_ (_18722_, _18721_, _18720_);
  and _50848_ (_18723_, _18722_, _02445_);
  or _50849_ (_18724_, _18723_, _18719_);
  and _50850_ (_18725_, _18724_, _02421_);
  or _50851_ (_18726_, _18725_, _18715_);
  and _50852_ (_18727_, _18726_, _02458_);
  or _50853_ (_18728_, _18727_, _18705_);
  and _50854_ (_18729_, _18728_, _02496_);
  or _50855_ (_18730_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or _50856_ (_18731_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and _50857_ (_18732_, _18731_, _18730_);
  and _50858_ (_18733_, _18732_, _02393_);
  or _50859_ (_18734_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or _50860_ (_18735_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and _50861_ (_18736_, _18735_, _18734_);
  and _50862_ (_18737_, _18736_, _02445_);
  or _50863_ (_18738_, _18737_, _18733_);
  and _50864_ (_18739_, _18738_, _02459_);
  or _50865_ (_18740_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or _50866_ (_18741_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and _50867_ (_18742_, _18741_, _18740_);
  and _50868_ (_18743_, _18742_, _02393_);
  or _50869_ (_18744_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or _50870_ (_18745_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and _50871_ (_18746_, _18745_, _18744_);
  and _50872_ (_18747_, _18746_, _02445_);
  or _50873_ (_18748_, _18747_, _18743_);
  and _50874_ (_18749_, _18748_, _02421_);
  or _50875_ (_18750_, _18749_, _18739_);
  and _50876_ (_18751_, _18750_, _02414_);
  and _50877_ (_18752_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and _50878_ (_18753_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or _50879_ (_18754_, _18753_, _18752_);
  and _50880_ (_18755_, _18754_, _02393_);
  and _50881_ (_18756_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and _50882_ (_18757_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or _50883_ (_18758_, _18757_, _18756_);
  and _50884_ (_18759_, _18758_, _02445_);
  or _50885_ (_18760_, _18759_, _18755_);
  and _50886_ (_18761_, _18760_, _02459_);
  and _50887_ (_18762_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and _50888_ (_18763_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or _50889_ (_18764_, _18763_, _18762_);
  and _50890_ (_18765_, _18764_, _02393_);
  and _50891_ (_18766_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and _50892_ (_18767_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or _50893_ (_18768_, _18767_, _18766_);
  and _50894_ (_18769_, _18768_, _02445_);
  or _50895_ (_18770_, _18769_, _18765_);
  and _50896_ (_18771_, _18770_, _02421_);
  or _50897_ (_18772_, _18771_, _18761_);
  and _50898_ (_18773_, _18772_, _02458_);
  or _50899_ (_18774_, _18773_, _18751_);
  and _50900_ (_18775_, _18774_, _02398_);
  or _50901_ (_18776_, _18775_, _18729_);
  and _50902_ (_18777_, _18776_, _02400_);
  and _50903_ (_18778_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and _50904_ (_18779_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or _50905_ (_18780_, _18779_, _18778_);
  and _50906_ (_18781_, _18780_, _02393_);
  and _50907_ (_18782_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and _50908_ (_18783_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or _50909_ (_18784_, _18783_, _18782_);
  and _50910_ (_18785_, _18784_, _02445_);
  or _50911_ (_18786_, _18785_, _18781_);
  or _50912_ (_18787_, _18786_, _02459_);
  and _50913_ (_18788_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and _50914_ (_18789_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or _50915_ (_18790_, _18789_, _18788_);
  and _50916_ (_18791_, _18790_, _02393_);
  and _50917_ (_18792_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and _50918_ (_18793_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or _50919_ (_18794_, _18793_, _18792_);
  and _50920_ (_18795_, _18794_, _02445_);
  or _50921_ (_18796_, _18795_, _18791_);
  or _50922_ (_18797_, _18796_, _02421_);
  and _50923_ (_18798_, _18797_, _02458_);
  and _50924_ (_18799_, _18798_, _18787_);
  or _50925_ (_18800_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or _50926_ (_18801_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and _50927_ (_18802_, _18801_, _18800_);
  and _50928_ (_18803_, _18802_, _02393_);
  or _50929_ (_18804_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or _50930_ (_18805_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and _50931_ (_18806_, _18805_, _18804_);
  and _50932_ (_18807_, _18806_, _02445_);
  or _50933_ (_18808_, _18807_, _18803_);
  or _50934_ (_18809_, _18808_, _02459_);
  or _50935_ (_18810_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or _50936_ (_18811_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and _50937_ (_18812_, _18811_, _18810_);
  and _50938_ (_18813_, _18812_, _02393_);
  or _50939_ (_18814_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or _50940_ (_18815_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and _50941_ (_18816_, _18815_, _18814_);
  and _50942_ (_18817_, _18816_, _02445_);
  or _50943_ (_18818_, _18817_, _18813_);
  or _50944_ (_18819_, _18818_, _02421_);
  and _50945_ (_18820_, _18819_, _02414_);
  and _50946_ (_18821_, _18820_, _18809_);
  or _50947_ (_18822_, _18821_, _18799_);
  and _50948_ (_18823_, _18822_, _02398_);
  and _50949_ (_18824_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and _50950_ (_18825_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or _50951_ (_18826_, _18825_, _18824_);
  and _50952_ (_18827_, _18826_, _02393_);
  and _50953_ (_18828_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and _50954_ (_18829_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or _50955_ (_18830_, _18829_, _18828_);
  and _50956_ (_18831_, _18830_, _02445_);
  or _50957_ (_18832_, _18831_, _18827_);
  or _50958_ (_18833_, _18832_, _02459_);
  and _50959_ (_18834_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and _50960_ (_18835_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or _50961_ (_18836_, _18835_, _18834_);
  and _50962_ (_18837_, _18836_, _02393_);
  and _50963_ (_18838_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and _50964_ (_18839_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or _50965_ (_18840_, _18839_, _18838_);
  and _50966_ (_18841_, _18840_, _02445_);
  or _50967_ (_18842_, _18841_, _18837_);
  or _50968_ (_18843_, _18842_, _02421_);
  and _50969_ (_18844_, _18843_, _02458_);
  and _50970_ (_18845_, _18844_, _18833_);
  or _50971_ (_18846_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or _50972_ (_18847_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and _50973_ (_18848_, _18847_, _02445_);
  and _50974_ (_18849_, _18848_, _18846_);
  or _50975_ (_18850_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or _50976_ (_18851_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and _50977_ (_18852_, _18851_, _02393_);
  and _50978_ (_18853_, _18852_, _18850_);
  or _50979_ (_18854_, _18853_, _18849_);
  or _50980_ (_18855_, _18854_, _02459_);
  or _50981_ (_18856_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or _50982_ (_18857_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and _50983_ (_18858_, _18857_, _02445_);
  and _50984_ (_18859_, _18858_, _18856_);
  or _50985_ (_18860_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or _50986_ (_18861_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and _50987_ (_18862_, _18861_, _02393_);
  and _50988_ (_18863_, _18862_, _18860_);
  or _50989_ (_18864_, _18863_, _18859_);
  or _50990_ (_18865_, _18864_, _02421_);
  and _50991_ (_18866_, _18865_, _02414_);
  and _50992_ (_18867_, _18866_, _18855_);
  or _50993_ (_18868_, _18867_, _18845_);
  and _50994_ (_18869_, _18868_, _02496_);
  or _50995_ (_18870_, _18869_, _18823_);
  and _50996_ (_18871_, _18870_, _02546_);
  or _50997_ (_18872_, _18871_, _18777_);
  and _50998_ (_18873_, _18872_, _02405_);
  or _50999_ (_18874_, _18873_, _18683_);
  and _51000_ (_18875_, _18874_, _26777_);
  and _51001_ (_18876_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and _51002_ (_18877_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or _51003_ (_18878_, _18877_, _18876_);
  and _51004_ (_18879_, _18878_, _02393_);
  and _51005_ (_18880_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and _51006_ (_18881_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or _51007_ (_18882_, _18881_, _18880_);
  and _51008_ (_18883_, _18882_, _02445_);
  or _51009_ (_18884_, _18883_, _18879_);
  and _51010_ (_18885_, _18884_, _02421_);
  and _51011_ (_18886_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  and _51012_ (_18887_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or _51013_ (_18888_, _18887_, _18886_);
  and _51014_ (_18889_, _18888_, _02393_);
  and _51015_ (_18890_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and _51016_ (_18891_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or _51017_ (_18892_, _18891_, _18890_);
  and _51018_ (_18893_, _18892_, _02445_);
  or _51019_ (_18894_, _18893_, _18889_);
  and _51020_ (_18895_, _18894_, _02459_);
  or _51021_ (_18896_, _18895_, _18885_);
  and _51022_ (_18897_, _18896_, _02458_);
  or _51023_ (_18898_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or _51024_ (_18899_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and _51025_ (_18900_, _18899_, _18898_);
  and _51026_ (_18901_, _18900_, _02393_);
  or _51027_ (_18902_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or _51028_ (_18903_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and _51029_ (_18904_, _18903_, _18902_);
  and _51030_ (_18905_, _18904_, _02445_);
  or _51031_ (_18906_, _18905_, _18901_);
  and _51032_ (_18907_, _18906_, _02421_);
  or _51033_ (_18908_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or _51034_ (_18909_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and _51035_ (_18910_, _18909_, _18908_);
  and _51036_ (_18911_, _18910_, _02393_);
  or _51037_ (_18912_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or _51038_ (_18913_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and _51039_ (_18914_, _18913_, _18912_);
  and _51040_ (_18915_, _18914_, _02445_);
  or _51041_ (_18916_, _18915_, _18911_);
  and _51042_ (_18917_, _18916_, _02459_);
  or _51043_ (_18918_, _18917_, _18907_);
  and _51044_ (_18919_, _18918_, _02414_);
  or _51045_ (_18920_, _18919_, _18897_);
  and _51046_ (_18921_, _18920_, _02398_);
  and _51047_ (_18922_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and _51048_ (_18923_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or _51049_ (_18924_, _18923_, _18922_);
  and _51050_ (_18925_, _18924_, _02393_);
  and _51051_ (_18926_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and _51052_ (_18927_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or _51053_ (_18928_, _18927_, _18926_);
  and _51054_ (_18929_, _18928_, _02445_);
  or _51055_ (_18930_, _18929_, _18925_);
  and _51056_ (_18931_, _18930_, _02421_);
  and _51057_ (_18932_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and _51058_ (_18933_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or _51059_ (_18934_, _18933_, _18932_);
  and _51060_ (_18935_, _18934_, _02393_);
  and _51061_ (_18936_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and _51062_ (_18937_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or _51063_ (_18938_, _18937_, _18936_);
  and _51064_ (_18939_, _18938_, _02445_);
  or _51065_ (_18940_, _18939_, _18935_);
  and _51066_ (_18941_, _18940_, _02459_);
  or _51067_ (_18942_, _18941_, _18931_);
  and _51068_ (_18943_, _18942_, _02458_);
  or _51069_ (_18944_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or _51070_ (_18945_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and _51071_ (_18946_, _18945_, _02445_);
  and _51072_ (_18947_, _18946_, _18944_);
  or _51073_ (_18948_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or _51074_ (_18949_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and _51075_ (_18950_, _18949_, _02393_);
  and _51076_ (_18951_, _18950_, _18948_);
  or _51077_ (_18952_, _18951_, _18947_);
  and _51078_ (_18953_, _18952_, _02421_);
  or _51079_ (_18954_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or _51080_ (_18955_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and _51081_ (_18956_, _18955_, _02445_);
  and _51082_ (_18957_, _18956_, _18954_);
  or _51083_ (_18958_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or _51084_ (_18959_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and _51085_ (_18960_, _18959_, _02393_);
  and _51086_ (_18961_, _18960_, _18958_);
  or _51087_ (_18962_, _18961_, _18957_);
  and _51088_ (_18963_, _18962_, _02459_);
  or _51089_ (_18964_, _18963_, _18953_);
  and _51090_ (_18965_, _18964_, _02414_);
  or _51091_ (_18966_, _18965_, _18943_);
  and _51092_ (_18967_, _18966_, _02496_);
  or _51093_ (_18968_, _18967_, _18921_);
  and _51094_ (_18969_, _18968_, _02400_);
  and _51095_ (_18970_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and _51096_ (_18971_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or _51097_ (_18972_, _18971_, _18970_);
  and _51098_ (_18973_, _18972_, _02393_);
  and _51099_ (_18974_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and _51100_ (_18975_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or _51101_ (_18976_, _18975_, _18974_);
  and _51102_ (_18977_, _18976_, _02445_);
  or _51103_ (_18978_, _18977_, _18973_);
  or _51104_ (_18979_, _18978_, _02459_);
  and _51105_ (_18980_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and _51106_ (_18981_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or _51107_ (_18982_, _18981_, _18980_);
  and _51108_ (_18983_, _18982_, _02393_);
  and _51109_ (_18984_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and _51110_ (_18985_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or _51111_ (_18986_, _18985_, _18984_);
  and _51112_ (_18987_, _18986_, _02445_);
  or _51113_ (_18988_, _18987_, _18983_);
  or _51114_ (_18989_, _18988_, _02421_);
  and _51115_ (_18990_, _18989_, _02458_);
  and _51116_ (_18991_, _18990_, _18979_);
  or _51117_ (_18992_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or _51118_ (_18993_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and _51119_ (_18994_, _18993_, _02445_);
  and _51120_ (_18995_, _18994_, _18992_);
  or _51121_ (_18996_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or _51122_ (_18997_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and _51123_ (_18998_, _18997_, _02393_);
  and _51124_ (_18999_, _18998_, _18996_);
  or _51125_ (_19000_, _18999_, _18995_);
  or _51126_ (_19001_, _19000_, _02459_);
  or _51127_ (_19002_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or _51128_ (_19003_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  and _51129_ (_19004_, _19003_, _02445_);
  and _51130_ (_19005_, _19004_, _19002_);
  or _51131_ (_19006_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or _51132_ (_19007_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  and _51133_ (_19008_, _19007_, _02393_);
  and _51134_ (_19009_, _19008_, _19006_);
  or _51135_ (_19010_, _19009_, _19005_);
  or _51136_ (_19011_, _19010_, _02421_);
  and _51137_ (_19012_, _19011_, _02414_);
  and _51138_ (_19013_, _19012_, _19001_);
  or _51139_ (_19014_, _19013_, _18991_);
  and _51140_ (_19015_, _19014_, _02496_);
  and _51141_ (_19016_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and _51142_ (_19017_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or _51143_ (_19018_, _19017_, _19016_);
  and _51144_ (_19019_, _19018_, _02393_);
  and _51145_ (_19020_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and _51146_ (_19021_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or _51147_ (_19022_, _19021_, _19020_);
  and _51148_ (_19023_, _19022_, _02445_);
  or _51149_ (_19024_, _19023_, _19019_);
  or _51150_ (_19025_, _19024_, _02459_);
  and _51151_ (_19026_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  and _51152_ (_19027_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or _51153_ (_19028_, _19027_, _19026_);
  and _51154_ (_19029_, _19028_, _02393_);
  and _51155_ (_19030_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and _51156_ (_19031_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or _51157_ (_19032_, _19031_, _19030_);
  and _51158_ (_19033_, _19032_, _02445_);
  or _51159_ (_19034_, _19033_, _19029_);
  or _51160_ (_19035_, _19034_, _02421_);
  and _51161_ (_19036_, _19035_, _02458_);
  and _51162_ (_19037_, _19036_, _19025_);
  or _51163_ (_19038_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or _51164_ (_19039_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and _51165_ (_19040_, _19039_, _19038_);
  and _51166_ (_19041_, _19040_, _02393_);
  or _51167_ (_19042_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or _51168_ (_19043_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and _51169_ (_19044_, _19043_, _19042_);
  and _51170_ (_19045_, _19044_, _02445_);
  or _51171_ (_19046_, _19045_, _19041_);
  or _51172_ (_19047_, _19046_, _02459_);
  or _51173_ (_19048_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or _51174_ (_19049_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and _51175_ (_19050_, _19049_, _19048_);
  and _51176_ (_19051_, _19050_, _02393_);
  or _51177_ (_19052_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or _51178_ (_19053_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  and _51179_ (_19054_, _19053_, _19052_);
  and _51180_ (_19055_, _19054_, _02445_);
  or _51181_ (_19056_, _19055_, _19051_);
  or _51182_ (_19057_, _19056_, _02421_);
  and _51183_ (_19058_, _19057_, _02414_);
  and _51184_ (_19059_, _19058_, _19047_);
  or _51185_ (_19060_, _19059_, _19037_);
  and _51186_ (_19061_, _19060_, _02398_);
  or _51187_ (_19062_, _19061_, _19015_);
  and _51188_ (_19063_, _19062_, _02546_);
  or _51189_ (_19064_, _19063_, _18969_);
  and _51190_ (_19065_, _19064_, _02646_);
  or _51191_ (_19066_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or _51192_ (_19067_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and _51193_ (_19068_, _19067_, _02445_);
  and _51194_ (_19069_, _19068_, _19066_);
  or _51195_ (_19070_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or _51196_ (_19071_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and _51197_ (_19072_, _19071_, _02393_);
  and _51198_ (_19073_, _19072_, _19070_);
  or _51199_ (_19074_, _19073_, _19069_);
  and _51200_ (_19075_, _19074_, _02459_);
  or _51201_ (_19076_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or _51202_ (_19077_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  and _51203_ (_19078_, _19077_, _02445_);
  and _51204_ (_19079_, _19078_, _19076_);
  or _51205_ (_19080_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or _51206_ (_19081_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and _51207_ (_19082_, _19081_, _02393_);
  and _51208_ (_19083_, _19082_, _19080_);
  or _51209_ (_19084_, _19083_, _19079_);
  and _51210_ (_19085_, _19084_, _02421_);
  or _51211_ (_19086_, _19085_, _19075_);
  and _51212_ (_19087_, _19086_, _02414_);
  and _51213_ (_19088_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  and _51214_ (_19089_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or _51215_ (_19090_, _19089_, _19088_);
  and _51216_ (_19091_, _19090_, _02393_);
  and _51217_ (_19092_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and _51218_ (_19093_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or _51219_ (_19094_, _19093_, _19092_);
  and _51220_ (_19095_, _19094_, _02445_);
  or _51221_ (_19096_, _19095_, _19091_);
  and _51222_ (_19097_, _19096_, _02459_);
  and _51223_ (_19098_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and _51224_ (_19099_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or _51225_ (_19100_, _19099_, _19098_);
  and _51226_ (_19101_, _19100_, _02393_);
  and _51227_ (_19102_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and _51228_ (_19103_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or _51229_ (_19104_, _19103_, _19102_);
  and _51230_ (_19105_, _19104_, _02445_);
  or _51231_ (_19106_, _19105_, _19101_);
  and _51232_ (_19107_, _19106_, _02421_);
  or _51233_ (_19108_, _19107_, _19097_);
  and _51234_ (_19109_, _19108_, _02458_);
  or _51235_ (_19110_, _19109_, _19087_);
  and _51236_ (_19111_, _19110_, _02496_);
  or _51237_ (_19112_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or _51238_ (_19113_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and _51239_ (_19114_, _19113_, _19112_);
  and _51240_ (_19115_, _19114_, _02393_);
  or _51241_ (_19116_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or _51242_ (_19117_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  and _51243_ (_19118_, _19117_, _19116_);
  and _51244_ (_19119_, _19118_, _02445_);
  or _51245_ (_19120_, _19119_, _19115_);
  and _51246_ (_19121_, _19120_, _02459_);
  or _51247_ (_19122_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or _51248_ (_19123_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and _51249_ (_19124_, _19123_, _19122_);
  and _51250_ (_19125_, _19124_, _02393_);
  or _51251_ (_19126_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or _51252_ (_19127_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and _51253_ (_19128_, _19127_, _19126_);
  and _51254_ (_19129_, _19128_, _02445_);
  or _51255_ (_19130_, _19129_, _19125_);
  and _51256_ (_19131_, _19130_, _02421_);
  or _51257_ (_19132_, _19131_, _19121_);
  and _51258_ (_19133_, _19132_, _02414_);
  and _51259_ (_19134_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and _51260_ (_19135_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or _51261_ (_19136_, _19135_, _19134_);
  and _51262_ (_19137_, _19136_, _02393_);
  and _51263_ (_19138_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and _51264_ (_19139_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or _51265_ (_19140_, _19139_, _19138_);
  and _51266_ (_19141_, _19140_, _02445_);
  or _51267_ (_19142_, _19141_, _19137_);
  and _51268_ (_19143_, _19142_, _02459_);
  and _51269_ (_19144_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  and _51270_ (_19145_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or _51271_ (_19146_, _19145_, _19144_);
  and _51272_ (_19147_, _19146_, _02393_);
  and _51273_ (_19148_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  and _51274_ (_19149_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or _51275_ (_19150_, _19149_, _19148_);
  and _51276_ (_19151_, _19150_, _02445_);
  or _51277_ (_19152_, _19151_, _19147_);
  and _51278_ (_19153_, _19152_, _02421_);
  or _51279_ (_19154_, _19153_, _19143_);
  and _51280_ (_19155_, _19154_, _02458_);
  or _51281_ (_19156_, _19155_, _19133_);
  and _51282_ (_19157_, _19156_, _02398_);
  or _51283_ (_19158_, _19157_, _19111_);
  and _51284_ (_19159_, _19158_, _02400_);
  and _51285_ (_19160_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and _51286_ (_19161_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or _51287_ (_19162_, _19161_, _19160_);
  and _51288_ (_19163_, _19162_, _02393_);
  and _51289_ (_19164_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and _51290_ (_19165_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or _51291_ (_19166_, _19165_, _19164_);
  and _51292_ (_19167_, _19166_, _02445_);
  or _51293_ (_19168_, _19167_, _19163_);
  or _51294_ (_19169_, _19168_, _02459_);
  and _51295_ (_19170_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and _51296_ (_19171_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or _51297_ (_19172_, _19171_, _19170_);
  and _51298_ (_19173_, _19172_, _02393_);
  and _51299_ (_19174_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and _51300_ (_19175_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or _51301_ (_19176_, _19175_, _19174_);
  and _51302_ (_19177_, _19176_, _02445_);
  or _51303_ (_19178_, _19177_, _19173_);
  or _51304_ (_19179_, _19178_, _02421_);
  and _51305_ (_19180_, _19179_, _02458_);
  and _51306_ (_19181_, _19180_, _19169_);
  or _51307_ (_19182_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or _51308_ (_19183_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and _51309_ (_19184_, _19183_, _19182_);
  and _51310_ (_19185_, _19184_, _02393_);
  or _51311_ (_19186_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or _51312_ (_19187_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and _51313_ (_19188_, _19187_, _19186_);
  and _51314_ (_19189_, _19188_, _02445_);
  or _51315_ (_19190_, _19189_, _19185_);
  or _51316_ (_19191_, _19190_, _02459_);
  or _51317_ (_19192_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or _51318_ (_19193_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and _51319_ (_19194_, _19193_, _19192_);
  and _51320_ (_19195_, _19194_, _02393_);
  or _51321_ (_19196_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or _51322_ (_19197_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and _51323_ (_19198_, _19197_, _19196_);
  and _51324_ (_19199_, _19198_, _02445_);
  or _51325_ (_19200_, _19199_, _19195_);
  or _51326_ (_19201_, _19200_, _02421_);
  and _51327_ (_19202_, _19201_, _02414_);
  and _51328_ (_19203_, _19202_, _19191_);
  or _51329_ (_19204_, _19203_, _19181_);
  and _51330_ (_19205_, _19204_, _02398_);
  and _51331_ (_19206_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  and _51332_ (_19207_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or _51333_ (_19208_, _19207_, _19206_);
  and _51334_ (_19209_, _19208_, _02393_);
  and _51335_ (_19210_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and _51336_ (_19211_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or _51337_ (_19212_, _19211_, _19210_);
  and _51338_ (_19213_, _19212_, _02445_);
  or _51339_ (_19214_, _19213_, _19209_);
  or _51340_ (_19215_, _19214_, _02459_);
  and _51341_ (_19216_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  and _51342_ (_19217_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or _51343_ (_19218_, _19217_, _19216_);
  and _51344_ (_19219_, _19218_, _02393_);
  and _51345_ (_19220_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and _51346_ (_19221_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or _51347_ (_19222_, _19221_, _19220_);
  and _51348_ (_19223_, _19222_, _02445_);
  or _51349_ (_19224_, _19223_, _19219_);
  or _51350_ (_19225_, _19224_, _02421_);
  and _51351_ (_19226_, _19225_, _02458_);
  and _51352_ (_19227_, _19226_, _19215_);
  or _51353_ (_19228_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or _51354_ (_19229_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and _51355_ (_19230_, _19229_, _02445_);
  and _51356_ (_19231_, _19230_, _19228_);
  or _51357_ (_19232_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or _51358_ (_19233_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  and _51359_ (_19234_, _19233_, _02393_);
  and _51360_ (_19235_, _19234_, _19232_);
  or _51361_ (_19236_, _19235_, _19231_);
  or _51362_ (_19237_, _19236_, _02459_);
  or _51363_ (_19238_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or _51364_ (_19239_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and _51365_ (_19240_, _19239_, _02445_);
  and _51366_ (_19241_, _19240_, _19238_);
  or _51367_ (_19242_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or _51368_ (_19243_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  and _51369_ (_19244_, _19243_, _02393_);
  and _51370_ (_19245_, _19244_, _19242_);
  or _51371_ (_19246_, _19245_, _19241_);
  or _51372_ (_19247_, _19246_, _02421_);
  and _51373_ (_19248_, _19247_, _02414_);
  and _51374_ (_19249_, _19248_, _19237_);
  or _51375_ (_19250_, _19249_, _19227_);
  and _51376_ (_19251_, _19250_, _02496_);
  or _51377_ (_19252_, _19251_, _19205_);
  and _51378_ (_19253_, _19252_, _02546_);
  or _51379_ (_19254_, _19253_, _19159_);
  and _51380_ (_19255_, _19254_, _02405_);
  or _51381_ (_19256_, _19255_, _19065_);
  and _51382_ (_19257_, _19256_, _02444_);
  or _51383_ (_19258_, _19257_, _18875_);
  or _51384_ (_19259_, _19258_, _02443_);
  or _51385_ (_19260_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and _51386_ (_19261_, _19260_, _22762_);
  and _51387_ (_11175_, _19261_, _19259_);
  and _51388_ (_19262_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  and _51389_ (_19263_, _24222_, _23898_);
  or _51390_ (_11183_, _19263_, _19262_);
  and _51391_ (_19264_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  and _51392_ (_19265_, _24222_, _23778_);
  or _51393_ (_11189_, _19265_, _19264_);
  and _51394_ (_19266_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  and _51395_ (_19267_, _17775_, _23747_);
  or _51396_ (_11193_, _19267_, _19266_);
  and _51397_ (_19268_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  and _51398_ (_19269_, _16371_, _23778_);
  or _51399_ (_11195_, _19269_, _19268_);
  and _51400_ (_19270_, _18167_, _23649_);
  and _51401_ (_19271_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  or _51402_ (_11200_, _19271_, _19270_);
  and _51403_ (_19272_, _18167_, _23747_);
  and _51404_ (_19273_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  or _51405_ (_11203_, _19273_, _19272_);
  and _51406_ (_19274_, _18167_, _23824_);
  and _51407_ (_19275_, _18169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  or _51408_ (_27221_, _19275_, _19274_);
  and _51409_ (_19276_, _06552_, _24050_);
  and _51410_ (_19277_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or _51411_ (_11207_, _19277_, _19276_);
  and _51412_ (_19278_, _16372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  and _51413_ (_19279_, _16371_, _23898_);
  or _51414_ (_26972_, _19279_, _19278_);
  and _51415_ (_19280_, _06552_, _23946_);
  and _51416_ (_19281_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or _51417_ (_11216_, _19281_, _19280_);
  and _51418_ (_19282_, _18217_, _23707_);
  and _51419_ (_19283_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or _51420_ (_11222_, _19283_, _19282_);
  and _51421_ (_19284_, _17215_, _23898_);
  and _51422_ (_19285_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  or _51423_ (_11228_, _19285_, _19284_);
  and _51424_ (_19286_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and _51425_ (_19287_, _17255_, _24050_);
  or _51426_ (_11230_, _19287_, _19286_);
  and _51427_ (_19288_, _17215_, _23778_);
  and _51428_ (_19289_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  or _51429_ (_11236_, _19289_, _19288_);
  and _51430_ (_19290_, _24006_, _23649_);
  and _51431_ (_19291_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  or _51432_ (_11242_, _19291_, _19290_);
  and _51433_ (_19292_, _23946_, _23790_);
  and _51434_ (_19293_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or _51435_ (_11244_, _19293_, _19292_);
  and _51436_ (_19294_, _02241_, _23898_);
  and _51437_ (_19295_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or _51438_ (_11246_, _19295_, _19294_);
  and _51439_ (_19296_, _24050_, _23987_);
  and _51440_ (_19297_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  or _51441_ (_26937_, _19297_, _19296_);
  and _51442_ (_19298_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and _51443_ (_19299_, _13763_, _23898_);
  or _51444_ (_27243_, _19299_, _19298_);
  and _51445_ (_19300_, _23987_, _23649_);
  and _51446_ (_19301_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  or _51447_ (_11252_, _19301_, _19300_);
  and _51448_ (_19302_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and _51449_ (_19303_, _13763_, _23778_);
  or _51450_ (_11255_, _19303_, _19302_);
  and _51451_ (_19304_, _02241_, _23778_);
  and _51452_ (_19305_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or _51453_ (_11258_, _19305_, _19304_);
  and _51454_ (_19306_, _23898_, _23790_);
  and _51455_ (_19307_, _23827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  or _51456_ (_11262_, _19307_, _19306_);
  and _51457_ (_19308_, _06552_, _23707_);
  and _51458_ (_19309_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or _51459_ (_11265_, _19309_, _19308_);
  and _51460_ (_19310_, _02326_, _23747_);
  and _51461_ (_19311_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or _51462_ (_11267_, _19311_, _19310_);
  and _51463_ (_19312_, _02241_, _23824_);
  and _51464_ (_19313_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or _51465_ (_27292_, _19313_, _19312_);
  and _51466_ (_19314_, _07743_, _23946_);
  and _51467_ (_19315_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or _51468_ (_11270_, _19315_, _19314_);
  and _51469_ (_19316_, _24086_, _23747_);
  and _51470_ (_19317_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or _51471_ (_11273_, _19317_, _19316_);
  and _51472_ (_19318_, _23987_, _23946_);
  and _51473_ (_19319_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  or _51474_ (_26936_, _19319_, _19318_);
  and _51475_ (_19320_, _01971_, _23707_);
  and _51476_ (_19321_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or _51477_ (_11280_, _19321_, _19320_);
  and _51478_ (_19322_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  and _51479_ (_19323_, _16319_, _23747_);
  or _51480_ (_11286_, _19323_, _19322_);
  and _51481_ (_19324_, _23907_, _23778_);
  and _51482_ (_19325_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or _51483_ (_11289_, _19325_, _19324_);
  and _51484_ (_19326_, _23907_, _23824_);
  and _51485_ (_19327_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or _51486_ (_11296_, _19327_, _19326_);
  and _51487_ (_19328_, _23912_, _23649_);
  and _51488_ (_19329_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  or _51489_ (_11299_, _19329_, _19328_);
  and _51490_ (_19330_, _02241_, _23946_);
  and _51491_ (_19331_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or _51492_ (_11307_, _19331_, _19330_);
  and _51493_ (_19332_, _02241_, _23707_);
  and _51494_ (_19333_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or _51495_ (_11312_, _19333_, _19332_);
  and _51496_ (_19334_, _24006_, _23778_);
  and _51497_ (_19335_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  or _51498_ (_11315_, _19335_, _19334_);
  and _51499_ (_19336_, _24006_, _23824_);
  and _51500_ (_19337_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  or _51501_ (_11317_, _19337_, _19336_);
  and _51502_ (_19338_, _23987_, _23707_);
  and _51503_ (_19339_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  or _51504_ (_11319_, _19339_, _19338_);
  and _51505_ (_19340_, _24086_, _24050_);
  and _51506_ (_19341_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or _51507_ (_27256_, _19341_, _19340_);
  and _51508_ (_19342_, _24011_, _23946_);
  and _51509_ (_19343_, _24013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or _51510_ (_11322_, _19343_, _19342_);
  and _51511_ (_19344_, _02241_, _23649_);
  and _51512_ (_19345_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or _51513_ (_27294_, _19345_, _19344_);
  and _51514_ (_19346_, _24006_, _23898_);
  and _51515_ (_19347_, _24008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  or _51516_ (_11329_, _19347_, _19346_);
  and _51517_ (_19348_, _02241_, _24050_);
  and _51518_ (_19349_, _02243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or _51519_ (_11331_, _19349_, _19348_);
  and _51520_ (_19350_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and _51521_ (_19351_, _07513_, _23747_);
  or _51522_ (_11335_, _19351_, _19350_);
  and _51523_ (_19352_, _23912_, _23778_);
  and _51524_ (_19353_, _23948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  or _51525_ (_11341_, _19353_, _19352_);
  and _51526_ (_19354_, _24050_, _23907_);
  and _51527_ (_19355_, _23909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or _51528_ (_11346_, _19355_, _19354_);
  and _51529_ (_19356_, _23992_, _23898_);
  and _51530_ (_19357_, _23994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or _51531_ (_11349_, _19357_, _19356_);
  and _51532_ (_19358_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and _51533_ (_19359_, _13763_, _23649_);
  or _51534_ (_27244_, _19359_, _19358_);
  and _51535_ (_19360_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  and _51536_ (_19361_, _24203_, _23898_);
  or _51537_ (_11353_, _19361_, _19360_);
  and _51538_ (_19362_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and _51539_ (_19363_, _24276_, _24050_);
  or _51540_ (_27251_, _19363_, _19362_);
  and _51541_ (_19364_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and _51542_ (_19365_, _24276_, _23778_);
  or _51543_ (_11356_, _19365_, _19364_);
  and _51544_ (_19366_, _01971_, _24050_);
  and _51545_ (_19367_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  or _51546_ (_11358_, _19367_, _19366_);
  and _51547_ (_19368_, _17378_, _23649_);
  and _51548_ (_19369_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  or _51549_ (_27291_, _19369_, _19368_);
  and _51550_ (_19370_, _17378_, _24050_);
  and _51551_ (_19371_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  or _51552_ (_11364_, _19371_, _19370_);
  and _51553_ (_19372_, _13764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  and _51554_ (_19373_, _13763_, _23747_);
  or _51555_ (_11368_, _19373_, _19372_);
  and _51556_ (_19374_, _23987_, _23898_);
  and _51557_ (_19375_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  or _51558_ (_11374_, _19375_, _19374_);
  and _51559_ (_19376_, _23987_, _23824_);
  and _51560_ (_19377_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  or _51561_ (_11376_, _19377_, _19376_);
  and _51562_ (_19378_, _17378_, _23707_);
  and _51563_ (_19379_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or _51564_ (_11388_, _19379_, _19378_);
  and _51565_ (_19380_, _24277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  and _51566_ (_19381_, _24276_, _23747_);
  or _51567_ (_11394_, _19381_, _19380_);
  and _51568_ (_19382_, _01971_, _23946_);
  and _51569_ (_19383_, _01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or _51570_ (_11396_, _19383_, _19382_);
  and _51571_ (_19384_, _17535_, _23707_);
  and _51572_ (_19385_, _17537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or _51573_ (_26935_, _19385_, _19384_);
  and _51574_ (_19386_, _07743_, _23649_);
  and _51575_ (_19387_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  or _51576_ (_11400_, _19387_, _19386_);
  and _51577_ (_19388_, _17378_, _23747_);
  and _51578_ (_19389_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  or _51579_ (_27290_, _19389_, _19388_);
  and _51580_ (_19390_, _24223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  and _51581_ (_19391_, _24222_, _24050_);
  or _51582_ (_11404_, _19391_, _19390_);
  and _51583_ (_19392_, _23987_, _23778_);
  and _51584_ (_19393_, _23989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  or _51585_ (_11406_, _19393_, _19392_);
  and _51586_ (_19394_, _17378_, _23946_);
  and _51587_ (_19395_, _17380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  or _51588_ (_11408_, _19395_, _19394_);
  and _51589_ (_19396_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  and _51590_ (_19397_, _16018_, _24050_);
  or _51591_ (_11410_, _19397_, _19396_);
  and _51592_ (_19398_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  and _51593_ (_19399_, _16319_, _23946_);
  or _51594_ (_11414_, _19399_, _19398_);
  and _51595_ (_19400_, _24204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  and _51596_ (_19401_, _24203_, _23649_);
  or _51597_ (_11418_, _19401_, _19400_);
  and _51598_ (_19402_, _17221_, _23747_);
  and _51599_ (_19403_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or _51600_ (_11425_, _19403_, _19402_);
  and _51601_ (_19404_, _06552_, _23747_);
  and _51602_ (_19405_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or _51603_ (_27144_, _19405_, _19404_);
  and _51604_ (_19406_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  and _51605_ (_19407_, _16018_, _23649_);
  or _51606_ (_26965_, _19407_, _19406_);
  and _51607_ (_19408_, _17215_, _23824_);
  and _51608_ (_19409_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  or _51609_ (_27217_, _19409_, _19408_);
  and _51610_ (_19410_, _06552_, _23824_);
  and _51611_ (_19411_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or _51612_ (_11454_, _19411_, _19410_);
  and _51613_ (_19412_, _25156_, _23946_);
  and _51614_ (_19413_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or _51615_ (_11456_, _19413_, _19412_);
  and _51616_ (_19414_, _25156_, _23747_);
  and _51617_ (_19415_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or _51618_ (_11458_, _19415_, _19414_);
  and _51619_ (_19416_, _25091_, _24050_);
  and _51620_ (_19417_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  or _51621_ (_11460_, _19417_, _19416_);
  and _51622_ (_19418_, _25091_, _23649_);
  and _51623_ (_19419_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  or _51624_ (_11463_, _19419_, _19418_);
  and _51625_ (_19420_, _17215_, _23649_);
  and _51626_ (_19422_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  or _51627_ (_11468_, _19422_, _19420_);
  and _51628_ (_19423_, _25079_, _23747_);
  and _51629_ (_19424_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  or _51630_ (_11471_, _19424_, _19423_);
  and _51631_ (_19425_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and _51632_ (_19426_, _17091_, _23747_);
  or _51633_ (_11473_, _19426_, _19425_);
  and _51634_ (_19427_, _24999_, _23649_);
  and _51635_ (_19428_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or _51636_ (_27184_, _19428_, _19427_);
  and _51637_ (_19429_, _24932_, _23649_);
  and _51638_ (_19430_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or _51639_ (_11478_, _19430_, _19429_);
  and _51640_ (_19431_, _24932_, _23778_);
  and _51641_ (_19432_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or _51642_ (_27179_, _19432_, _19431_);
  and _51643_ (_19433_, _08198_, _24050_);
  and _51644_ (_19434_, _08200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or _51645_ (_11483_, _19434_, _19433_);
  and _51646_ (_19435_, _24858_, _23946_);
  and _51647_ (_19436_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  or _51648_ (_11485_, _19436_, _19435_);
  and _51649_ (_19437_, _24858_, _23824_);
  and _51650_ (_19438_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  or _51651_ (_11487_, _19438_, _19437_);
  and _51652_ (_19439_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  and _51653_ (_19440_, _17091_, _23824_);
  or _51654_ (_11489_, _19440_, _19439_);
  and _51655_ (_19441_, _24839_, _23707_);
  and _51656_ (_19442_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  or _51657_ (_11491_, _19442_, _19441_);
  and _51658_ (_19443_, _24839_, _23747_);
  and _51659_ (_19444_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  or _51660_ (_11493_, _19444_, _19443_);
  and _51661_ (_19445_, _17215_, _23747_);
  and _51662_ (_19446_, _17217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  or _51663_ (_11497_, _19446_, _19445_);
  and _51664_ (_19447_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and _51665_ (_19448_, _16375_, _23707_);
  or _51666_ (_11499_, _19448_, _19447_);
  and _51667_ (_19449_, _24789_, _23946_);
  and _51668_ (_19450_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or _51669_ (_11502_, _19450_, _19449_);
  and _51670_ (_19451_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and _51671_ (_19452_, _16375_, _24050_);
  or _51672_ (_26970_, _19452_, _19451_);
  and _51673_ (_19453_, _24789_, _23898_);
  and _51674_ (_19454_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or _51675_ (_11505_, _19454_, _19453_);
  and _51676_ (_19455_, _24722_, _24050_);
  and _51677_ (_19456_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  or _51678_ (_11506_, _19456_, _19455_);
  and _51679_ (_19457_, _24722_, _23824_);
  and _51680_ (_19458_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  or _51681_ (_11510_, _19458_, _19457_);
  and _51682_ (_19459_, _24121_, _23816_);
  nor _51683_ (_19460_, _14722_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _51684_ (_19461_, _19460_, _14723_);
  nand _51685_ (_19462_, _19461_, _24174_);
  or _51686_ (_19463_, _24174_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _51687_ (_19464_, _19463_, _19462_);
  nand _51688_ (_19465_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _51689_ (_19466_, _19465_, _24127_);
  or _51690_ (_19467_, _19466_, _19464_);
  and _51691_ (_19468_, _19467_, _24166_);
  or _51692_ (_11512_, _19468_, _19459_);
  and _51693_ (_19469_, _07743_, _23747_);
  and _51694_ (_19470_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  or _51695_ (_11515_, _19470_, _19469_);
  and _51696_ (_19471_, _24688_, _24050_);
  and _51697_ (_19472_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  or _51698_ (_11519_, _19472_, _19471_);
  and _51699_ (_19473_, _24688_, _23824_);
  and _51700_ (_19474_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  or _51701_ (_11522_, _19474_, _19473_);
  and _51702_ (_19475_, _24688_, _23778_);
  and _51703_ (_19476_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  or _51704_ (_11524_, _19476_, _19475_);
  and _51705_ (_19477_, _17221_, _23824_);
  and _51706_ (_19478_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or _51707_ (_11526_, _19478_, _19477_);
  and _51708_ (_19479_, _24639_, _23707_);
  and _51709_ (_19480_, _24641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or _51710_ (_11528_, _19480_, _19479_);
  and _51711_ (_19481_, _24375_, _23649_);
  and _51712_ (_19482_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or _51713_ (_11532_, _19482_, _19481_);
  and _51714_ (_19483_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and _51715_ (_19484_, _17091_, _24050_);
  or _51716_ (_11534_, _19484_, _19483_);
  and _51717_ (_19485_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and _51718_ (_19486_, _01967_, _23649_);
  or _51719_ (_11538_, _19486_, _19485_);
  and _51720_ (_19487_, _25091_, _23778_);
  and _51721_ (_19488_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  or _51722_ (_11539_, _19488_, _19487_);
  and _51723_ (_19489_, _25079_, _23946_);
  and _51724_ (_19490_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  or _51725_ (_11541_, _19490_, _19489_);
  and _51726_ (_19491_, _25079_, _23898_);
  and _51727_ (_19492_, _25081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  or _51728_ (_11543_, _19492_, _19491_);
  and _51729_ (_19493_, _24999_, _24050_);
  and _51730_ (_19494_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or _51731_ (_11545_, _19494_, _19493_);
  and _51732_ (_19495_, _24999_, _23898_);
  and _51733_ (_19496_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or _51734_ (_11548_, _19496_, _19495_);
  and _51735_ (_19497_, _24932_, _24050_);
  and _51736_ (_19498_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or _51737_ (_27181_, _19498_, _19497_);
  and _51738_ (_19499_, _24932_, _23824_);
  and _51739_ (_19500_, _24934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or _51740_ (_27180_, _19500_, _19499_);
  and _51741_ (_19501_, _24858_, _23707_);
  and _51742_ (_19502_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  or _51743_ (_11562_, _19502_, _19501_);
  and _51744_ (_19503_, _24950_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _51745_ (_19504_, _24865_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _51746_ (_19505_, _24865_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _51747_ (_19506_, _19505_, _19504_);
  nor _51748_ (_19507_, _19506_, _02137_);
  or _51749_ (_19508_, _19507_, _24862_);
  or _51750_ (_19509_, _19508_, _19503_);
  or _51751_ (_19510_, _19506_, _24954_);
  and _51752_ (_19511_, _19510_, _22762_);
  and _51753_ (_11565_, _19511_, _19509_);
  and _51754_ (_19512_, _15004_, _23778_);
  and _51755_ (_19513_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or _51756_ (_11568_, _19513_, _19512_);
  and _51757_ (_19514_, _24839_, _23778_);
  and _51758_ (_19515_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  or _51759_ (_11569_, _19515_, _19514_);
  and _51760_ (_19516_, _24645_, _24076_);
  and _51761_ (_19517_, _19516_, _24064_);
  nand _51762_ (_19518_, _19517_, _23711_);
  or _51763_ (_19519_, _25039_, _24961_);
  and _51764_ (_19520_, _19519_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and _51765_ (_19521_, _19520_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and _51766_ (_19522_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _24865_);
  and _51767_ (_19523_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _51768_ (_19524_, _19523_, _19522_);
  nor _51769_ (_19525_, _19524_, _24864_);
  nor _51770_ (_19526_, _02156_, _02121_);
  nor _51771_ (_19527_, _19526_, _24864_);
  nor _51772_ (_19528_, _19527_, _19525_);
  nand _51773_ (_19529_, _19528_, _19521_);
  nand _51774_ (_19530_, _19529_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _51775_ (_19531_, _19530_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _51776_ (_19532_, _19531_, _19517_);
  and _51777_ (_19533_, _19532_, _19518_);
  nand _51778_ (_19534_, _19533_, _24817_);
  or _51779_ (_19535_, _24817_, _23892_);
  and _51780_ (_19536_, _19535_, _22762_);
  and _51781_ (_11577_, _19536_, _19534_);
  and _51782_ (_19537_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and _51783_ (_19538_, _17091_, _23946_);
  or _51784_ (_11591_, _19538_, _19537_);
  and _51785_ (_19539_, _06552_, _23649_);
  and _51786_ (_19540_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or _51787_ (_11595_, _19540_, _19539_);
  and _51788_ (_11604_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _22762_);
  and _51789_ (_19541_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and _51790_ (_19542_, _17091_, _23649_);
  or _51791_ (_27242_, _19542_, _19541_);
  and _51792_ (_19543_, _24688_, _23649_);
  and _51793_ (_19544_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  or _51794_ (_11609_, _19544_, _19543_);
  and _51795_ (_19545_, _24375_, _23898_);
  and _51796_ (_19546_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or _51797_ (_11613_, _19546_, _19545_);
  and _51798_ (_19547_, _25156_, _23707_);
  and _51799_ (_19548_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or _51800_ (_11615_, _19548_, _19547_);
  and _51801_ (_19549_, _25156_, _23778_);
  and _51802_ (_19550_, _25158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or _51803_ (_11617_, _19550_, _19549_);
  and _51804_ (_19551_, _24858_, _23747_);
  and _51805_ (_19552_, _24860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  or _51806_ (_11621_, _19552_, _19551_);
  and _51807_ (_19553_, _24839_, _23649_);
  and _51808_ (_19554_, _24841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  or _51809_ (_11622_, _19554_, _19553_);
  and _51810_ (_19555_, _24789_, _23824_);
  and _51811_ (_19556_, _24791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or _51812_ (_11625_, _19556_, _19555_);
  and _51813_ (_19557_, _24722_, _23747_);
  and _51814_ (_19558_, _24724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  or _51815_ (_27174_, _19558_, _19557_);
  and _51816_ (_19559_, _24375_, _23946_);
  and _51817_ (_19560_, _24377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or _51818_ (_11628_, _19560_, _19559_);
  and _51819_ (_19561_, _25091_, _23898_);
  and _51820_ (_19562_, _25093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  or _51821_ (_27186_, _19562_, _19561_);
  and _51822_ (_19563_, _24999_, _23824_);
  and _51823_ (_19564_, _25001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or _51824_ (_27182_, _19564_, _19563_);
  not _51825_ (_19565_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _51826_ (_19566_, _19520_, _19565_);
  nand _51827_ (_19567_, _19526_, _19525_);
  or _51828_ (_19568_, _19567_, _19566_);
  and _51829_ (_19569_, _19568_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _51830_ (_19570_, _19569_, _06778_);
  and _51831_ (_19571_, _24813_, _24654_);
  or _51832_ (_19572_, _19571_, _19570_);
  nand _51833_ (_19573_, _19571_, _23594_);
  and _51834_ (_19574_, _19573_, _19572_);
  or _51835_ (_19575_, _19574_, _24816_);
  nand _51836_ (_19576_, _24816_, _23702_);
  and _51837_ (_19577_, _19576_, _22762_);
  and _51838_ (_11637_, _19577_, _19575_);
  and _51839_ (_11643_, _26274_, _22762_);
  and _51840_ (_19578_, _16320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  and _51841_ (_19579_, _16319_, _23778_);
  or _51842_ (_11645_, _19579_, _19578_);
  nand _51843_ (_19580_, _23018_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _51844_ (_19581_, _19580_, _24653_);
  or _51845_ (_19582_, _19581_, _05827_);
  and _51846_ (_19583_, _19582_, _24813_);
  nand _51847_ (_19584_, _24813_, _23018_);
  and _51848_ (_19585_, _19584_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _51849_ (_19586_, _19585_, _24816_);
  or _51850_ (_19587_, _19586_, _19583_);
  or _51851_ (_19588_, _24817_, _24043_);
  and _51852_ (_19589_, _19588_, _22762_);
  and _51853_ (_11651_, _19589_, _19587_);
  and _51854_ (_19590_, _24892_, _24880_);
  nand _51855_ (_19591_, _24895_, _19590_);
  nand _51856_ (_19592_, _24905_, _24902_);
  and _51857_ (_19593_, _19592_, _24896_);
  or _51858_ (_19594_, _19593_, _24895_);
  and _51859_ (_19595_, _19594_, _24938_);
  and _51860_ (_19596_, _19595_, _19591_);
  or _51861_ (_19597_, _19596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not _51862_ (_19598_, _24938_);
  not _51863_ (_19599_, _24918_);
  or _51864_ (_19600_, _19599_, _24914_);
  or _51865_ (_19601_, _24889_, _24870_);
  and _51866_ (_19602_, _19601_, _19600_);
  or _51867_ (_19603_, _19602_, _19598_);
  and _51868_ (_19604_, _19603_, _22762_);
  and _51869_ (_11656_, _19604_, _19597_);
  and _51870_ (_19605_, _04922_, _23778_);
  and _51871_ (_19606_, _04925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  or _51872_ (_11659_, _19606_, _19605_);
  and _51873_ (_11662_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _22762_);
  and _51874_ (_19607_, _19594_, _24863_);
  and _51875_ (_19608_, _19607_, _19591_);
  or _51876_ (_19609_, _19608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  not _51877_ (_19610_, _24863_);
  or _51878_ (_19611_, _19602_, _19610_);
  and _51879_ (_19612_, _19611_, _22762_);
  and _51880_ (_11663_, _19612_, _19609_);
  and _51881_ (_11665_, _26366_, _22762_);
  and _51882_ (_19613_, _25142_, _23707_);
  and _51883_ (_19614_, _25144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or _51884_ (_27201_, _19614_, _19613_);
  not _51885_ (_19615_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and _51886_ (_19616_, _19615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  not _51887_ (_19617_, _19525_);
  and _51888_ (_19618_, _19527_, _19617_);
  not _51889_ (_19619_, _19618_);
  or _51890_ (_19620_, _19619_, _19566_);
  and _51891_ (_19621_, _19620_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _51892_ (_19622_, _19621_, _19616_);
  and _51893_ (_19623_, _24813_, _24125_);
  or _51894_ (_19624_, _19623_, _19622_);
  nand _51895_ (_19625_, _19623_, _23594_);
  and _51896_ (_19626_, _19625_, _19624_);
  or _51897_ (_19627_, _19626_, _24816_);
  or _51898_ (_19628_, _24817_, _23939_);
  and _51899_ (_19629_, _19628_, _22762_);
  and _51900_ (_11677_, _19629_, _19627_);
  nand _51901_ (_19630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _51902_ (_19631_, _19618_, _19521_);
  nor _51903_ (_19632_, _19631_, _19630_);
  and _51904_ (_19633_, _24118_, _23003_);
  and _51905_ (_19634_, _19633_, _24064_);
  nand _51906_ (_19635_, _24645_, _19634_);
  nand _51907_ (_19636_, _19635_, _19632_);
  or _51908_ (_19637_, _19635_, _23594_);
  and _51909_ (_19638_, _19637_, _19636_);
  nand _51910_ (_19639_, _19638_, _24817_);
  or _51911_ (_19640_, _24817_, _23738_);
  and _51912_ (_19641_, _19640_, _22762_);
  and _51913_ (_11683_, _19641_, _19639_);
  and _51914_ (_19642_, _16019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  and _51915_ (_19643_, _16018_, _23946_);
  or _51916_ (_11684_, _19643_, _19642_);
  and _51917_ (_19644_, _24654_, _24648_);
  nand _51918_ (_19645_, _19644_, _23594_);
  or _51919_ (_19646_, _19644_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _51920_ (_19647_, _19646_, _24659_);
  and _51921_ (_19648_, _19647_, _19645_);
  nor _51922_ (_19649_, _24659_, _23702_);
  or _51923_ (_19650_, _19649_, _19648_);
  and _51924_ (_11687_, _19650_, _22762_);
  nor _51925_ (_19651_, _14721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _51926_ (_19652_, _19651_, _14722_);
  and _51927_ (_19653_, _19652_, _24174_);
  and _51928_ (_19654_, _14719_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand _51929_ (_19655_, _24185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _51930_ (_19656_, _19655_, _24127_);
  or _51931_ (_19657_, _19656_, _19654_);
  or _51932_ (_19658_, _19657_, _19653_);
  and _51933_ (_19659_, _19658_, _24171_);
  and _51934_ (_19660_, _24120_, _23892_);
  or _51935_ (_19661_, _19660_, _19659_);
  and _51936_ (_11690_, _19661_, _22762_);
  and _51937_ (_19662_, _17221_, _23898_);
  and _51938_ (_19663_, _17223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or _51939_ (_11694_, _19663_, _19662_);
  and _51940_ (_19664_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  and _51941_ (_19665_, _02306_, _24050_);
  or _51942_ (_11696_, _19665_, _19664_);
  and _51943_ (_19666_, _05119_, _23747_);
  and _51944_ (_19667_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  or _51945_ (_11698_, _19667_, _19666_);
  nand _51946_ (_19668_, _24950_, _24864_);
  nand _51947_ (_19669_, _19504_, _24862_);
  and _51948_ (_19670_, _19669_, _22762_);
  and _51949_ (_11704_, _19670_, _19668_);
  and _51950_ (_19671_, _25754_, _23778_);
  and _51951_ (_19672_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  or _51952_ (_27033_, _19672_, _19671_);
  and _51953_ (_19673_, _01759_, _23747_);
  and _51954_ (_19674_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or _51955_ (_11707_, _19674_, _19673_);
  and _51956_ (_19675_, _24730_, _24654_);
  nand _51957_ (_19676_, _19675_, _23594_);
  or _51958_ (_19677_, _19675_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _51959_ (_19678_, _19677_, _19676_);
  or _51960_ (_19679_, _19678_, _24736_);
  nand _51961_ (_19680_, _24736_, _23702_);
  and _51962_ (_19681_, _19680_, _22762_);
  and _51963_ (_11710_, _19681_, _19679_);
  and _51964_ (_19682_, _02215_, _24050_);
  and _51965_ (_19683_, _02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or _51966_ (_11711_, _19683_, _19682_);
  and _51967_ (_19684_, _02350_, _23824_);
  and _51968_ (_19685_, _02352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or _51969_ (_11715_, _19685_, _19684_);
  and _51970_ (_19686_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  and _51971_ (_19687_, _02306_, _23946_);
  or _51972_ (_11718_, _19687_, _19686_);
  and _51973_ (_19688_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  and _51974_ (_19689_, _02306_, _23649_);
  or _51975_ (_11721_, _19689_, _19688_);
  and _51976_ (_19690_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and _51977_ (_19691_, _16375_, _23824_);
  or _51978_ (_11723_, _19691_, _19690_);
  and _51979_ (_19692_, _08642_, _23707_);
  and _51980_ (_19693_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  or _51981_ (_11724_, _19693_, _19692_);
  and _51982_ (_19694_, _05298_, _23898_);
  and _51983_ (_19695_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or _51984_ (_11726_, _19695_, _19694_);
  and _51985_ (_19696_, _05346_, _23649_);
  and _51986_ (_19697_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or _51987_ (_11728_, _19697_, _19696_);
  and _51988_ (_19698_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and _51989_ (_19699_, _16375_, _23747_);
  or _51990_ (_26969_, _19699_, _19698_);
  and _51991_ (_19700_, _08642_, _24050_);
  and _51992_ (_19701_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  or _51993_ (_11733_, _19701_, _19700_);
  and _51994_ (_19702_, _05429_, _23898_);
  and _51995_ (_19703_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or _51996_ (_11734_, _19703_, _19702_);
  and _51997_ (_19704_, _06615_, _23707_);
  and _51998_ (_19705_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or _51999_ (_11738_, _19705_, _19704_);
  or _52000_ (_19706_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and _52001_ (_11754_, _19706_, _05482_);
  and _52002_ (_19707_, _15004_, _23898_);
  and _52003_ (_19708_, _15006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or _52004_ (_11755_, _19708_, _19707_);
  nor _52005_ (_11758_, _00759_, rst);
  and _52006_ (_11759_, _00341_, _22762_);
  and _52007_ (_11762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _22762_);
  and _52008_ (_19709_, _05119_, _23649_);
  and _52009_ (_19710_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  or _52010_ (_11783_, _19710_, _19709_);
  and _52011_ (_19711_, _25571_, _24050_);
  and _52012_ (_19712_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or _52013_ (_11787_, _19712_, _19711_);
  and _52014_ (_19713_, _02087_, _23946_);
  and _52015_ (_19714_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or _52016_ (_27009_, _19714_, _19713_);
  and _52017_ (_19715_, _17092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and _52018_ (_19716_, _17091_, _23778_);
  or _52019_ (_27241_, _19716_, _19715_);
  and _52020_ (_19717_, _04656_, _23946_);
  and _52021_ (_19718_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or _52022_ (_11791_, _19718_, _19717_);
  and _52023_ (_19719_, _04832_, _23898_);
  and _52024_ (_19720_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or _52025_ (_11793_, _19720_, _19719_);
  or _52026_ (_19721_, _05223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and _52027_ (_11795_, _19721_, _05224_);
  and _52028_ (_19722_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and _52029_ (_19723_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or _52030_ (_19724_, _19723_, _19722_);
  and _52031_ (_19725_, _19724_, _02393_);
  and _52032_ (_19726_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and _52033_ (_19727_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or _52034_ (_19728_, _19727_, _19726_);
  and _52035_ (_19729_, _19728_, _02445_);
  or _52036_ (_19730_, _19729_, _19725_);
  and _52037_ (_19731_, _19730_, _02421_);
  and _52038_ (_19732_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and _52039_ (_19733_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or _52040_ (_19734_, _19733_, _19732_);
  and _52041_ (_19735_, _19734_, _02393_);
  and _52042_ (_19736_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and _52043_ (_19737_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or _52044_ (_19738_, _19737_, _19736_);
  and _52045_ (_19739_, _19738_, _02445_);
  or _52046_ (_19740_, _19739_, _19735_);
  and _52047_ (_19741_, _19740_, _02459_);
  or _52048_ (_19742_, _19741_, _19731_);
  and _52049_ (_19743_, _19742_, _02458_);
  or _52050_ (_19744_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or _52051_ (_19745_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and _52052_ (_19746_, _19745_, _19744_);
  and _52053_ (_19747_, _19746_, _02393_);
  or _52054_ (_19748_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or _52055_ (_19749_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and _52056_ (_19750_, _19749_, _19748_);
  and _52057_ (_19751_, _19750_, _02445_);
  or _52058_ (_19752_, _19751_, _19747_);
  and _52059_ (_19753_, _19752_, _02421_);
  or _52060_ (_19754_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or _52061_ (_19755_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and _52062_ (_19756_, _19755_, _19754_);
  and _52063_ (_19757_, _19756_, _02393_);
  or _52064_ (_19758_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or _52065_ (_19759_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and _52066_ (_19760_, _19759_, _19758_);
  and _52067_ (_19761_, _19760_, _02445_);
  or _52068_ (_19762_, _19761_, _19757_);
  and _52069_ (_19763_, _19762_, _02459_);
  or _52070_ (_19764_, _19763_, _19753_);
  and _52071_ (_19765_, _19764_, _02414_);
  or _52072_ (_19766_, _19765_, _19743_);
  and _52073_ (_19767_, _19766_, _02398_);
  and _52074_ (_19768_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and _52075_ (_19769_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or _52076_ (_19770_, _19769_, _19768_);
  and _52077_ (_19771_, _19770_, _02393_);
  and _52078_ (_19772_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and _52079_ (_19773_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or _52080_ (_19774_, _19773_, _19772_);
  and _52081_ (_19775_, _19774_, _02445_);
  or _52082_ (_19776_, _19775_, _19771_);
  and _52083_ (_19777_, _19776_, _02421_);
  and _52084_ (_19778_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and _52085_ (_19779_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or _52086_ (_19780_, _19779_, _19778_);
  and _52087_ (_19781_, _19780_, _02393_);
  and _52088_ (_19782_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and _52089_ (_19783_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or _52090_ (_19784_, _19783_, _19782_);
  and _52091_ (_19785_, _19784_, _02445_);
  or _52092_ (_19786_, _19785_, _19781_);
  and _52093_ (_19787_, _19786_, _02459_);
  or _52094_ (_19788_, _19787_, _19777_);
  and _52095_ (_19789_, _19788_, _02458_);
  or _52096_ (_19790_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or _52097_ (_19791_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and _52098_ (_19792_, _19791_, _02445_);
  and _52099_ (_19793_, _19792_, _19790_);
  or _52100_ (_19794_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or _52101_ (_19795_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and _52102_ (_19796_, _19795_, _02393_);
  and _52103_ (_19797_, _19796_, _19794_);
  or _52104_ (_19798_, _19797_, _19793_);
  and _52105_ (_19799_, _19798_, _02421_);
  or _52106_ (_19800_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or _52107_ (_19801_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and _52108_ (_19802_, _19801_, _02445_);
  and _52109_ (_19803_, _19802_, _19800_);
  or _52110_ (_19804_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or _52111_ (_19805_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and _52112_ (_19806_, _19805_, _02393_);
  and _52113_ (_19807_, _19806_, _19804_);
  or _52114_ (_19808_, _19807_, _19803_);
  and _52115_ (_19809_, _19808_, _02459_);
  or _52116_ (_19810_, _19809_, _19799_);
  and _52117_ (_19811_, _19810_, _02414_);
  or _52118_ (_19812_, _19811_, _19789_);
  and _52119_ (_19813_, _19812_, _02496_);
  or _52120_ (_19814_, _19813_, _19767_);
  and _52121_ (_19815_, _19814_, _02400_);
  and _52122_ (_19816_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and _52123_ (_19817_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or _52124_ (_19818_, _19817_, _19816_);
  and _52125_ (_19819_, _19818_, _02393_);
  and _52126_ (_19820_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and _52127_ (_19821_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or _52128_ (_19822_, _19821_, _19820_);
  and _52129_ (_19823_, _19822_, _02445_);
  or _52130_ (_19824_, _19823_, _19819_);
  or _52131_ (_19825_, _19824_, _02459_);
  and _52132_ (_19826_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and _52133_ (_19827_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or _52134_ (_19828_, _19827_, _19826_);
  and _52135_ (_19829_, _19828_, _02393_);
  and _52136_ (_19830_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and _52137_ (_19831_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or _52138_ (_19832_, _19831_, _19830_);
  and _52139_ (_19833_, _19832_, _02445_);
  or _52140_ (_19834_, _19833_, _19829_);
  or _52141_ (_19835_, _19834_, _02421_);
  and _52142_ (_19836_, _19835_, _02458_);
  and _52143_ (_19837_, _19836_, _19825_);
  or _52144_ (_19838_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or _52145_ (_19839_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and _52146_ (_19840_, _19839_, _02445_);
  and _52147_ (_19841_, _19840_, _19838_);
  or _52148_ (_19842_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or _52149_ (_19843_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and _52150_ (_19844_, _19843_, _02393_);
  and _52151_ (_19845_, _19844_, _19842_);
  or _52152_ (_19846_, _19845_, _19841_);
  or _52153_ (_19847_, _19846_, _02459_);
  or _52154_ (_19848_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or _52155_ (_19849_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and _52156_ (_19850_, _19849_, _02445_);
  and _52157_ (_19851_, _19850_, _19848_);
  or _52158_ (_19852_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or _52159_ (_19853_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and _52160_ (_19854_, _19853_, _02393_);
  and _52161_ (_19855_, _19854_, _19852_);
  or _52162_ (_19856_, _19855_, _19851_);
  or _52163_ (_19857_, _19856_, _02421_);
  and _52164_ (_19858_, _19857_, _02414_);
  and _52165_ (_19859_, _19858_, _19847_);
  or _52166_ (_19860_, _19859_, _19837_);
  and _52167_ (_19861_, _19860_, _02496_);
  and _52168_ (_19862_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and _52169_ (_19863_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or _52170_ (_19864_, _19863_, _19862_);
  and _52171_ (_19865_, _19864_, _02393_);
  and _52172_ (_19866_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and _52173_ (_19867_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or _52174_ (_19868_, _19867_, _19866_);
  and _52175_ (_19869_, _19868_, _02445_);
  or _52176_ (_19870_, _19869_, _19865_);
  or _52177_ (_19871_, _19870_, _02459_);
  and _52178_ (_19872_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and _52179_ (_19873_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or _52180_ (_19874_, _19873_, _19872_);
  and _52181_ (_19875_, _19874_, _02393_);
  and _52182_ (_19876_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and _52183_ (_19877_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or _52184_ (_19878_, _19877_, _19876_);
  and _52185_ (_19879_, _19878_, _02445_);
  or _52186_ (_19880_, _19879_, _19875_);
  or _52187_ (_19881_, _19880_, _02421_);
  and _52188_ (_19882_, _19881_, _02458_);
  and _52189_ (_19883_, _19882_, _19871_);
  or _52190_ (_19884_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or _52191_ (_19885_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and _52192_ (_19886_, _19885_, _19884_);
  and _52193_ (_19887_, _19886_, _02393_);
  or _52194_ (_19888_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or _52195_ (_19889_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and _52196_ (_19890_, _19889_, _19888_);
  and _52197_ (_19891_, _19890_, _02445_);
  or _52198_ (_19892_, _19891_, _19887_);
  or _52199_ (_19893_, _19892_, _02459_);
  or _52200_ (_19894_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or _52201_ (_19895_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and _52202_ (_19896_, _19895_, _19894_);
  and _52203_ (_19897_, _19896_, _02393_);
  or _52204_ (_19898_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or _52205_ (_19899_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and _52206_ (_19900_, _19899_, _19898_);
  and _52207_ (_19901_, _19900_, _02445_);
  or _52208_ (_19902_, _19901_, _19897_);
  or _52209_ (_19903_, _19902_, _02421_);
  and _52210_ (_19904_, _19903_, _02414_);
  and _52211_ (_19905_, _19904_, _19893_);
  or _52212_ (_19906_, _19905_, _19883_);
  and _52213_ (_19907_, _19906_, _02398_);
  or _52214_ (_19908_, _19907_, _19861_);
  and _52215_ (_19909_, _19908_, _02546_);
  or _52216_ (_19910_, _19909_, _19815_);
  and _52217_ (_19911_, _19910_, _02646_);
  or _52218_ (_19912_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or _52219_ (_19913_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and _52220_ (_19914_, _19913_, _02445_);
  and _52221_ (_19915_, _19914_, _19912_);
  or _52222_ (_19916_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or _52223_ (_19917_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and _52224_ (_19918_, _19917_, _02393_);
  and _52225_ (_19919_, _19918_, _19916_);
  or _52226_ (_19921_, _19919_, _19915_);
  and _52227_ (_19922_, _19921_, _02459_);
  or _52228_ (_19923_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or _52229_ (_19924_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and _52230_ (_19925_, _19924_, _02445_);
  and _52231_ (_19926_, _19925_, _19923_);
  or _52232_ (_19927_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or _52233_ (_19928_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and _52234_ (_19929_, _19928_, _02393_);
  and _52235_ (_19930_, _19929_, _19927_);
  or _52236_ (_19931_, _19930_, _19926_);
  and _52237_ (_19932_, _19931_, _02421_);
  or _52238_ (_19933_, _19932_, _19922_);
  and _52239_ (_19934_, _19933_, _02414_);
  and _52240_ (_19935_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and _52241_ (_19936_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or _52242_ (_19937_, _19936_, _19935_);
  and _52243_ (_19938_, _19937_, _02393_);
  and _52244_ (_19939_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and _52245_ (_19940_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or _52246_ (_19942_, _19940_, _19939_);
  and _52247_ (_19943_, _19942_, _02445_);
  or _52248_ (_19944_, _19943_, _19938_);
  and _52249_ (_19945_, _19944_, _02459_);
  and _52250_ (_19946_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and _52251_ (_19947_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or _52252_ (_19948_, _19947_, _19946_);
  and _52253_ (_19949_, _19948_, _02393_);
  and _52254_ (_19950_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and _52255_ (_19951_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or _52256_ (_19952_, _19951_, _19950_);
  and _52257_ (_19953_, _19952_, _02445_);
  or _52258_ (_19954_, _19953_, _19949_);
  and _52259_ (_19955_, _19954_, _02421_);
  or _52260_ (_19956_, _19955_, _19945_);
  and _52261_ (_19957_, _19956_, _02458_);
  or _52262_ (_19958_, _19957_, _19934_);
  and _52263_ (_19959_, _19958_, _02496_);
  or _52264_ (_19960_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or _52265_ (_19961_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and _52266_ (_19962_, _19961_, _19960_);
  and _52267_ (_19963_, _19962_, _02393_);
  or _52268_ (_19964_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or _52269_ (_19965_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and _52270_ (_19966_, _19965_, _19964_);
  and _52271_ (_19967_, _19966_, _02445_);
  or _52272_ (_19968_, _19967_, _19963_);
  and _52273_ (_19969_, _19968_, _02459_);
  or _52274_ (_19970_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or _52275_ (_19971_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and _52276_ (_19973_, _19971_, _19970_);
  and _52277_ (_19974_, _19973_, _02393_);
  or _52278_ (_19975_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or _52279_ (_19976_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and _52280_ (_19977_, _19976_, _19975_);
  and _52281_ (_19978_, _19977_, _02445_);
  or _52282_ (_19979_, _19978_, _19974_);
  and _52283_ (_19980_, _19979_, _02421_);
  or _52284_ (_19981_, _19980_, _19969_);
  and _52285_ (_19982_, _19981_, _02414_);
  and _52286_ (_19983_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and _52287_ (_19984_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or _52288_ (_19985_, _19984_, _19983_);
  and _52289_ (_19986_, _19985_, _02393_);
  and _52290_ (_19987_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and _52291_ (_19988_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or _52292_ (_19989_, _19988_, _19987_);
  and _52293_ (_19990_, _19989_, _02445_);
  or _52294_ (_19991_, _19990_, _19986_);
  and _52295_ (_19992_, _19991_, _02459_);
  and _52296_ (_19993_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and _52297_ (_19994_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or _52298_ (_19995_, _19994_, _19993_);
  and _52299_ (_19996_, _19995_, _02393_);
  and _52300_ (_19997_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and _52301_ (_19998_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or _52302_ (_19999_, _19998_, _19997_);
  and _52303_ (_20000_, _19999_, _02445_);
  or _52304_ (_20001_, _20000_, _19996_);
  and _52305_ (_20002_, _20001_, _02421_);
  or _52306_ (_20003_, _20002_, _19992_);
  and _52307_ (_20004_, _20003_, _02458_);
  or _52308_ (_20005_, _20004_, _19982_);
  and _52309_ (_20006_, _20005_, _02398_);
  or _52310_ (_20007_, _20006_, _19959_);
  and _52311_ (_20008_, _20007_, _02400_);
  and _52312_ (_20009_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and _52313_ (_20010_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or _52314_ (_20011_, _20010_, _20009_);
  and _52315_ (_20012_, _20011_, _02393_);
  and _52316_ (_20013_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and _52317_ (_20014_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or _52318_ (_20015_, _20014_, _20013_);
  and _52319_ (_20016_, _20015_, _02445_);
  or _52320_ (_20017_, _20016_, _20012_);
  or _52321_ (_20018_, _20017_, _02459_);
  and _52322_ (_20019_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and _52323_ (_20020_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or _52324_ (_20021_, _20020_, _20019_);
  and _52325_ (_20022_, _20021_, _02393_);
  and _52326_ (_20023_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and _52327_ (_20024_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or _52328_ (_20025_, _20024_, _20023_);
  and _52329_ (_20026_, _20025_, _02445_);
  or _52330_ (_20027_, _20026_, _20022_);
  or _52331_ (_20028_, _20027_, _02421_);
  and _52332_ (_20029_, _20028_, _02458_);
  and _52333_ (_20030_, _20029_, _20018_);
  or _52334_ (_20031_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or _52335_ (_20032_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and _52336_ (_20033_, _20032_, _20031_);
  and _52337_ (_20034_, _20033_, _02393_);
  or _52338_ (_20035_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or _52339_ (_20036_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and _52340_ (_20037_, _20036_, _20035_);
  and _52341_ (_20038_, _20037_, _02445_);
  or _52342_ (_20039_, _20038_, _20034_);
  or _52343_ (_20040_, _20039_, _02459_);
  or _52344_ (_20041_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or _52345_ (_20042_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and _52346_ (_20044_, _20042_, _20041_);
  and _52347_ (_20045_, _20044_, _02393_);
  or _52348_ (_20046_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or _52349_ (_20047_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and _52350_ (_20048_, _20047_, _20046_);
  and _52351_ (_20049_, _20048_, _02445_);
  or _52352_ (_20050_, _20049_, _20045_);
  or _52353_ (_20051_, _20050_, _02421_);
  and _52354_ (_20052_, _20051_, _02414_);
  and _52355_ (_20053_, _20052_, _20040_);
  or _52356_ (_20054_, _20053_, _20030_);
  and _52357_ (_20055_, _20054_, _02398_);
  and _52358_ (_20056_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and _52359_ (_20057_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or _52360_ (_20058_, _20057_, _20056_);
  and _52361_ (_20059_, _20058_, _02393_);
  and _52362_ (_20060_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and _52363_ (_20061_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or _52364_ (_20062_, _20061_, _20060_);
  and _52365_ (_20063_, _20062_, _02445_);
  or _52366_ (_20064_, _20063_, _20059_);
  or _52367_ (_20065_, _20064_, _02459_);
  and _52368_ (_20066_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and _52369_ (_20067_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or _52370_ (_20068_, _20067_, _20066_);
  and _52371_ (_20069_, _20068_, _02393_);
  and _52372_ (_20070_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and _52373_ (_20071_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or _52374_ (_20072_, _20071_, _20070_);
  and _52375_ (_20073_, _20072_, _02445_);
  or _52376_ (_20074_, _20073_, _20069_);
  or _52377_ (_20075_, _20074_, _02421_);
  and _52378_ (_20076_, _20075_, _02458_);
  and _52379_ (_20077_, _20076_, _20065_);
  or _52380_ (_20078_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or _52381_ (_20079_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and _52382_ (_20080_, _20079_, _02445_);
  and _52383_ (_20081_, _20080_, _20078_);
  or _52384_ (_20082_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or _52385_ (_20083_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and _52386_ (_20084_, _20083_, _02393_);
  and _52387_ (_20085_, _20084_, _20082_);
  or _52388_ (_20086_, _20085_, _20081_);
  or _52389_ (_20087_, _20086_, _02459_);
  or _52390_ (_20088_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or _52391_ (_20089_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and _52392_ (_20090_, _20089_, _02445_);
  and _52393_ (_20091_, _20090_, _20088_);
  or _52394_ (_20092_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or _52395_ (_20093_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and _52396_ (_20094_, _20093_, _02393_);
  and _52397_ (_20095_, _20094_, _20092_);
  or _52398_ (_20096_, _20095_, _20091_);
  or _52399_ (_20097_, _20096_, _02421_);
  and _52400_ (_20098_, _20097_, _02414_);
  and _52401_ (_20099_, _20098_, _20087_);
  or _52402_ (_20100_, _20099_, _20077_);
  and _52403_ (_20101_, _20100_, _02496_);
  or _52404_ (_20102_, _20101_, _20055_);
  and _52405_ (_20103_, _20102_, _02546_);
  or _52406_ (_20104_, _20103_, _20008_);
  and _52407_ (_20105_, _20104_, _02405_);
  or _52408_ (_20106_, _20105_, _19911_);
  and _52409_ (_20107_, _20106_, _26777_);
  and _52410_ (_20108_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and _52411_ (_20109_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or _52412_ (_20110_, _20109_, _20108_);
  and _52413_ (_20111_, _20110_, _02393_);
  and _52414_ (_20112_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  and _52415_ (_20113_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or _52416_ (_20114_, _20113_, _20112_);
  and _52417_ (_20115_, _20114_, _02445_);
  or _52418_ (_20116_, _20115_, _20111_);
  and _52419_ (_20117_, _20116_, _02421_);
  and _52420_ (_20118_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and _52421_ (_20119_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or _52422_ (_20120_, _20119_, _20118_);
  and _52423_ (_20121_, _20120_, _02393_);
  and _52424_ (_20122_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and _52425_ (_20123_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or _52426_ (_20124_, _20123_, _20122_);
  and _52427_ (_20125_, _20124_, _02445_);
  or _52428_ (_20126_, _20125_, _20121_);
  and _52429_ (_20127_, _20126_, _02459_);
  or _52430_ (_20128_, _20127_, _20117_);
  and _52431_ (_20129_, _20128_, _02458_);
  or _52432_ (_20130_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or _52433_ (_20131_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and _52434_ (_20132_, _20131_, _20130_);
  and _52435_ (_20133_, _20132_, _02393_);
  or _52436_ (_20134_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or _52437_ (_20135_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and _52438_ (_20136_, _20135_, _20134_);
  and _52439_ (_20137_, _20136_, _02445_);
  or _52440_ (_20138_, _20137_, _20133_);
  and _52441_ (_20139_, _20138_, _02421_);
  or _52442_ (_20140_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or _52443_ (_20141_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and _52444_ (_20142_, _20141_, _20140_);
  and _52445_ (_20143_, _20142_, _02393_);
  or _52446_ (_20144_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or _52447_ (_20145_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and _52448_ (_20146_, _20145_, _20144_);
  and _52449_ (_20147_, _20146_, _02445_);
  or _52450_ (_20148_, _20147_, _20143_);
  and _52451_ (_20149_, _20148_, _02459_);
  or _52452_ (_20150_, _20149_, _20139_);
  and _52453_ (_20151_, _20150_, _02414_);
  or _52454_ (_20152_, _20151_, _20129_);
  and _52455_ (_20153_, _20152_, _02398_);
  and _52456_ (_20154_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and _52457_ (_20155_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or _52458_ (_20156_, _20155_, _20154_);
  and _52459_ (_20157_, _20156_, _02393_);
  and _52460_ (_20158_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and _52461_ (_20159_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or _52462_ (_20160_, _20159_, _20158_);
  and _52463_ (_20161_, _20160_, _02445_);
  or _52464_ (_20162_, _20161_, _20157_);
  and _52465_ (_20163_, _20162_, _02421_);
  and _52466_ (_20164_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and _52467_ (_20165_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _52468_ (_20166_, _20165_, _20164_);
  and _52469_ (_20167_, _20166_, _02393_);
  and _52470_ (_20168_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and _52471_ (_20169_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or _52472_ (_20170_, _20169_, _20168_);
  and _52473_ (_20171_, _20170_, _02445_);
  or _52474_ (_20172_, _20171_, _20167_);
  and _52475_ (_20173_, _20172_, _02459_);
  or _52476_ (_20174_, _20173_, _20163_);
  and _52477_ (_20175_, _20174_, _02458_);
  or _52478_ (_20176_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or _52479_ (_20177_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and _52480_ (_20178_, _20177_, _02445_);
  and _52481_ (_20179_, _20178_, _20176_);
  or _52482_ (_20180_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or _52483_ (_20181_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and _52484_ (_20182_, _20181_, _02393_);
  and _52485_ (_20183_, _20182_, _20180_);
  or _52486_ (_20184_, _20183_, _20179_);
  and _52487_ (_20185_, _20184_, _02421_);
  or _52488_ (_20186_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or _52489_ (_20187_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and _52490_ (_20188_, _20187_, _02445_);
  and _52491_ (_20189_, _20188_, _20186_);
  or _52492_ (_20190_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or _52493_ (_20191_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and _52494_ (_20192_, _20191_, _02393_);
  and _52495_ (_20193_, _20192_, _20190_);
  or _52496_ (_20194_, _20193_, _20189_);
  and _52497_ (_20195_, _20194_, _02459_);
  or _52498_ (_20196_, _20195_, _20185_);
  and _52499_ (_20197_, _20196_, _02414_);
  or _52500_ (_20198_, _20197_, _20175_);
  and _52501_ (_20199_, _20198_, _02496_);
  or _52502_ (_20200_, _20199_, _20153_);
  and _52503_ (_20201_, _20200_, _02400_);
  and _52504_ (_20202_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and _52505_ (_20203_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or _52506_ (_20204_, _20203_, _20202_);
  and _52507_ (_20205_, _20204_, _02393_);
  and _52508_ (_20206_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and _52509_ (_20207_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or _52510_ (_20208_, _20207_, _20206_);
  and _52511_ (_20209_, _20208_, _02445_);
  or _52512_ (_20210_, _20209_, _20205_);
  or _52513_ (_20211_, _20210_, _02459_);
  and _52514_ (_20212_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and _52515_ (_20213_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or _52516_ (_20214_, _20213_, _20212_);
  and _52517_ (_20215_, _20214_, _02393_);
  and _52518_ (_20216_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and _52519_ (_20217_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or _52520_ (_20218_, _20217_, _20216_);
  and _52521_ (_20219_, _20218_, _02445_);
  or _52522_ (_20220_, _20219_, _20215_);
  or _52523_ (_20221_, _20220_, _02421_);
  and _52524_ (_20222_, _20221_, _02458_);
  and _52525_ (_20223_, _20222_, _20211_);
  or _52526_ (_20224_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or _52527_ (_20225_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  and _52528_ (_20226_, _20225_, _02445_);
  and _52529_ (_20227_, _20226_, _20224_);
  or _52530_ (_20228_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or _52531_ (_20229_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  and _52532_ (_20230_, _20229_, _02393_);
  and _52533_ (_20231_, _20230_, _20228_);
  or _52534_ (_20232_, _20231_, _20227_);
  or _52535_ (_20233_, _20232_, _02459_);
  or _52536_ (_20234_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or _52537_ (_20235_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and _52538_ (_20236_, _20235_, _02445_);
  and _52539_ (_20237_, _20236_, _20234_);
  or _52540_ (_20238_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or _52541_ (_20239_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and _52542_ (_20240_, _20239_, _02393_);
  and _52543_ (_20241_, _20240_, _20238_);
  or _52544_ (_20242_, _20241_, _20237_);
  or _52545_ (_20243_, _20242_, _02421_);
  and _52546_ (_20244_, _20243_, _02414_);
  and _52547_ (_20245_, _20244_, _20233_);
  or _52548_ (_20246_, _20245_, _20223_);
  and _52549_ (_20247_, _20246_, _02496_);
  and _52550_ (_20248_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and _52551_ (_20249_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or _52552_ (_20250_, _20249_, _20248_);
  and _52553_ (_20251_, _20250_, _02393_);
  and _52554_ (_20252_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and _52555_ (_20253_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or _52556_ (_20254_, _20253_, _20252_);
  and _52557_ (_20255_, _20254_, _02445_);
  or _52558_ (_20256_, _20255_, _20251_);
  or _52559_ (_20257_, _20256_, _02459_);
  and _52560_ (_20258_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and _52561_ (_20259_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or _52562_ (_20260_, _20259_, _20258_);
  and _52563_ (_20261_, _20260_, _02393_);
  and _52564_ (_20262_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and _52565_ (_20263_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or _52566_ (_20264_, _20263_, _20262_);
  and _52567_ (_20265_, _20264_, _02445_);
  or _52568_ (_20266_, _20265_, _20261_);
  or _52569_ (_20267_, _20266_, _02421_);
  and _52570_ (_20268_, _20267_, _02458_);
  and _52571_ (_20269_, _20268_, _20257_);
  or _52572_ (_20270_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or _52573_ (_20271_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and _52574_ (_20272_, _20271_, _20270_);
  and _52575_ (_20273_, _20272_, _02393_);
  or _52576_ (_20274_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or _52577_ (_20275_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and _52578_ (_20276_, _20275_, _20274_);
  and _52579_ (_20277_, _20276_, _02445_);
  or _52580_ (_20278_, _20277_, _20273_);
  or _52581_ (_20279_, _20278_, _02459_);
  or _52582_ (_20280_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or _52583_ (_20281_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and _52584_ (_20282_, _20281_, _20280_);
  and _52585_ (_20283_, _20282_, _02393_);
  or _52586_ (_20284_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or _52587_ (_20285_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and _52588_ (_20286_, _20285_, _20284_);
  and _52589_ (_20287_, _20286_, _02445_);
  or _52590_ (_20288_, _20287_, _20283_);
  or _52591_ (_20289_, _20288_, _02421_);
  and _52592_ (_20290_, _20289_, _02414_);
  and _52593_ (_20291_, _20290_, _20279_);
  or _52594_ (_20292_, _20291_, _20269_);
  and _52595_ (_20293_, _20292_, _02398_);
  or _52596_ (_20294_, _20293_, _20247_);
  and _52597_ (_20295_, _20294_, _02546_);
  or _52598_ (_20296_, _20295_, _20201_);
  and _52599_ (_20297_, _20296_, _02646_);
  or _52600_ (_20298_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or _52601_ (_20299_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  and _52602_ (_20300_, _20299_, _02445_);
  and _52603_ (_20301_, _20300_, _20298_);
  or _52604_ (_20302_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or _52605_ (_20303_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and _52606_ (_20304_, _20303_, _02393_);
  and _52607_ (_20305_, _20304_, _20302_);
  or _52608_ (_20306_, _20305_, _20301_);
  and _52609_ (_20307_, _20306_, _02459_);
  or _52610_ (_20308_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or _52611_ (_20309_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  and _52612_ (_20310_, _20309_, _02445_);
  and _52613_ (_20311_, _20310_, _20308_);
  or _52614_ (_20312_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or _52615_ (_20313_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and _52616_ (_20314_, _20313_, _02393_);
  and _52617_ (_20315_, _20314_, _20312_);
  or _52618_ (_20316_, _20315_, _20311_);
  and _52619_ (_20317_, _20316_, _02421_);
  or _52620_ (_20318_, _20317_, _20307_);
  and _52621_ (_20319_, _20318_, _02414_);
  and _52622_ (_20320_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and _52623_ (_20321_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or _52624_ (_20322_, _20321_, _20320_);
  and _52625_ (_20323_, _20322_, _02393_);
  and _52626_ (_20324_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  and _52627_ (_20325_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or _52628_ (_20326_, _20325_, _20324_);
  and _52629_ (_20327_, _20326_, _02445_);
  or _52630_ (_20328_, _20327_, _20323_);
  and _52631_ (_20329_, _20328_, _02459_);
  and _52632_ (_20330_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  and _52633_ (_20331_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or _52634_ (_20332_, _20331_, _20330_);
  and _52635_ (_20333_, _20332_, _02393_);
  and _52636_ (_20334_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and _52637_ (_20335_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or _52638_ (_20336_, _20335_, _20334_);
  and _52639_ (_20337_, _20336_, _02445_);
  or _52640_ (_20338_, _20337_, _20333_);
  and _52641_ (_20339_, _20338_, _02421_);
  or _52642_ (_20340_, _20339_, _20329_);
  and _52643_ (_20341_, _20340_, _02458_);
  or _52644_ (_20342_, _20341_, _20319_);
  and _52645_ (_20343_, _20342_, _02496_);
  or _52646_ (_20344_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or _52647_ (_20345_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and _52648_ (_20346_, _20345_, _20344_);
  and _52649_ (_20347_, _20346_, _02393_);
  or _52650_ (_20348_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or _52651_ (_20349_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  and _52652_ (_20350_, _20349_, _20348_);
  and _52653_ (_20351_, _20350_, _02445_);
  or _52654_ (_20352_, _20351_, _20347_);
  and _52655_ (_20353_, _20352_, _02459_);
  or _52656_ (_20354_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or _52657_ (_20355_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and _52658_ (_20356_, _20355_, _20354_);
  and _52659_ (_20357_, _20356_, _02393_);
  or _52660_ (_20358_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or _52661_ (_20359_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and _52662_ (_20360_, _20359_, _20358_);
  and _52663_ (_20361_, _20360_, _02445_);
  or _52664_ (_20362_, _20361_, _20357_);
  and _52665_ (_20363_, _20362_, _02421_);
  or _52666_ (_20364_, _20363_, _20353_);
  and _52667_ (_20365_, _20364_, _02414_);
  and _52668_ (_20366_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and _52669_ (_20367_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or _52670_ (_20368_, _20367_, _20366_);
  and _52671_ (_20369_, _20368_, _02393_);
  and _52672_ (_20370_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and _52673_ (_20371_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or _52674_ (_20372_, _20371_, _20370_);
  and _52675_ (_20373_, _20372_, _02445_);
  or _52676_ (_20374_, _20373_, _20369_);
  and _52677_ (_20375_, _20374_, _02459_);
  and _52678_ (_20376_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and _52679_ (_20377_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or _52680_ (_20378_, _20377_, _20376_);
  and _52681_ (_20379_, _20378_, _02393_);
  and _52682_ (_20380_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and _52683_ (_20381_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or _52684_ (_20382_, _20381_, _20380_);
  and _52685_ (_20383_, _20382_, _02445_);
  or _52686_ (_20384_, _20383_, _20379_);
  and _52687_ (_20385_, _20384_, _02421_);
  or _52688_ (_20386_, _20385_, _20375_);
  and _52689_ (_20387_, _20386_, _02458_);
  or _52690_ (_20388_, _20387_, _20365_);
  and _52691_ (_20389_, _20388_, _02398_);
  or _52692_ (_20390_, _20389_, _20343_);
  and _52693_ (_20391_, _20390_, _02400_);
  and _52694_ (_20392_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and _52695_ (_20393_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or _52696_ (_20394_, _20393_, _20392_);
  and _52697_ (_20395_, _20394_, _02393_);
  and _52698_ (_20396_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and _52699_ (_20397_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or _52700_ (_20398_, _20397_, _20396_);
  and _52701_ (_20399_, _20398_, _02445_);
  or _52702_ (_20400_, _20399_, _20395_);
  or _52703_ (_20401_, _20400_, _02459_);
  and _52704_ (_20402_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and _52705_ (_20403_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or _52706_ (_20404_, _20403_, _20402_);
  and _52707_ (_20405_, _20404_, _02393_);
  and _52708_ (_20406_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and _52709_ (_20407_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or _52710_ (_20408_, _20407_, _20406_);
  and _52711_ (_20409_, _20408_, _02445_);
  or _52712_ (_20410_, _20409_, _20405_);
  or _52713_ (_20411_, _20410_, _02421_);
  and _52714_ (_20412_, _20411_, _02458_);
  and _52715_ (_20413_, _20412_, _20401_);
  or _52716_ (_20414_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or _52717_ (_20415_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and _52718_ (_20416_, _20415_, _20414_);
  and _52719_ (_20417_, _20416_, _02393_);
  or _52720_ (_20418_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or _52721_ (_20419_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and _52722_ (_20420_, _20419_, _20418_);
  and _52723_ (_20421_, _20420_, _02445_);
  or _52724_ (_20422_, _20421_, _20417_);
  or _52725_ (_20423_, _20422_, _02459_);
  or _52726_ (_20424_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or _52727_ (_20425_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and _52728_ (_20426_, _20425_, _20424_);
  and _52729_ (_20427_, _20426_, _02393_);
  or _52730_ (_20428_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or _52731_ (_20429_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and _52732_ (_20430_, _20429_, _20428_);
  and _52733_ (_20431_, _20430_, _02445_);
  or _52734_ (_20432_, _20431_, _20427_);
  or _52735_ (_20433_, _20432_, _02421_);
  and _52736_ (_20434_, _20433_, _02414_);
  and _52737_ (_20435_, _20434_, _20423_);
  or _52738_ (_20436_, _20435_, _20413_);
  and _52739_ (_20437_, _20436_, _02398_);
  and _52740_ (_20438_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and _52741_ (_20439_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or _52742_ (_20440_, _20439_, _20438_);
  and _52743_ (_20441_, _20440_, _02393_);
  and _52744_ (_20442_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and _52745_ (_20443_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or _52746_ (_20444_, _20443_, _20442_);
  and _52747_ (_20445_, _20444_, _02445_);
  or _52748_ (_20446_, _20445_, _20441_);
  or _52749_ (_20447_, _20446_, _02459_);
  and _52750_ (_20448_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and _52751_ (_20449_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or _52752_ (_20450_, _20449_, _20448_);
  and _52753_ (_20451_, _20450_, _02393_);
  and _52754_ (_20452_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and _52755_ (_20453_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or _52756_ (_20454_, _20453_, _20452_);
  and _52757_ (_20455_, _20454_, _02445_);
  or _52758_ (_20456_, _20455_, _20451_);
  or _52759_ (_20457_, _20456_, _02421_);
  and _52760_ (_20458_, _20457_, _02458_);
  and _52761_ (_20459_, _20458_, _20447_);
  or _52762_ (_20460_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or _52763_ (_20461_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and _52764_ (_20462_, _20461_, _02445_);
  and _52765_ (_20463_, _20462_, _20460_);
  or _52766_ (_20464_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or _52767_ (_20465_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and _52768_ (_20466_, _20465_, _02393_);
  and _52769_ (_20467_, _20466_, _20464_);
  or _52770_ (_20468_, _20467_, _20463_);
  or _52771_ (_20469_, _20468_, _02459_);
  or _52772_ (_20470_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or _52773_ (_20471_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and _52774_ (_20472_, _20471_, _02445_);
  and _52775_ (_20473_, _20472_, _20470_);
  or _52776_ (_20474_, _02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or _52777_ (_20475_, _02429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  and _52778_ (_20476_, _20475_, _02393_);
  and _52779_ (_20477_, _20476_, _20474_);
  or _52780_ (_20478_, _20477_, _20473_);
  or _52781_ (_20479_, _20478_, _02421_);
  and _52782_ (_20480_, _20479_, _02414_);
  and _52783_ (_20481_, _20480_, _20469_);
  or _52784_ (_20482_, _20481_, _20459_);
  and _52785_ (_20483_, _20482_, _02496_);
  or _52786_ (_20484_, _20483_, _20437_);
  and _52787_ (_20485_, _20484_, _02546_);
  or _52788_ (_20486_, _20485_, _20391_);
  and _52789_ (_20487_, _20486_, _02405_);
  or _52790_ (_20488_, _20487_, _20297_);
  and _52791_ (_20489_, _20488_, _02444_);
  or _52792_ (_20490_, _20489_, _20107_);
  or _52793_ (_20491_, _20490_, _02443_);
  or _52794_ (_20492_, _03267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and _52795_ (_20493_, _20492_, _22762_);
  and _52796_ (_11797_, _20493_, _20491_);
  and _52797_ (_20494_, _06615_, _23824_);
  and _52798_ (_20495_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or _52799_ (_11803_, _20495_, _20494_);
  and _52800_ (_11817_, _00520_, _22762_);
  and _52801_ (_11828_, _03305_, _24862_);
  and _52802_ (_11830_, _00422_, _22762_);
  and _52803_ (_20496_, _06651_, _23707_);
  and _52804_ (_20497_, _06653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  or _52805_ (_11834_, _20497_, _20496_);
  and _52806_ (_20498_, _05346_, _23946_);
  and _52807_ (_20499_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or _52808_ (_11849_, _20499_, _20498_);
  and _52809_ (_20500_, _02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  and _52810_ (_20501_, _02306_, _23707_);
  or _52811_ (_11853_, _20501_, _20500_);
  and _52812_ (_20502_, _16376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and _52813_ (_20503_, _16375_, _23649_);
  or _52814_ (_11855_, _20503_, _20502_);
  and _52815_ (_11857_, _00673_, _22762_);
  and _52816_ (_11859_, _26370_, _22762_);
  and _52817_ (_20504_, _06552_, _23778_);
  and _52818_ (_20505_, _06554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or _52819_ (_11863_, _20505_, _20504_);
  and _52820_ (_20506_, _02087_, _24050_);
  and _52821_ (_20507_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or _52822_ (_11867_, _20507_, _20506_);
  or _52823_ (_20508_, _22770_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nand _52824_ (_20509_, _22770_, _14710_);
  and _52825_ (_20510_, _20509_, _22762_);
  and _52826_ (_26883_[15], _20510_, _20508_);
  and _52827_ (_11872_, _00595_, _22762_);
  and _52828_ (_20511_, _18217_, _23824_);
  and _52829_ (_20512_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or _52830_ (_11882_, _20512_, _20511_);
  and _52831_ (_20513_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and _52832_ (_20514_, _06507_, _23747_);
  or _52833_ (_11884_, _20514_, _20513_);
  and _52834_ (_20515_, _07743_, _24050_);
  and _52835_ (_20516_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  or _52836_ (_27073_, _20516_, _20515_);
  nand _52837_ (_20517_, _02077_, _23702_);
  and _52838_ (_20518_, _02076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _52839_ (_20519_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _52840_ (_20520_, _20519_, _20518_);
  or _52841_ (_20521_, _20520_, _02077_);
  and _52842_ (_20522_, _20521_, _12675_);
  and _52843_ (_20523_, _20522_, _20517_);
  and _52844_ (_20524_, _02073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _52845_ (_20525_, _20524_, _20523_);
  and _52846_ (_11891_, _20525_, _22762_);
  and _52847_ (_20526_, _07743_, _23707_);
  and _52848_ (_20527_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  or _52849_ (_27074_, _20527_, _20526_);
  and _52850_ (_20528_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and _52851_ (_20529_, _17255_, _23824_);
  or _52852_ (_11911_, _20529_, _20528_);
  and _52853_ (_20530_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and _52854_ (_20531_, _17255_, _23898_);
  or _52855_ (_11924_, _20531_, _20530_);
  and _52856_ (_20532_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and _52857_ (_20533_, _16325_, _24050_);
  or _52858_ (_11962_, _20533_, _20532_);
  and _52859_ (_20534_, _08642_, _23898_);
  and _52860_ (_20535_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  or _52861_ (_11964_, _20535_, _20534_);
  and _52862_ (_20536_, _03339_, _23707_);
  and _52863_ (_20537_, _03342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or _52864_ (_11998_, _20537_, _20536_);
  and _52865_ (_20538_, _08642_, _23824_);
  and _52866_ (_20539_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  or _52867_ (_12002_, _20539_, _20538_);
  and _52868_ (_20540_, _24086_, _23824_);
  and _52869_ (_20541_, _24088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or _52870_ (_12009_, _20541_, _20540_);
  and _52871_ (_20542_, _05459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or _52872_ (_26914_, _20542_, _05461_);
  and _52873_ (_20543_, _08642_, _23778_);
  and _52874_ (_20544_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  or _52875_ (_27141_, _20544_, _20543_);
  nor _52876_ (_20545_, _23596_, _26375_);
  and _52877_ (_20546_, _23596_, _26375_);
  or _52878_ (_20547_, _20546_, _20545_);
  and _52879_ (_12022_, _20547_, _22762_);
  or _52880_ (_20548_, _05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and _52881_ (_12024_, _20548_, _05470_);
  and _52882_ (_12026_, _01169_, _22762_);
  and _52883_ (_20549_, _06615_, _23898_);
  and _52884_ (_20550_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or _52885_ (_12028_, _20550_, _20549_);
  and _52886_ (_12035_, _00919_, _22762_);
  and _52887_ (_12037_, _00428_, _22762_);
  and _52888_ (_12040_, _01048_, _22762_);
  and _52889_ (_12042_, _01231_, _22762_);
  and _52890_ (_12044_, _00334_, _22762_);
  and _52891_ (_12048_, _01290_, _22762_);
  and _52892_ (_12050_, _26541_, _22762_);
  and _52893_ (_12052_, _01107_, _22762_);
  and _52894_ (_12054_, _04279_, _22762_);
  and _52895_ (_12056_, _00600_, _22762_);
  and _52896_ (_12060_, _00511_, _22762_);
  and _52897_ (_20551_, _05454_, _23747_);
  and _52898_ (_20552_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _52899_ (_12063_, _20552_, _20551_);
  and _52900_ (_20553_, _05454_, _23707_);
  and _52901_ (_20554_, _05457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _52902_ (_12066_, _20554_, _20553_);
  and _52903_ (_20555_, _05429_, _23707_);
  and _52904_ (_20556_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or _52905_ (_12068_, _20556_, _20555_);
  and _52906_ (_20557_, _05429_, _23946_);
  and _52907_ (_20558_, _05431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or _52908_ (_12070_, _20558_, _20557_);
  and _52909_ (_20559_, _05379_, _23649_);
  and _52910_ (_20560_, _05381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _52911_ (_12072_, _20560_, _20559_);
  and _52912_ (_12086_, _00679_, _22762_);
  and _52913_ (_20561_, _08642_, _23649_);
  and _52914_ (_20562_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  or _52915_ (_27142_, _20562_, _20561_);
  and _52916_ (_20563_, _17263_, _24050_);
  and _52917_ (_20564_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  or _52918_ (_12101_, _20564_, _20563_);
  and _52919_ (_20565_, _05200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  and _52920_ (_20566_, _05199_, _24050_);
  or _52921_ (_27232_, _20566_, _20565_);
  and _52922_ (_20567_, _05319_, _23824_);
  and _52923_ (_20568_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _52924_ (_12105_, _20568_, _20567_);
  and _52925_ (_20569_, _05346_, _23707_);
  and _52926_ (_20571_, _05348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or _52927_ (_12107_, _20571_, _20569_);
  and _52928_ (_20572_, _05319_, _24050_);
  and _52929_ (_20573_, _05322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or _52930_ (_12109_, _20573_, _20572_);
  and _52931_ (_20574_, _05298_, _23946_);
  and _52932_ (_20575_, _05301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or _52933_ (_12111_, _20575_, _20574_);
  and _52934_ (_20576_, _02107_, _23898_);
  and _52935_ (_20577_, _02109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  or _52936_ (_12113_, _20577_, _20576_);
  and _52937_ (_20578_, _05223_, _24050_);
  and _52938_ (_20579_, _05276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or _52939_ (_12116_, _20579_, _20578_);
  and _52940_ (_20580_, _07536_, _24050_);
  and _52941_ (_20581_, _07539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  or _52942_ (_27114_, _20581_, _20580_);
  and _52943_ (_20582_, _05119_, _23778_);
  and _52944_ (_20583_, _05121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  or _52945_ (_12185_, _20583_, _20582_);
  and _52946_ (_20584_, _05102_, _23649_);
  and _52947_ (_20585_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or _52948_ (_27301_, _20585_, _20584_);
  and _52949_ (_20586_, _05102_, _23824_);
  and _52950_ (_20587_, _05105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or _52951_ (_12224_, _20587_, _20586_);
  and _52952_ (_20588_, _04832_, _23778_);
  and _52953_ (_20589_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or _52954_ (_12226_, _20589_, _20588_);
  and _52955_ (_20590_, _04832_, _24050_);
  and _52956_ (_20591_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or _52957_ (_12228_, _20591_, _20590_);
  and _52958_ (_20592_, _08642_, _23747_);
  and _52959_ (_20593_, _08644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  or _52960_ (_12230_, _20593_, _20592_);
  and _52961_ (_20594_, _04832_, _23649_);
  and _52962_ (_20595_, _04834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _52963_ (_12232_, _20595_, _20594_);
  and _52964_ (_20596_, _04656_, _23649_);
  and _52965_ (_20597_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or _52966_ (_12234_, _20597_, _20596_);
  and _52967_ (_20598_, _04656_, _23898_);
  and _52968_ (_20599_, _04660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or _52969_ (_12237_, _20599_, _20598_);
  and _52970_ (_20600_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  and _52971_ (_20601_, _17775_, _23707_);
  or _52972_ (_12239_, _20601_, _20600_);
  and _52973_ (_20602_, _02087_, _23649_);
  and _52974_ (_20603_, _02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _52975_ (_12241_, _20603_, _20602_);
  and _52976_ (_20604_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  and _52977_ (_20605_, _17775_, _24050_);
  or _52978_ (_12243_, _20605_, _20604_);
  and _52979_ (_20606_, _01759_, _24050_);
  and _52980_ (_20607_, _01762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or _52981_ (_12245_, _20607_, _20606_);
  and _52982_ (_20608_, _25754_, _23707_);
  and _52983_ (_20609_, _25756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  or _52984_ (_12247_, _20609_, _20608_);
  and _52985_ (_20610_, _07514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and _52986_ (_20611_, _07513_, _23946_);
  or _52987_ (_12249_, _20611_, _20610_);
  and _52988_ (_20612_, _25571_, _23946_);
  and _52989_ (_20613_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or _52990_ (_27058_, _20613_, _20612_);
  and _52991_ (_20614_, _25571_, _23824_);
  and _52992_ (_20615_, _25573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or _52993_ (_12252_, _20615_, _20614_);
  and _52994_ (_20616_, _25488_, _23649_);
  and _52995_ (_20617_, _25490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or _52996_ (_12254_, _20617_, _20616_);
  and _52997_ (_20618_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  and _52998_ (_20619_, _17775_, _23946_);
  or _52999_ (_12256_, _20619_, _20618_);
  and _53000_ (_20620_, _25340_, _23898_);
  and _53001_ (_20621_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  or _53002_ (_12258_, _20621_, _20620_);
  and _53003_ (_20622_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and _53004_ (_20623_, _16325_, _23747_);
  or _53005_ (_12260_, _20623_, _20622_);
  and _53006_ (_20624_, _25340_, _23946_);
  and _53007_ (_20625_, _25342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  or _53008_ (_12264_, _20625_, _20624_);
  and _53009_ (_20626_, _17776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  and _53010_ (_20627_, _17775_, _23824_);
  or _53011_ (_12266_, _20627_, _20626_);
  and _53012_ (_20628_, _24358_, _23946_);
  and _53013_ (_20629_, _24360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  or _53014_ (_12268_, _20629_, _20628_);
  and _53015_ (_20630_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and _53016_ (_20631_, _16325_, _23824_);
  or _53017_ (_26967_, _20631_, _20630_);
  and _53018_ (_20632_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and _53019_ (_20633_, _17255_, _23747_);
  or _53020_ (_12273_, _20633_, _20632_);
  and _53021_ (_20634_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and _53022_ (_20635_, _17255_, _23946_);
  or _53023_ (_12277_, _20635_, _20634_);
  and _53024_ (_20636_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and _53025_ (_20637_, _16325_, _23649_);
  or _53026_ (_12280_, _20637_, _20636_);
  and _53027_ (_20638_, _08548_, _23649_);
  and _53028_ (_20639_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  or _53029_ (_12282_, _20639_, _20638_);
  and _53030_ (_20640_, _06602_, _23824_);
  and _53031_ (_20641_, _06604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  or _53032_ (_12284_, _20641_, _20640_);
  and _53033_ (_20642_, _18217_, _23898_);
  and _53034_ (_20643_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or _53035_ (_12288_, _20643_, _20642_);
  and _53036_ (_12290_, _00984_, _22762_);
  and _53037_ (_20644_, _17263_, _23707_);
  and _53038_ (_20645_, _17265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  or _53039_ (_12292_, _20645_, _20644_);
  and _53040_ (_20646_, _17256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and _53041_ (_20647_, _17255_, _23649_);
  or _53042_ (_12294_, _20647_, _20646_);
  and _53043_ (_20648_, _18217_, _23778_);
  and _53044_ (_20649_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or _53045_ (_12477_, _20649_, _20648_);
  and _53046_ (_20650_, _08548_, _24050_);
  and _53047_ (_20651_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  or _53048_ (_27137_, _20651_, _20650_);
  and _53049_ (_20652_, _25739_, _23649_);
  and _53050_ (_20653_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  or _53051_ (_12509_, _20653_, _20652_);
  and _53052_ (_20654_, _07743_, _23778_);
  and _53053_ (_20655_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  or _53054_ (_27071_, _20655_, _20654_);
  and _53055_ (_20656_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _53056_ (_20657_, _20656_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _53057_ (_20658_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and _53058_ (_20659_, _20658_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and _53059_ (_20660_, _20659_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and _53060_ (_20661_, _20660_, _20657_);
  and _53061_ (_20662_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _53062_ (_20663_, _20662_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and _53063_ (_20664_, _20663_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _53064_ (_20665_, _20664_, _20661_);
  and _53065_ (_20666_, _20665_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _53066_ (_20667_, _20666_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _53067_ (_20668_, _20667_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and _53068_ (_20669_, _20667_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _53069_ (_20670_, _20669_, _20668_);
  nor _53070_ (_20671_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not _53071_ (_20672_, _20671_);
  and _53072_ (_20673_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _22841_);
  and _53073_ (_20674_, _20656_, _22854_);
  nor _53074_ (_20675_, _20656_, _22854_);
  nor _53075_ (_20676_, _20675_, _20674_);
  nor _53076_ (_20677_, _20676_, _22841_);
  nor _53077_ (_20678_, _20677_, _20673_);
  not _53078_ (_20679_, _20678_);
  nor _53079_ (_20680_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53080_ (_20681_, _22849_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _53081_ (_20682_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _22845_);
  nor _53082_ (_20683_, _20682_, _20681_);
  and _53083_ (_20684_, _20683_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53084_ (_20685_, _20684_, _20680_);
  nor _53085_ (_20686_, _20685_, _08039_);
  and _53086_ (_20687_, _20685_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor _53087_ (_20688_, _20687_, _20686_);
  nor _53088_ (_20689_, _20688_, _20679_);
  nor _53089_ (_20690_, _20685_, _07621_);
  and _53090_ (_20691_, _20685_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _53091_ (_20692_, _20691_, _20690_);
  nor _53092_ (_20693_, _20692_, _20678_);
  nor _53093_ (_20694_, _20693_, _20689_);
  nor _53094_ (_20695_, _20694_, _20672_);
  and _53095_ (_20696_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _22841_);
  not _53096_ (_20697_, _20696_);
  nor _53097_ (_20698_, _20685_, _07600_);
  and _53098_ (_20699_, _20685_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _53099_ (_20700_, _20699_, _20698_);
  nor _53100_ (_20701_, _20700_, _20679_);
  not _53101_ (_20702_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _53102_ (_20703_, _20685_, _20702_);
  and _53103_ (_20704_, _20685_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _53104_ (_20705_, _20704_, _20703_);
  nor _53105_ (_20706_, _20705_, _20678_);
  nor _53106_ (_20707_, _20706_, _20701_);
  nor _53107_ (_20708_, _20707_, _20697_);
  nor _53108_ (_20709_, _20708_, _20695_);
  and _53109_ (_20710_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not _53110_ (_20711_, _20710_);
  not _53111_ (_20712_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _53112_ (_20713_, _20685_, _20712_);
  and _53113_ (_20714_, _20685_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _53114_ (_20715_, _20714_, _20713_);
  nor _53115_ (_20716_, _20715_, _20679_);
  nor _53116_ (_20717_, _20685_, _07665_);
  and _53117_ (_20718_, _20685_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _53118_ (_20719_, _20718_, _20717_);
  nor _53119_ (_20720_, _20719_, _20678_);
  nor _53120_ (_20721_, _20720_, _20716_);
  nor _53121_ (_20722_, _20721_, _20711_);
  and _53122_ (_20723_, _22845_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not _53123_ (_20724_, _20723_);
  nor _53124_ (_20725_, _20685_, _07657_);
  and _53125_ (_20726_, _20685_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _53126_ (_20727_, _20726_, _20725_);
  nor _53127_ (_20728_, _20727_, _20679_);
  nor _53128_ (_20729_, _20685_, _08225_);
  and _53129_ (_20730_, _20685_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _53130_ (_20731_, _20730_, _20729_);
  nor _53131_ (_20732_, _20731_, _20678_);
  nor _53132_ (_20733_, _20732_, _20728_);
  nor _53133_ (_20734_, _20733_, _20724_);
  nor _53134_ (_20735_, _20734_, _20722_);
  and _53135_ (_20736_, _20735_, _20709_);
  not _53136_ (_20737_, _20685_);
  and _53137_ (_20738_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _53138_ (_20739_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _53139_ (_20740_, _20739_, _20738_);
  and _53140_ (_20741_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _53141_ (_20742_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _53142_ (_20743_, _20742_, _20741_);
  and _53143_ (_20744_, _20743_, _20740_);
  and _53144_ (_20745_, _20744_, _20737_);
  and _53145_ (_20746_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _53146_ (_20747_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor _53147_ (_20748_, _20747_, _20746_);
  and _53148_ (_20749_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _53149_ (_20750_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _53150_ (_20751_, _20750_, _20749_);
  and _53151_ (_20752_, _20751_, _20748_);
  and _53152_ (_20753_, _20752_, _20685_);
  or _53153_ (_20754_, _20753_, _20679_);
  nor _53154_ (_20755_, _20754_, _20745_);
  and _53155_ (_20756_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _53156_ (_20757_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor _53157_ (_20758_, _20757_, _20756_);
  and _53158_ (_20759_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _53159_ (_20760_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor _53160_ (_20761_, _20760_, _20759_);
  and _53161_ (_20762_, _20761_, _20758_);
  nor _53162_ (_20763_, _20762_, _20685_);
  and _53163_ (_20764_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _53164_ (_20765_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _53165_ (_20766_, _20765_, _20764_);
  and _53166_ (_20767_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _53167_ (_20768_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _53168_ (_20769_, _20768_, _20767_);
  and _53169_ (_20770_, _20769_, _20766_);
  nor _53170_ (_20771_, _20770_, _20737_);
  or _53171_ (_20772_, _20771_, _20763_);
  and _53172_ (_20773_, _20772_, _20679_);
  nor _53173_ (_20774_, _20773_, _20755_);
  nor _53174_ (_20775_, _20774_, _20736_);
  and _53175_ (_20776_, _20775_, _20670_);
  nor _53176_ (_20777_, _20666_, _22897_);
  and _53177_ (_20778_, _20663_, _20661_);
  and _53178_ (_20779_, _20778_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _53179_ (_20780_, _20779_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _53180_ (_20781_, _20780_, _22897_);
  nor _53181_ (_20782_, _20781_, _20777_);
  not _53182_ (_20783_, _20782_);
  and _53183_ (_20784_, _20783_, _20775_);
  nor _53184_ (_20785_, _20665_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _53185_ (_20786_, _20785_, _20666_);
  and _53186_ (_20787_, _20786_, _20775_);
  nor _53187_ (_20788_, _20783_, _20775_);
  nor _53188_ (_20789_, _20788_, _20784_);
  nor _53189_ (_20790_, _20778_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _53190_ (_20791_, _20790_, _20779_);
  and _53191_ (_20792_, _20791_, _20775_);
  nor _53192_ (_20793_, _20791_, _20775_);
  and _53193_ (_20794_, _20662_, _20661_);
  nor _53194_ (_20795_, _20794_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _53195_ (_20796_, _20795_, _20778_);
  and _53196_ (_20797_, _20796_, _20775_);
  nor _53197_ (_20798_, _20796_, _20775_);
  nor _53198_ (_20799_, _20798_, _20797_);
  and _53199_ (_20800_, _20661_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _53200_ (_20801_, _20800_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _53201_ (_20802_, _20801_, _20794_);
  and _53202_ (_20803_, _20802_, _20775_);
  nor _53203_ (_20804_, _20802_, _20775_);
  nor _53204_ (_20805_, _20661_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _53205_ (_20806_, _20805_, _20800_);
  and _53206_ (_20807_, _20806_, _20775_);
  and _53207_ (_20808_, _20659_, _20657_);
  nor _53208_ (_20809_, _20808_, _22874_);
  and _53209_ (_20810_, _20808_, _22874_);
  nor _53210_ (_20811_, _20810_, _20809_);
  not _53211_ (_20812_, _20811_);
  and _53212_ (_20813_, _20812_, _20775_);
  nor _53213_ (_20814_, _20812_, _20775_);
  and _53214_ (_20815_, _20658_, _20657_);
  nor _53215_ (_20816_, _20815_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _53216_ (_20817_, _20816_, _20808_);
  and _53217_ (_20818_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _53218_ (_20819_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _53219_ (_20820_, _20819_, _20818_);
  and _53220_ (_20821_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _53221_ (_20822_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _53222_ (_20823_, _20822_, _20821_);
  and _53223_ (_20824_, _20823_, _20820_);
  and _53224_ (_20825_, _20824_, _20685_);
  and _53225_ (_20826_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _53226_ (_20827_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _53227_ (_20828_, _20827_, _20826_);
  and _53228_ (_20829_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _53229_ (_20830_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _53230_ (_20831_, _20830_, _20829_);
  and _53231_ (_20832_, _20831_, _20828_);
  and _53232_ (_20833_, _20832_, _20737_);
  or _53233_ (_20834_, _20833_, _20679_);
  nor _53234_ (_20835_, _20834_, _20825_);
  and _53235_ (_20836_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _53236_ (_20837_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _53237_ (_20838_, _20837_, _20836_);
  and _53238_ (_20839_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _53239_ (_20840_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _53240_ (_20841_, _20840_, _20839_);
  and _53241_ (_20842_, _20841_, _20838_);
  nor _53242_ (_20843_, _20842_, _20685_);
  and _53243_ (_20844_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _53244_ (_20845_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _53245_ (_20846_, _20845_, _20844_);
  and _53246_ (_20847_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _53247_ (_20848_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _53248_ (_20849_, _20848_, _20847_);
  and _53249_ (_20850_, _20849_, _20846_);
  nor _53250_ (_20851_, _20850_, _20737_);
  or _53251_ (_20852_, _20851_, _20843_);
  and _53252_ (_20853_, _20852_, _20679_);
  nor _53253_ (_20854_, _20853_, _20835_);
  nor _53254_ (_20855_, _20854_, _20736_);
  and _53255_ (_20856_, _20855_, _20817_);
  nor _53256_ (_20857_, _20855_, _20817_);
  nor _53257_ (_20858_, _20857_, _20856_);
  not _53258_ (_20859_, _20858_);
  and _53259_ (_20860_, _20657_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _53260_ (_20861_, _20860_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _53261_ (_20862_, _20861_, _20815_);
  and _53262_ (_20863_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _53263_ (_20864_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _53264_ (_20865_, _20864_, _20863_);
  and _53265_ (_20866_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _53266_ (_20867_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _53267_ (_20868_, _20867_, _20866_);
  and _53268_ (_20869_, _20868_, _20865_);
  and _53269_ (_20870_, _20869_, _20737_);
  and _53270_ (_20871_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _53271_ (_20872_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _53272_ (_20873_, _20872_, _20871_);
  and _53273_ (_20874_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _53274_ (_20875_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _53275_ (_20876_, _20875_, _20874_);
  and _53276_ (_20877_, _20876_, _20873_);
  and _53277_ (_20878_, _20877_, _20685_);
  or _53278_ (_20879_, _20878_, _20679_);
  nor _53279_ (_20880_, _20879_, _20870_);
  and _53280_ (_20881_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _53281_ (_20882_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _53282_ (_20883_, _20882_, _20881_);
  and _53283_ (_20884_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _53284_ (_20885_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _53285_ (_20886_, _20885_, _20884_);
  and _53286_ (_20887_, _20886_, _20883_);
  and _53287_ (_20888_, _20887_, _20737_);
  and _53288_ (_20889_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _53289_ (_20890_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _53290_ (_20891_, _20890_, _20889_);
  and _53291_ (_20892_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _53292_ (_20893_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _53293_ (_20894_, _20893_, _20892_);
  and _53294_ (_20895_, _20894_, _20891_);
  and _53295_ (_20896_, _20895_, _20685_);
  nor _53296_ (_20897_, _20896_, _20888_);
  and _53297_ (_20898_, _20897_, _20679_);
  nor _53298_ (_20899_, _20898_, _20880_);
  nor _53299_ (_20900_, _20899_, _20736_);
  and _53300_ (_20901_, _20900_, _20862_);
  nor _53301_ (_20902_, _20900_, _20862_);
  nor _53302_ (_20903_, _20902_, _20901_);
  not _53303_ (_20904_, _20903_);
  and _53304_ (_20905_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _53305_ (_20906_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _53306_ (_20907_, _20906_, _20905_);
  and _53307_ (_20908_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _53308_ (_20909_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _53309_ (_20910_, _20909_, _20908_);
  and _53310_ (_20911_, _20910_, _20907_);
  and _53311_ (_20912_, _20911_, _20737_);
  and _53312_ (_20913_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _53313_ (_20914_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _53314_ (_20915_, _20914_, _20913_);
  and _53315_ (_20916_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _53316_ (_20917_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _53317_ (_20918_, _20917_, _20916_);
  and _53318_ (_20919_, _20918_, _20915_);
  and _53319_ (_20920_, _20919_, _20685_);
  or _53320_ (_20921_, _20920_, _20679_);
  nor _53321_ (_20922_, _20921_, _20912_);
  and _53322_ (_20923_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _53323_ (_20924_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _53324_ (_20925_, _20924_, _20923_);
  and _53325_ (_20926_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _53326_ (_20927_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _53327_ (_20928_, _20927_, _20926_);
  and _53328_ (_20929_, _20928_, _20925_);
  nor _53329_ (_20930_, _20929_, _20685_);
  and _53330_ (_20931_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _53331_ (_20932_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _53332_ (_20933_, _20932_, _20931_);
  and _53333_ (_20934_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _53334_ (_20935_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _53335_ (_20936_, _20935_, _20934_);
  and _53336_ (_20937_, _20936_, _20933_);
  nor _53337_ (_20938_, _20937_, _20737_);
  or _53338_ (_20939_, _20938_, _20930_);
  and _53339_ (_20940_, _20939_, _20679_);
  nor _53340_ (_20941_, _20940_, _20922_);
  nor _53341_ (_20942_, _20941_, _20736_);
  nor _53342_ (_20943_, _20657_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _53343_ (_20944_, _20943_, _20860_);
  and _53344_ (_20945_, _20944_, _20942_);
  not _53345_ (_20946_, _20676_);
  and _53346_ (_20947_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _53347_ (_20948_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _53348_ (_20949_, _20948_, _20947_);
  and _53349_ (_20950_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _53350_ (_20951_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _53351_ (_20952_, _20951_, _20950_);
  and _53352_ (_20953_, _20952_, _20949_);
  and _53353_ (_20954_, _20953_, _20737_);
  and _53354_ (_20955_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _53355_ (_20956_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _53356_ (_20957_, _20956_, _20955_);
  and _53357_ (_20958_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _53358_ (_20959_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _53359_ (_20960_, _20959_, _20958_);
  and _53360_ (_20961_, _20960_, _20957_);
  and _53361_ (_20962_, _20961_, _20685_);
  or _53362_ (_20963_, _20962_, _20679_);
  nor _53363_ (_20964_, _20963_, _20954_);
  and _53364_ (_20965_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _53365_ (_20966_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _53366_ (_20967_, _20966_, _20965_);
  and _53367_ (_20968_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _53368_ (_20969_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _53369_ (_20970_, _20969_, _20968_);
  and _53370_ (_20971_, _20970_, _20967_);
  nor _53371_ (_20972_, _20971_, _20685_);
  and _53372_ (_20973_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _53373_ (_20974_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _53374_ (_20975_, _20974_, _20973_);
  and _53375_ (_20976_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _53376_ (_20977_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _53377_ (_20978_, _20977_, _20976_);
  and _53378_ (_20979_, _20978_, _20975_);
  nor _53379_ (_20980_, _20979_, _20737_);
  or _53380_ (_20981_, _20980_, _20972_);
  and _53381_ (_20982_, _20981_, _20679_);
  nor _53382_ (_20983_, _20982_, _20964_);
  nor _53383_ (_20984_, _20983_, _20736_);
  and _53384_ (_20985_, _20984_, _20946_);
  nor _53385_ (_20986_, _20984_, _20946_);
  nor _53386_ (_20987_, _20986_, _20985_);
  not _53387_ (_20988_, _20987_);
  not _53388_ (_20989_, _20683_);
  and _53389_ (_20990_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _53390_ (_20991_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _53391_ (_20992_, _20991_, _20990_);
  and _53392_ (_20993_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _53393_ (_20994_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _53394_ (_20995_, _20994_, _20993_);
  and _53395_ (_20996_, _20995_, _20992_);
  and _53396_ (_20997_, _20996_, _20737_);
  and _53397_ (_20998_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _53398_ (_20999_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _53399_ (_21000_, _20999_, _20998_);
  and _53400_ (_21001_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _53401_ (_21002_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _53402_ (_21003_, _21002_, _21001_);
  and _53403_ (_21004_, _21003_, _21000_);
  and _53404_ (_21005_, _21004_, _20685_);
  or _53405_ (_21006_, _21005_, _20679_);
  nor _53406_ (_21007_, _21006_, _20997_);
  and _53407_ (_21008_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _53408_ (_21009_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _53409_ (_21010_, _21009_, _21008_);
  and _53410_ (_21011_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _53411_ (_21012_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _53412_ (_21013_, _21012_, _21011_);
  and _53413_ (_21014_, _21013_, _21010_);
  and _53414_ (_21015_, _21014_, _20737_);
  and _53415_ (_21016_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _53416_ (_21017_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _53417_ (_21018_, _21017_, _21016_);
  and _53418_ (_21019_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _53419_ (_21020_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _53420_ (_21021_, _21020_, _21019_);
  and _53421_ (_21022_, _21021_, _21018_);
  and _53422_ (_21023_, _21022_, _20685_);
  nor _53423_ (_21024_, _21023_, _21015_);
  and _53424_ (_21025_, _21024_, _20679_);
  nor _53425_ (_21026_, _21025_, _21007_);
  nor _53426_ (_21027_, _21026_, _20736_);
  and _53427_ (_21028_, _21027_, _20989_);
  and _53428_ (_21029_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _53429_ (_21030_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _53430_ (_21031_, _21030_, _21029_);
  and _53431_ (_21032_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _53432_ (_21033_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _53433_ (_21034_, _21033_, _21032_);
  and _53434_ (_21035_, _21034_, _21031_);
  and _53435_ (_21036_, _21035_, _20737_);
  and _53436_ (_21037_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _53437_ (_21038_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _53438_ (_21039_, _21038_, _21037_);
  and _53439_ (_21040_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _53440_ (_21041_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _53441_ (_21042_, _21041_, _21040_);
  and _53442_ (_21043_, _21042_, _21039_);
  and _53443_ (_21044_, _21043_, _20685_);
  or _53444_ (_21045_, _21044_, _20679_);
  nor _53445_ (_21046_, _21045_, _21036_);
  and _53446_ (_21047_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _53447_ (_21048_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _53448_ (_21049_, _21048_, _21047_);
  and _53449_ (_21050_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _53450_ (_21051_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _53451_ (_21052_, _21051_, _21050_);
  and _53452_ (_21053_, _21052_, _21049_);
  nor _53453_ (_21054_, _21053_, _20685_);
  and _53454_ (_21055_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _53455_ (_21056_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _53456_ (_21057_, _21056_, _21055_);
  and _53457_ (_21058_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _53458_ (_21059_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _53459_ (_21060_, _21059_, _21058_);
  and _53460_ (_21061_, _21060_, _21057_);
  nor _53461_ (_21062_, _21061_, _20737_);
  or _53462_ (_21063_, _21062_, _21054_);
  and _53463_ (_21064_, _21063_, _20679_);
  nor _53464_ (_21065_, _21064_, _21046_);
  nor _53465_ (_21066_, _21065_, _20736_);
  and _53466_ (_21067_, _21066_, _22845_);
  and _53467_ (_21068_, _20696_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _53468_ (_21069_, _20710_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _53469_ (_21070_, _21069_, _21068_);
  and _53470_ (_21071_, _20723_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _53471_ (_21072_, _20671_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor _53472_ (_21073_, _21072_, _21071_);
  and _53473_ (_21074_, _21073_, _21070_);
  and _53474_ (_21075_, _21074_, _20737_);
  and _53475_ (_21076_, _20696_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _53476_ (_21077_, _20671_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _53477_ (_21078_, _21077_, _21076_);
  and _53478_ (_21079_, _20723_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _53479_ (_21080_, _20710_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _53480_ (_21081_, _21080_, _21079_);
  and _53481_ (_21082_, _21081_, _21078_);
  and _53482_ (_21083_, _21082_, _20685_);
  or _53483_ (_21084_, _21083_, _20679_);
  nor _53484_ (_21085_, _21084_, _21075_);
  and _53485_ (_21086_, _20696_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _53486_ (_21087_, _20671_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _53487_ (_21088_, _21087_, _21086_);
  and _53488_ (_21089_, _20723_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _53489_ (_21090_, _20710_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _53490_ (_21091_, _21090_, _21089_);
  and _53491_ (_21092_, _21091_, _21088_);
  and _53492_ (_21093_, _21092_, _20737_);
  and _53493_ (_21094_, _20723_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _53494_ (_21095_, _20710_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _53495_ (_21096_, _21095_, _21094_);
  and _53496_ (_21097_, _20696_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _53497_ (_21098_, _20671_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _53498_ (_21099_, _21098_, _21097_);
  and _53499_ (_21100_, _21099_, _21096_);
  and _53500_ (_21101_, _21100_, _20685_);
  nor _53501_ (_21102_, _21101_, _21093_);
  and _53502_ (_21103_, _21102_, _20679_);
  nor _53503_ (_21104_, _21103_, _21085_);
  nor _53504_ (_21105_, _21104_, _20736_);
  and _53505_ (_21106_, _21105_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53506_ (_21107_, _21066_, _22845_);
  nor _53507_ (_21108_, _21107_, _21067_);
  and _53508_ (_21109_, _21108_, _21106_);
  nor _53509_ (_21110_, _21109_, _21067_);
  nor _53510_ (_21111_, _21027_, _20989_);
  nor _53511_ (_21112_, _21111_, _21028_);
  not _53512_ (_21113_, _21112_);
  nor _53513_ (_21114_, _21113_, _21110_);
  nor _53514_ (_21115_, _21114_, _21028_);
  nor _53515_ (_21116_, _21115_, _20988_);
  nor _53516_ (_21117_, _21116_, _20985_);
  nor _53517_ (_21118_, _20944_, _20942_);
  nor _53518_ (_21119_, _21118_, _20945_);
  not _53519_ (_21120_, _21119_);
  nor _53520_ (_21121_, _21120_, _21117_);
  nor _53521_ (_21122_, _21121_, _20945_);
  nor _53522_ (_21123_, _21122_, _20904_);
  nor _53523_ (_21124_, _21123_, _20901_);
  nor _53524_ (_21125_, _21124_, _20859_);
  nor _53525_ (_21126_, _21125_, _20856_);
  nor _53526_ (_21127_, _21126_, _20814_);
  or _53527_ (_21128_, _21127_, _20813_);
  nor _53528_ (_21129_, _20806_, _20775_);
  nor _53529_ (_21130_, _21129_, _20807_);
  and _53530_ (_21131_, _21130_, _21128_);
  nor _53531_ (_21132_, _21131_, _20807_);
  nor _53532_ (_21133_, _21132_, _20804_);
  or _53533_ (_21134_, _21133_, _20803_);
  and _53534_ (_21135_, _21134_, _20799_);
  nor _53535_ (_21136_, _21135_, _20797_);
  nor _53536_ (_21137_, _21136_, _20793_);
  or _53537_ (_21138_, _21137_, _20792_);
  nor _53538_ (_21139_, _20786_, _20775_);
  nor _53539_ (_21140_, _21139_, _20787_);
  and _53540_ (_21141_, _21140_, _21138_);
  and _53541_ (_21142_, _21141_, _20789_);
  or _53542_ (_21143_, _21142_, _20787_);
  nor _53543_ (_21144_, _21143_, _20784_);
  nor _53544_ (_21145_, _20775_, _20670_);
  nor _53545_ (_21146_, _21145_, _20776_);
  not _53546_ (_21147_, _21146_);
  nor _53547_ (_21148_, _21147_, _21144_);
  nor _53548_ (_21149_, _21148_, _20776_);
  nor _53549_ (_21150_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _53550_ (_21151_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _53551_ (_21152_, _21151_, _21150_);
  not _53552_ (_21153_, _21152_);
  nor _53553_ (_21154_, _21153_, _20669_);
  and _53554_ (_21155_, _21153_, _20669_);
  nor _53555_ (_21156_, _21155_, _21154_);
  not _53556_ (_21157_, _21156_);
  and _53557_ (_21158_, _21157_, _20775_);
  nor _53558_ (_21159_, _21157_, _20775_);
  nor _53559_ (_21160_, _21159_, _21158_);
  not _53560_ (_21161_, _21160_);
  nand _53561_ (_21162_, _21161_, _21149_);
  or _53562_ (_21163_, _21161_, _21149_);
  and _53563_ (_21164_, _21163_, _21162_);
  and _53564_ (_21165_, _21147_, _21144_);
  nor _53565_ (_21166_, _21165_, _21148_);
  nor _53566_ (_21167_, _21166_, _22837_);
  and _53567_ (_21168_, _21166_, _22837_);
  nor _53568_ (_21169_, _21141_, _20787_);
  and _53569_ (_21170_, _20789_, _22832_);
  nor _53570_ (_21171_, _20789_, _22832_);
  nor _53571_ (_21172_, _21171_, _21170_);
  nand _53572_ (_21173_, _21172_, _21169_);
  or _53573_ (_21174_, _21172_, _21169_);
  and _53574_ (_21175_, _21174_, _21173_);
  nor _53575_ (_21176_, _21140_, _21138_);
  nor _53576_ (_21177_, _21176_, _21141_);
  nor _53577_ (_21178_, _21177_, _22827_);
  and _53578_ (_21179_, _21177_, _22827_);
  nor _53579_ (_21180_, _20791_, _22823_);
  and _53580_ (_21181_, _20791_, _22823_);
  or _53581_ (_21182_, _21181_, _21180_);
  nand _53582_ (_21183_, _21182_, _20775_);
  or _53583_ (_21184_, _21182_, _20775_);
  and _53584_ (_21185_, _21184_, _21183_);
  not _53585_ (_21186_, _21185_);
  nand _53586_ (_21187_, _21186_, _21136_);
  or _53587_ (_21188_, _21186_, _21136_);
  and _53588_ (_21189_, _21188_, _21187_);
  nor _53589_ (_21190_, _21134_, _20799_);
  nor _53590_ (_21191_, _21190_, _21135_);
  nor _53591_ (_21192_, _21191_, _22819_);
  and _53592_ (_21193_, _21191_, _22819_);
  not _53593_ (_21194_, _20775_);
  nor _53594_ (_21195_, _20802_, _22814_);
  and _53595_ (_21196_, _20802_, _22814_);
  or _53596_ (_21197_, _21196_, _21195_);
  nand _53597_ (_21198_, _21197_, _21194_);
  or _53598_ (_21199_, _21197_, _21194_);
  and _53599_ (_21200_, _21199_, _21198_);
  or _53600_ (_21201_, _21200_, _21132_);
  nand _53601_ (_21202_, _21200_, _21132_);
  and _53602_ (_21203_, _21202_, _21201_);
  nor _53603_ (_21204_, _20813_, _20814_);
  nor _53604_ (_21205_, _21204_, _21126_);
  and _53605_ (_21206_, _21204_, _21126_);
  or _53606_ (_21207_, _21206_, _21205_);
  nor _53607_ (_21208_, _21207_, _22806_);
  and _53608_ (_21209_, _21207_, _22806_);
  and _53609_ (_21210_, _21124_, _20859_);
  nor _53610_ (_21211_, _21210_, _21125_);
  and _53611_ (_21212_, _21211_, _22802_);
  nor _53612_ (_21213_, _21211_, _22802_);
  and _53613_ (_21214_, _21122_, _20904_);
  nor _53614_ (_21215_, _21214_, _21123_);
  nor _53615_ (_21216_, _21215_, _22798_);
  and _53616_ (_21217_, _21215_, _22798_);
  and _53617_ (_21218_, _21120_, _21117_);
  nor _53618_ (_21219_, _21218_, _21121_);
  and _53619_ (_21220_, _21219_, _22794_);
  and _53620_ (_21221_, _21115_, _20988_);
  nor _53621_ (_21222_, _21221_, _21116_);
  and _53622_ (_21223_, _21222_, _22788_);
  nor _53623_ (_21224_, _21222_, _22788_);
  and _53624_ (_21225_, _21113_, _21110_);
  nor _53625_ (_21226_, _21225_, _21114_);
  nor _53626_ (_21227_, _21226_, _22783_);
  nor _53627_ (_21228_, _21108_, _21106_);
  nor _53628_ (_21229_, _21228_, _21109_);
  nor _53629_ (_21230_, _21229_, _22778_);
  and _53630_ (_21231_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _53631_ (_21232_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _53632_ (_21233_, _21232_, _21231_);
  and _53633_ (_21234_, _21233_, _21105_);
  nor _53634_ (_21235_, _21233_, _21105_);
  or _53635_ (_21236_, _21235_, _21234_);
  and _53636_ (_21237_, _21229_, _22778_);
  or _53637_ (_21238_, _21237_, _21236_);
  or _53638_ (_21239_, _21238_, _21230_);
  and _53639_ (_21240_, _21226_, _22783_);
  or _53640_ (_21241_, _21240_, _21239_);
  or _53641_ (_21242_, _21241_, _21227_);
  or _53642_ (_21243_, _21242_, _21224_);
  or _53643_ (_21244_, _21243_, _21223_);
  nor _53644_ (_21245_, _21219_, _22794_);
  or _53645_ (_21246_, _21245_, _21244_);
  or _53646_ (_21248_, _21246_, _21220_);
  or _53647_ (_21249_, _21248_, _21217_);
  or _53648_ (_21250_, _21249_, _21216_);
  or _53649_ (_21251_, _21250_, _21213_);
  or _53650_ (_21252_, _21251_, _21212_);
  or _53651_ (_21253_, _21252_, _21209_);
  or _53652_ (_21254_, _21253_, _21208_);
  nor _53653_ (_21255_, _21130_, _21128_);
  nor _53654_ (_21256_, _21255_, _21131_);
  nor _53655_ (_21257_, _21256_, _22810_);
  and _53656_ (_21258_, _21256_, _22810_);
  or _53657_ (_21259_, _21258_, _21257_);
  or _53658_ (_21260_, _21259_, _21254_);
  or _53659_ (_21261_, _21260_, _21203_);
  or _53660_ (_21262_, _21261_, _21193_);
  or _53661_ (_21263_, _21262_, _21192_);
  or _53662_ (_21264_, _21263_, _21189_);
  or _53663_ (_21265_, _21264_, _21179_);
  or _53664_ (_21266_, _21265_, _21178_);
  or _53665_ (_21267_, _21266_, _21175_);
  or _53666_ (_21268_, _21267_, _21168_);
  or _53667_ (_21269_, _21268_, _21167_);
  or _53668_ (_21270_, _21269_, _21164_);
  and _53669_ (_21271_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _53670_ (_21272_, _21271_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _53671_ (_21273_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _53672_ (_21274_, _21273_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _53673_ (_21275_, _21274_, _21272_);
  not _53674_ (_21276_, _21275_);
  nor _53675_ (_21277_, _21272_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _53676_ (_21278_, _21272_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _53677_ (_21279_, _21278_, _21277_);
  nand _53678_ (_21280_, _21279_, _20702_);
  or _53679_ (_21281_, _21279_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _53680_ (_21282_, _21281_, _21280_);
  and _53681_ (_21283_, _21282_, _21276_);
  nand _53682_ (_21284_, _21279_, _07612_);
  or _53683_ (_21285_, _21279_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _53684_ (_21286_, _21285_, _21275_);
  and _53685_ (_21287_, _21286_, _21284_);
  or _53686_ (_21288_, _21287_, _21283_);
  or _53687_ (_21289_, _21288_, _22778_);
  and _53688_ (_21290_, _22783_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _53689_ (_21291_, \oc8051_symbolic_cxrom1.regvalid [5], _22788_);
  and _53690_ (_21292_, \oc8051_symbolic_cxrom1.regvalid [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _53691_ (_21293_, _21292_, _21291_);
  and _53692_ (_21294_, _21293_, _21290_);
  or _53693_ (_21295_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _53694_ (_21296_, \oc8051_symbolic_cxrom1.regvalid [1], _22788_);
  and _53695_ (_21297_, _21296_, _21271_);
  and _53696_ (_21298_, _21297_, _21295_);
  or _53697_ (_21299_, _21298_, _21294_);
  nor _53698_ (_21300_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _53699_ (_21301_, _21300_, _22783_);
  nor _53700_ (_21302_, _21301_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _53701_ (_21303_, _21301_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _53702_ (_21304_, _21303_, _21302_);
  and _53703_ (_21305_, _21304_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _53704_ (_21306_, _21300_, _22783_);
  nor _53705_ (_21307_, _21306_, _21301_);
  or _53706_ (_21308_, _08145_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _53707_ (_21309_, _21308_, _21307_);
  or _53708_ (_21310_, _21309_, _21305_);
  and _53709_ (_21311_, _21310_, _22778_);
  nor _53710_ (_21312_, _21304_, _07600_);
  and _53711_ (_21313_, _21304_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _53712_ (_21314_, _21313_, _21312_);
  or _53713_ (_21315_, _21314_, _21307_);
  and _53714_ (_21316_, _21315_, _21311_);
  or _53715_ (_21317_, _21316_, _21299_);
  and _53716_ (_21318_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _53717_ (_21319_, \oc8051_symbolic_cxrom1.regvalid [0], _22788_);
  or _53718_ (_21320_, _21319_, _21318_);
  and _53719_ (_21321_, _21320_, _22783_);
  and _53720_ (_21322_, \oc8051_symbolic_cxrom1.regvalid [4], _22788_);
  and _53721_ (_21323_, \oc8051_symbolic_cxrom1.regvalid [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _53722_ (_21324_, _21323_, _21322_);
  and _53723_ (_21325_, _21324_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _53724_ (_21326_, _21325_, _21321_);
  or _53725_ (_21327_, _21326_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _53726_ (_21328_, _21290_, _21324_);
  or _53727_ (_21329_, \oc8051_symbolic_cxrom1.regvalid [0], _22788_);
  or _53728_ (_21330_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _53729_ (_21331_, _21330_, _21271_);
  and _53730_ (_21332_, _21331_, _21329_);
  or _53731_ (_21333_, _21332_, _21328_);
  and _53732_ (_21334_, \oc8051_symbolic_cxrom1.regvalid [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _53733_ (_21335_, \oc8051_symbolic_cxrom1.regvalid [6], _22788_);
  or _53734_ (_21336_, _21335_, _22783_);
  or _53735_ (_21337_, _21336_, _21334_);
  or _53736_ (_21338_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _53737_ (_21339_, \oc8051_symbolic_cxrom1.regvalid [10], _22788_);
  and _53738_ (_21340_, _21339_, _21338_);
  or _53739_ (_21341_, _21340_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _53740_ (_21342_, _21341_, _21337_);
  and _53741_ (_21343_, _21342_, _22778_);
  or _53742_ (_21344_, _21343_, _21333_);
  or _53743_ (_21345_, _21342_, _22778_);
  and _53744_ (_21346_, _21345_, _22772_);
  and _53745_ (_21347_, _21346_, _21344_);
  and _53746_ (_21349_, _21347_, _21327_);
  nand _53747_ (_21350_, _21279_, _07621_);
  or _53748_ (_21351_, _21279_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _53749_ (_21352_, _21351_, _21350_);
  and _53750_ (_21353_, _21352_, _21276_);
  nand _53751_ (_21354_, _21279_, _07572_);
  or _53752_ (_21355_, _21279_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _53753_ (_21356_, _21355_, _21275_);
  and _53754_ (_21357_, _21356_, _21354_);
  or _53755_ (_21358_, _21357_, _21353_);
  or _53756_ (_21359_, _21358_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _53757_ (_21360_, _21359_, _21349_);
  and _53758_ (_21361_, _21360_, _21317_);
  and _53759_ (_21362_, _21361_, _21289_);
  or _53760_ (_21363_, \oc8051_symbolic_cxrom1.regvalid [10], _22778_);
  or _53761_ (_21364_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _53762_ (_21365_, _21364_, _21363_);
  nand _53763_ (_21366_, _21365_, _21304_);
  or _53764_ (_21367_, \oc8051_symbolic_cxrom1.regvalid [2], _22778_);
  or _53765_ (_21368_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _53766_ (_21369_, _21368_, _21367_);
  or _53767_ (_21370_, _21369_, _21304_);
  and _53768_ (_21371_, _21370_, _21366_);
  or _53769_ (_21372_, _21371_, _21307_);
  nor _53770_ (_21373_, _21279_, _20712_);
  and _53771_ (_21374_, _21279_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _53772_ (_21375_, _21374_, _21373_);
  and _53773_ (_21376_, _21375_, _21276_);
  or _53774_ (_21377_, _21279_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _53775_ (_21378_, \oc8051_symbolic_cxrom1.regvalid [12], _22788_);
  and _53776_ (_21379_, _21378_, _21275_);
  and _53777_ (_21380_, _21379_, _21377_);
  or _53778_ (_21381_, _21380_, _22778_);
  or _53779_ (_21382_, _21381_, _21376_);
  nand _53780_ (_21383_, \oc8051_symbolic_cxrom1.regvalid [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _53781_ (_21384_, _21383_, _21308_);
  or _53782_ (_21385_, _21384_, _22783_);
  or _53783_ (_21386_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _53784_ (_21387_, \oc8051_symbolic_cxrom1.regvalid [11], _22788_);
  and _53785_ (_21388_, _21387_, _21386_);
  or _53786_ (_21389_, _21388_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _53787_ (_21390_, _21389_, _21385_);
  and _53788_ (_21391_, _21390_, _21273_);
  and _53789_ (_21392_, _22778_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _53790_ (_21393_, _21293_, _22783_);
  or _53791_ (_21394_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _53792_ (_21395_, \oc8051_symbolic_cxrom1.regvalid [9], _22788_);
  and _53793_ (_21396_, _21395_, _21394_);
  or _53794_ (_21397_, _21396_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _53795_ (_21398_, _21397_, _21393_);
  and _53796_ (_21399_, _21398_, _21392_);
  or _53797_ (_21400_, _21399_, _21391_);
  and _53798_ (_21401_, _21390_, _22778_);
  or _53799_ (_21402_, _21401_, _21299_);
  and _53800_ (_21403_, _21402_, _21400_);
  and _53801_ (_21404_, _21403_, _21382_);
  and _53802_ (_21405_, _21404_, _21372_);
  or _53803_ (_21406_, _21279_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _53804_ (_21407_, \oc8051_symbolic_cxrom1.regvalid [14], _22788_);
  and _53805_ (_21408_, _21407_, _21406_);
  or _53806_ (_21409_, _21408_, _21276_);
  nand _53807_ (_21410_, _21279_, _08225_);
  or _53808_ (_21411_, _21279_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _53809_ (_21412_, _21411_, _21410_);
  or _53810_ (_21413_, _21412_, _21275_);
  and _53811_ (_21414_, _21413_, _21409_);
  or _53812_ (_21415_, _21414_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _53813_ (_21416_, _21304_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or _53814_ (_21417_, _21335_, _22778_);
  or _53815_ (_21418_, _21417_, _21416_);
  and _53816_ (_21420_, _21304_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _53817_ (_21421_, _21322_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _53818_ (_21422_, _21421_, _21420_);
  nand _53819_ (_21423_, _21422_, _21418_);
  nand _53820_ (_21424_, _21423_, _21307_);
  and _53821_ (_21425_, _21424_, _21415_);
  and _53822_ (_21426_, _21425_, _21405_);
  or _53823_ (_21427_, _21426_, _21362_);
  nor _53824_ (_21428_, _20671_, _22849_);
  and _53825_ (_21429_, _20680_, _22845_);
  nor _53826_ (_21430_, _21429_, _21428_);
  not _53827_ (_21431_, _21430_);
  and _53828_ (_21432_, _21428_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53829_ (_21433_, _21428_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53830_ (_21434_, _21433_, _21432_);
  and _53831_ (_21435_, _21434_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _53832_ (_21436_, _21434_, _07600_);
  or _53833_ (_21437_, _21436_, _21435_);
  and _53834_ (_21438_, _21437_, _21431_);
  nand _53835_ (_21439_, _21434_, _07612_);
  nor _53836_ (_21440_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53837_ (_21441_, _21440_, _21431_);
  and _53838_ (_21442_, _21441_, _21439_);
  or _53839_ (_21443_, _21442_, _21438_);
  and _53840_ (_21444_, _21443_, _20671_);
  and _53841_ (_21445_, _21434_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _53842_ (_21446_, _21434_, _20712_);
  or _53843_ (_21447_, _21446_, _21445_);
  and _53844_ (_21448_, _21447_, _21431_);
  or _53845_ (_21449_, _21434_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _53846_ (_21450_, \oc8051_symbolic_cxrom1.regvalid [12], _22854_);
  nor _53847_ (_21451_, _21450_, _21431_);
  and _53848_ (_21452_, _21451_, _21449_);
  or _53849_ (_21453_, _21452_, _21448_);
  and _53850_ (_21454_, _21453_, _20723_);
  or _53851_ (_21455_, _21454_, _21444_);
  and _53852_ (_21456_, _21434_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _53853_ (_21457_, _21434_, _07657_);
  or _53854_ (_21458_, _21457_, _21456_);
  and _53855_ (_21459_, _21458_, _21431_);
  or _53856_ (_21460_, _21434_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _53857_ (_21461_, _07637_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53858_ (_21462_, _21461_, _21431_);
  and _53859_ (_21463_, _21462_, _21460_);
  or _53860_ (_21464_, _21463_, _21459_);
  and _53861_ (_21465_, _21464_, _20710_);
  and _53862_ (_21466_, _21434_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _53863_ (_21467_, _21434_, _08039_);
  or _53864_ (_21468_, _21467_, _21466_);
  and _53865_ (_21469_, _21468_, _21431_);
  nand _53866_ (_21470_, _21434_, _07572_);
  nor _53867_ (_21471_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53868_ (_21472_, _21471_, _21431_);
  and _53869_ (_21473_, _21472_, _21470_);
  or _53870_ (_21474_, _21473_, _21469_);
  and _53871_ (_21475_, _21474_, _20696_);
  or _53872_ (_21476_, _21475_, _21465_);
  or _53873_ (_21477_, _21476_, _21455_);
  and _53874_ (_21478_, _07612_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _53875_ (_21479_, _21478_);
  nor _53876_ (_21480_, _21440_, _22849_);
  and _53877_ (_21481_, _21480_, _21479_);
  and _53878_ (_21482_, _20702_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53879_ (_21483_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53880_ (_21484_, _21483_, _21482_);
  and _53881_ (_21485_, _21484_, _22849_);
  nor _53882_ (_21486_, _21485_, _21481_);
  nor _53883_ (_21487_, _21486_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _53884_ (_21488_, _07572_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53885_ (_21489_, _21488_, _21471_);
  and _53886_ (_21490_, _21489_, _20681_);
  and _53887_ (_21491_, _08039_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53888_ (_21492_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _53889_ (_21493_, _21492_, _22849_);
  nor _53890_ (_21494_, _21493_, _21491_);
  and _53891_ (_21495_, _21494_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _53892_ (_21496_, _21495_, _21490_);
  not _53893_ (_21497_, _21496_);
  nor _53894_ (_21498_, _21497_, _21487_);
  nor _53895_ (_21499_, _21498_, _22841_);
  not _53896_ (_21500_, _21499_);
  nor _53897_ (_21501_, \oc8051_symbolic_cxrom1.regvalid [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _53898_ (_21502_, _21501_);
  nor _53899_ (_21503_, _21461_, _22849_);
  and _53900_ (_21504_, _21503_, _21502_);
  and _53901_ (_21505_, _08225_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53902_ (_21506_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53903_ (_21507_, _21506_, _21505_);
  and _53904_ (_21508_, _21507_, _22849_);
  nor _53905_ (_21509_, _21508_, _21504_);
  nor _53906_ (_21510_, _21509_, _20672_);
  and _53907_ (_21511_, _20696_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _53908_ (_21512_, _20712_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53909_ (_21513_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53910_ (_21514_, _21513_, _21512_);
  and _53911_ (_21515_, _21514_, _21511_);
  nor _53912_ (_21516_, \oc8051_symbolic_cxrom1.regvalid [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53913_ (_21517_, _21516_, _21450_);
  and _53914_ (_21518_, _20681_, _22841_);
  and _53915_ (_21519_, _21518_, _21517_);
  nor _53916_ (_21520_, _21519_, _21515_);
  not _53917_ (_21521_, _21520_);
  nor _53918_ (_21522_, _21521_, _21510_);
  and _53919_ (_21523_, _21522_, _21500_);
  and _53920_ (_21524_, _21489_, _20682_);
  nor _53921_ (_21525_, _21524_, _22841_);
  nor _53922_ (_21526_, _21486_, _22845_);
  nor _53923_ (_21527_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _53924_ (_21528_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _53925_ (_21529_, _07621_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53926_ (_21530_, _21529_, _21528_);
  and _53927_ (_21531_, _21530_, _21527_);
  nor _53928_ (_21532_, _21531_, _21526_);
  and _53929_ (_21533_, _21532_, _21525_);
  nor _53930_ (_21534_, _21509_, _22845_);
  nor _53931_ (_21535_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _53932_ (_21536_, _07665_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53933_ (_21537_, _21536_, _21535_);
  and _53934_ (_21538_, _21537_, _21527_);
  and _53935_ (_21539_, _21517_, _20682_);
  or _53936_ (_21540_, _21539_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _53937_ (_21541_, _21540_, _21538_);
  nor _53938_ (_21542_, _21541_, _21534_);
  nor _53939_ (_21543_, _21542_, _21533_);
  not _53940_ (_21544_, _22770_);
  nor _53941_ (_21545_, _21544_, first_instr);
  nand _53942_ (_21546_, _21545_, _21543_);
  nor _53943_ (_21547_, _21546_, _21523_);
  nand _53944_ (_21548_, _21547_, _21477_);
  nor _53945_ (_21549_, _21548_, _20736_);
  and _53946_ (_21550_, _21549_, _21427_);
  nor _53947_ (_21551_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53948_ (_21552_, _08575_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53949_ (_21553_, _21552_, _21551_);
  and _53950_ (_21554_, _21553_, _21527_);
  nor _53951_ (_21555_, _21554_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53952_ (_21556_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53953_ (_21557_, _09098_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53954_ (_21558_, _21557_, _21556_);
  and _53955_ (_21559_, _21558_, _20682_);
  not _53956_ (_21560_, _21559_);
  nor _53957_ (_21561_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53958_ (_21562_, _08830_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53959_ (_21563_, _21562_, _21561_);
  and _53960_ (_21564_, _21563_, _20681_);
  nor _53961_ (_21565_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53962_ (_21566_, _09352_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53963_ (_21567_, _21566_, _21565_);
  and _53964_ (_21568_, _21567_, _20656_);
  nor _53965_ (_21569_, _21568_, _21564_);
  and _53966_ (_21570_, _21569_, _21560_);
  and _53967_ (_21571_, _21570_, _21555_);
  nor _53968_ (_21572_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53969_ (_21573_, _09586_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53970_ (_21574_, _21573_, _21572_);
  and _53971_ (_21575_, _21574_, _21527_);
  nor _53972_ (_21576_, _21575_, _22854_);
  nor _53973_ (_21577_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53974_ (_21578_, _10084_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53975_ (_21579_, _21578_, _21577_);
  and _53976_ (_21580_, _21579_, _20682_);
  not _53977_ (_21581_, _21580_);
  nor _53978_ (_21582_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53979_ (_21583_, _09819_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53980_ (_21584_, _21583_, _21582_);
  and _53981_ (_21585_, _21584_, _20681_);
  nor _53982_ (_21586_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53983_ (_21587_, _10388_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53984_ (_21588_, _21587_, _21586_);
  and _53985_ (_21589_, _21588_, _20656_);
  nor _53986_ (_21590_, _21589_, _21585_);
  and _53987_ (_21591_, _21590_, _21581_);
  and _53988_ (_21592_, _21591_, _21576_);
  nor _53989_ (_21593_, _21592_, _21571_);
  and _53990_ (_21594_, _21593_, _21543_);
  nor _53991_ (_21595_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53992_ (_21596_, _09333_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53993_ (_21597_, _21596_, _21595_);
  and _53994_ (_21598_, _21597_, _20656_);
  nor _53995_ (_21599_, _21598_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _53996_ (_21600_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _53997_ (_21601_, _08809_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _53998_ (_21602_, _21601_, _21600_);
  and _53999_ (_21603_, _21602_, _20681_);
  not _54000_ (_21604_, _21603_);
  nor _54001_ (_21605_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54002_ (_21606_, _09080_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54003_ (_21607_, _21606_, _21605_);
  and _54004_ (_21608_, _21607_, _20682_);
  nor _54005_ (_21609_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54006_ (_21610_, _08556_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54007_ (_21611_, _21610_, _21609_);
  and _54008_ (_21612_, _21611_, _21527_);
  nor _54009_ (_21613_, _21612_, _21608_);
  and _54010_ (_21614_, _21613_, _21604_);
  and _54011_ (_21615_, _21614_, _21599_);
  nor _54012_ (_21616_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54013_ (_21617_, _10369_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54014_ (_21618_, _21617_, _21616_);
  and _54015_ (_21619_, _21618_, _20656_);
  nor _54016_ (_21620_, _21619_, _22854_);
  nor _54017_ (_21621_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54018_ (_21622_, _09802_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54019_ (_21623_, _21622_, _21621_);
  and _54020_ (_21624_, _21623_, _20681_);
  not _54021_ (_21625_, _21624_);
  nor _54022_ (_21626_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54023_ (_21627_, _10069_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54024_ (_21628_, _21627_, _21626_);
  and _54025_ (_21629_, _21628_, _20682_);
  nor _54026_ (_21630_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54027_ (_21631_, _09570_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54028_ (_21632_, _21631_, _21630_);
  and _54029_ (_21633_, _21632_, _21527_);
  nor _54030_ (_21634_, _21633_, _21629_);
  and _54031_ (_21635_, _21634_, _21625_);
  and _54032_ (_21636_, _21635_, _21620_);
  nor _54033_ (_21637_, _21636_, _21615_);
  and _54034_ (_21638_, _21637_, _21543_);
  nor _54035_ (_21639_, _21638_, _21594_);
  nor _54036_ (_21640_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54037_ (_21641_, _08857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54038_ (_21642_, _21641_, _21640_);
  and _54039_ (_21643_, _21642_, _20681_);
  nor _54040_ (_21644_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54041_ (_21645_, _09128_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54042_ (_21646_, _21645_, _21644_);
  and _54043_ (_21647_, _21646_, _20682_);
  nor _54044_ (_21648_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54045_ (_21649_, _08602_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54046_ (_21650_, _21649_, _21648_);
  and _54047_ (_21651_, _21650_, _21527_);
  nor _54048_ (_21652_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54049_ (_21653_, _09389_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54050_ (_21654_, _21653_, _21652_);
  and _54051_ (_21655_, _21654_, _20656_);
  or _54052_ (_21656_, _21655_, _21651_);
  or _54053_ (_21657_, _21656_, _21647_);
  or _54054_ (_21658_, _21657_, _21643_);
  and _54055_ (_21659_, _21658_, _22854_);
  nor _54056_ (_21660_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54057_ (_21661_, _09849_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54058_ (_21662_, _21661_, _21660_);
  and _54059_ (_21663_, _21662_, _20681_);
  nor _54060_ (_21664_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54061_ (_21665_, _10118_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54062_ (_21666_, _21665_, _21664_);
  and _54063_ (_21667_, _21666_, _20682_);
  nor _54064_ (_21668_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54065_ (_21669_, _09613_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54066_ (_21670_, _21669_, _21668_);
  and _54067_ (_21671_, _21670_, _21527_);
  nor _54068_ (_21672_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54069_ (_21673_, _10426_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54070_ (_21674_, _21673_, _21672_);
  and _54071_ (_21675_, _21674_, _20656_);
  or _54072_ (_21676_, _21675_, _21671_);
  or _54073_ (_21677_, _21676_, _21667_);
  or _54074_ (_21678_, _21677_, _21663_);
  and _54075_ (_21679_, _21678_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _54076_ (_21680_, _21679_, _21659_);
  and _54077_ (_21681_, _21680_, _21543_);
  nor _54078_ (_21682_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54079_ (_21683_, _08844_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54080_ (_21684_, _21683_, _21682_);
  and _54081_ (_21685_, _21684_, _20681_);
  nor _54082_ (_21686_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54083_ (_21687_, _09113_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54084_ (_21688_, _21687_, _21686_);
  and _54085_ (_21689_, _21688_, _20682_);
  nor _54086_ (_21690_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54087_ (_21691_, _08589_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54088_ (_21692_, _21691_, _21690_);
  and _54089_ (_21693_, _21692_, _21527_);
  nor _54090_ (_21694_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54091_ (_21695_, _09371_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54092_ (_21696_, _21695_, _21694_);
  and _54093_ (_21697_, _21696_, _20656_);
  or _54094_ (_21698_, _21697_, _21693_);
  or _54095_ (_21699_, _21698_, _21689_);
  or _54096_ (_21700_, _21699_, _21685_);
  and _54097_ (_21701_, _21700_, _22854_);
  nor _54098_ (_21702_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54099_ (_21703_, _09834_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54100_ (_21704_, _21703_, _21702_);
  and _54101_ (_21705_, _21704_, _20681_);
  nor _54102_ (_21706_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54103_ (_21707_, _10102_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54104_ (_21708_, _21707_, _21706_);
  and _54105_ (_21709_, _21708_, _20682_);
  nor _54106_ (_21710_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54107_ (_21711_, _09598_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54108_ (_21712_, _21711_, _21710_);
  and _54109_ (_21713_, _21712_, _21527_);
  nor _54110_ (_21714_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54111_ (_21715_, _10410_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54112_ (_21716_, _21715_, _21714_);
  and _54113_ (_21717_, _21716_, _20656_);
  or _54114_ (_21718_, _21717_, _21713_);
  or _54115_ (_21719_, _21718_, _21709_);
  or _54116_ (_21720_, _21719_, _21705_);
  and _54117_ (_21721_, _21720_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _54118_ (_21722_, _21721_, _21701_);
  and _54119_ (_21723_, _21722_, _21543_);
  nor _54120_ (_21724_, _21723_, _21681_);
  and _54121_ (_21725_, _21724_, _21639_);
  nor _54122_ (_21726_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54123_ (_21727_, _08883_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54124_ (_21728_, _21727_, _21726_);
  and _54125_ (_21729_, _21728_, _20681_);
  nor _54126_ (_21730_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54127_ (_21731_, _09153_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54128_ (_21732_, _21731_, _21730_);
  and _54129_ (_21733_, _21732_, _20682_);
  nor _54130_ (_21734_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54131_ (_21735_, _08630_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54132_ (_21736_, _21735_, _21734_);
  and _54133_ (_21737_, _21736_, _21527_);
  nor _54134_ (_21738_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54135_ (_21739_, _09415_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54136_ (_21740_, _21739_, _21738_);
  and _54137_ (_21741_, _21740_, _20656_);
  or _54138_ (_21742_, _21741_, _21737_);
  or _54139_ (_21743_, _21742_, _21733_);
  or _54140_ (_21744_, _21743_, _21729_);
  and _54141_ (_21745_, _21744_, _22854_);
  nor _54142_ (_21746_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54143_ (_21747_, _09875_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54144_ (_21748_, _21747_, _21746_);
  and _54145_ (_21749_, _21748_, _20681_);
  nor _54146_ (_21750_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54147_ (_21751_, _10150_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54148_ (_21752_, _21751_, _21750_);
  and _54149_ (_21753_, _21752_, _20682_);
  nor _54150_ (_21754_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54151_ (_21755_, _09641_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54152_ (_21756_, _21755_, _21754_);
  and _54153_ (_21757_, _21756_, _21527_);
  nor _54154_ (_21758_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54155_ (_21759_, _10453_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54156_ (_21760_, _21759_, _21758_);
  and _54157_ (_21761_, _21760_, _20656_);
  or _54158_ (_21762_, _21761_, _21757_);
  or _54159_ (_21763_, _21762_, _21753_);
  or _54160_ (_21764_, _21763_, _21749_);
  and _54161_ (_21765_, _21764_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _54162_ (_21766_, _21765_, _21745_);
  and _54163_ (_21767_, _21766_, _21543_);
  nor _54164_ (_21768_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54165_ (_21769_, _08617_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54166_ (_21770_, _21769_, _21768_);
  and _54167_ (_21771_, _21770_, _21527_);
  nor _54168_ (_21772_, _21771_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _54169_ (_21773_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54170_ (_21774_, _09141_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54171_ (_21775_, _21774_, _21773_);
  and _54172_ (_21776_, _21775_, _20682_);
  not _54173_ (_21777_, _21776_);
  nor _54174_ (_21778_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54175_ (_21779_, _08870_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54176_ (_21780_, _21779_, _21778_);
  and _54177_ (_21781_, _21780_, _20681_);
  nor _54178_ (_21782_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54179_ (_21783_, _09402_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54180_ (_21784_, _21783_, _21782_);
  and _54181_ (_21785_, _21784_, _20656_);
  nor _54182_ (_21786_, _21785_, _21781_);
  and _54183_ (_21787_, _21786_, _21777_);
  and _54184_ (_21788_, _21787_, _21772_);
  nor _54185_ (_21789_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54186_ (_21790_, _09627_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54187_ (_21791_, _21790_, _21789_);
  and _54188_ (_21792_, _21791_, _21527_);
  nor _54189_ (_21793_, _21792_, _22854_);
  nor _54190_ (_21794_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54191_ (_21795_, _10135_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54192_ (_21796_, _21795_, _21794_);
  and _54193_ (_21797_, _21796_, _20682_);
  not _54194_ (_21798_, _21797_);
  nor _54195_ (_21799_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54196_ (_21800_, _09863_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54197_ (_21801_, _21800_, _21799_);
  and _54198_ (_21802_, _21801_, _20681_);
  nor _54199_ (_21803_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54200_ (_21804_, _10441_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54201_ (_21805_, _21804_, _21803_);
  and _54202_ (_21806_, _21805_, _20656_);
  nor _54203_ (_21807_, _21806_, _21802_);
  and _54204_ (_21808_, _21807_, _21798_);
  and _54205_ (_21809_, _21808_, _21793_);
  nor _54206_ (_21810_, _21809_, _21788_);
  and _54207_ (_21811_, _21810_, _21543_);
  nor _54208_ (_21812_, _21811_, _21767_);
  nor _54209_ (_21813_, \oc8051_symbolic_cxrom1.regarray[0] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54210_ (_21814_, _07675_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54211_ (_21815_, _21814_, _21813_);
  and _54212_ (_21816_, _21815_, _21527_);
  nor _54213_ (_21817_, _21816_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _54214_ (_21818_, \oc8051_symbolic_cxrom1.regarray[4] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54215_ (_21819_, _07689_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54216_ (_21821_, _21819_, _21818_);
  and _54217_ (_21822_, _21821_, _20682_);
  not _54218_ (_21823_, _21822_);
  nor _54219_ (_21824_, \oc8051_symbolic_cxrom1.regarray[2] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54220_ (_21825_, _07696_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54221_ (_21826_, _21825_, _21824_);
  and _54222_ (_21827_, _21826_, _20681_);
  nor _54223_ (_21828_, \oc8051_symbolic_cxrom1.regarray[6] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54224_ (_21829_, _07682_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54225_ (_21830_, _21829_, _21828_);
  and _54226_ (_21831_, _21830_, _20656_);
  nor _54227_ (_21832_, _21831_, _21827_);
  and _54228_ (_21833_, _21832_, _21823_);
  and _54229_ (_21834_, _21833_, _21817_);
  nor _54230_ (_21835_, \oc8051_symbolic_cxrom1.regarray[8] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54231_ (_21836_, _07709_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54232_ (_21837_, _21836_, _21835_);
  and _54233_ (_21838_, _21837_, _21527_);
  nor _54234_ (_21839_, _21838_, _22854_);
  nor _54235_ (_21840_, \oc8051_symbolic_cxrom1.regarray[12] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54236_ (_21841_, _07717_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54237_ (_21842_, _21841_, _21840_);
  and _54238_ (_21843_, _21842_, _20682_);
  not _54239_ (_21844_, _21843_);
  nor _54240_ (_21845_, \oc8051_symbolic_cxrom1.regarray[10] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54241_ (_21846_, _07731_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54242_ (_21847_, _21846_, _21845_);
  and _54243_ (_21848_, _21847_, _20681_);
  nor _54244_ (_21849_, \oc8051_symbolic_cxrom1.regarray[14] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54245_ (_21850_, _07723_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54246_ (_21851_, _21850_, _21849_);
  and _54247_ (_21852_, _21851_, _20656_);
  nor _54248_ (_21853_, _21852_, _21848_);
  and _54249_ (_21854_, _21853_, _21844_);
  and _54250_ (_21855_, _21854_, _21839_);
  nor _54251_ (_21856_, _21855_, _21834_);
  and _54252_ (_21857_, _21856_, _21543_);
  nor _54253_ (_21858_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54254_ (_21859_, _08646_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54255_ (_21860_, _21859_, _21858_);
  and _54256_ (_21861_, _21860_, _21527_);
  nor _54257_ (_21862_, _21861_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _54258_ (_21863_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54259_ (_21864_, _09166_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54260_ (_21865_, _21864_, _21863_);
  and _54261_ (_21866_, _21865_, _20682_);
  not _54262_ (_21867_, _21866_);
  nor _54263_ (_21868_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54264_ (_21869_, _08898_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54265_ (_21870_, _21869_, _21868_);
  and _54266_ (_21871_, _21870_, _20681_);
  nor _54267_ (_21872_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54268_ (_21873_, _09428_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54269_ (_21874_, _21873_, _21872_);
  and _54270_ (_21875_, _21874_, _20656_);
  nor _54271_ (_21876_, _21875_, _21871_);
  and _54272_ (_21877_, _21876_, _21867_);
  and _54273_ (_21878_, _21877_, _21862_);
  nor _54274_ (_21879_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54275_ (_21880_, _09654_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54276_ (_21881_, _21880_, _21879_);
  and _54277_ (_21882_, _21881_, _21527_);
  nor _54278_ (_21883_, _21882_, _22854_);
  nor _54279_ (_21884_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54280_ (_21885_, _10166_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54281_ (_21886_, _21885_, _21884_);
  and _54282_ (_21887_, _21886_, _20682_);
  not _54283_ (_21888_, _21887_);
  nor _54284_ (_21889_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54285_ (_21890_, _09888_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54286_ (_21891_, _21890_, _21889_);
  and _54287_ (_21892_, _21891_, _20681_);
  nor _54288_ (_21893_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54289_ (_21894_, _10467_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54290_ (_21895_, _21894_, _21893_);
  and _54291_ (_21896_, _21895_, _20656_);
  nor _54292_ (_21897_, _21896_, _21892_);
  and _54293_ (_21898_, _21897_, _21888_);
  and _54294_ (_21899_, _21898_, _21883_);
  nor _54295_ (_21900_, _21899_, _21878_);
  not _54296_ (_21901_, _21900_);
  and _54297_ (_21902_, _21901_, _21857_);
  and _54298_ (_21903_, _21902_, _21812_);
  and _54299_ (_21904_, _21903_, _21725_);
  and _54300_ (_21905_, _21904_, _21550_);
  and _54301_ (_21906_, _21905_, _21270_);
  not _54302_ (_21907_, _21857_);
  and _54303_ (_21908_, _21900_, _21543_);
  nand _54304_ (_21909_, _21811_, _21766_);
  and _54305_ (_21910_, _21723_, _21594_);
  nor _54306_ (_21911_, _21910_, _21680_);
  nor _54307_ (_21912_, _21911_, _21909_);
  not _54308_ (_21913_, _21638_);
  and _54309_ (_21914_, _21724_, _21913_);
  and _54310_ (_21915_, _21914_, _21594_);
  not _54311_ (_21916_, _21637_);
  not _54312_ (_21917_, _21593_);
  not _54313_ (_21918_, _21680_);
  and _54314_ (_21919_, _21723_, _21918_);
  and _54315_ (_21920_, _21919_, _21917_);
  and _54316_ (_21921_, _21920_, _21916_);
  or _54317_ (_21922_, _21921_, _21915_);
  or _54318_ (_21923_, _21922_, _21912_);
  and _54319_ (_21924_, _21923_, _21908_);
  and _54320_ (_21925_, _21901_, _21767_);
  and _54321_ (_21926_, _21925_, _21920_);
  not _54322_ (_21927_, _21767_);
  and _54323_ (_21928_, _21920_, _21638_);
  and _54324_ (_21929_, _21928_, _21927_);
  or _54325_ (_21930_, _21929_, _21926_);
  or _54326_ (_21931_, _21930_, _21924_);
  and _54327_ (_21932_, _21931_, _21907_);
  and _54328_ (_21933_, _21915_, _21927_);
  not _54329_ (_21934_, _21908_);
  nor _54330_ (_21935_, _21934_, _21766_);
  and _54331_ (_21936_, _21935_, _21914_);
  and _54332_ (_21937_, _21908_, _21766_);
  and _54333_ (_21938_, _21937_, _21928_);
  or _54334_ (_21939_, _21938_, _21936_);
  or _54335_ (_21940_, _21939_, _21933_);
  and _54336_ (_21941_, _21940_, _21857_);
  not _54337_ (_21942_, _21810_);
  and _54338_ (_21943_, _21908_, _21942_);
  and _54339_ (_21944_, _21943_, _21928_);
  and _54340_ (_21945_, _21811_, _21927_);
  and _54341_ (_21946_, _21945_, _21920_);
  and _54342_ (_21947_, _21767_, _21914_);
  and _54343_ (_21948_, _21942_, _21681_);
  not _54344_ (_21949_, _21811_);
  and _54345_ (_21950_, _21910_, _21949_);
  or _54346_ (_21951_, _21950_, _21948_);
  or _54347_ (_21952_, _21951_, _21947_);
  or _54348_ (_21953_, _21952_, _21946_);
  and _54349_ (_21954_, _21953_, _21902_);
  or _54350_ (_21955_, _21954_, _21944_);
  or _54351_ (_21956_, _21955_, _21941_);
  or _54352_ (_21957_, _21956_, _21932_);
  nor _54353_ (_21958_, _20782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _54354_ (_21959_, _20782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or _54355_ (_21960_, _21959_, _21958_);
  nor _54356_ (_21961_, _20786_, _22827_);
  and _54357_ (_21962_, _20786_, _22827_);
  or _54358_ (_21963_, _21962_, _21961_);
  or _54359_ (_21964_, _21963_, _21960_);
  and _54360_ (_21965_, _20670_, _22837_);
  nor _54361_ (_21966_, _20670_, _22837_);
  or _54362_ (_21967_, _21966_, _21965_);
  or _54363_ (_21968_, _21967_, _21157_);
  or _54364_ (_21969_, _21968_, _21964_);
  or _54365_ (_21970_, _20796_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _54366_ (_21971_, _20796_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _54367_ (_21972_, _21971_, _21970_);
  or _54368_ (_21973_, _21197_, _21182_);
  and _54369_ (_21974_, _20817_, _22802_);
  nor _54370_ (_21975_, _20683_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _54371_ (_21976_, _20683_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _54372_ (_21977_, _21976_, _21975_);
  nor _54373_ (_21978_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _54374_ (_21979_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _54375_ (_21980_, _21979_, _21978_);
  not _54376_ (_21981_, _21980_);
  and _54377_ (_21982_, _21981_, _20657_);
  or _54378_ (_21983_, _21982_, _21977_);
  and _54379_ (_21984_, _20676_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _54380_ (_21985_, _20676_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _54381_ (_21986_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _54382_ (_21987_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _54383_ (_21988_, _21987_, _21986_);
  nand _54384_ (_21989_, _21988_, _21233_);
  nor _54385_ (_21990_, _21981_, _20657_);
  or _54386_ (_21991_, _21990_, _21989_);
  or _54387_ (_21992_, _21991_, _21985_);
  or _54388_ (_21993_, _21992_, _21984_);
  or _54389_ (_21994_, _21993_, _21983_);
  nor _54390_ (_21995_, _20817_, _22802_);
  or _54391_ (_21996_, _21995_, _21994_);
  or _54392_ (_21997_, _21996_, _21974_);
  or _54393_ (_21998_, _20806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _54394_ (_21999_, _20806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _54395_ (_22000_, _21999_, _21998_);
  nor _54396_ (_22001_, _20862_, _22798_);
  and _54397_ (_22002_, _20862_, _22798_);
  or _54398_ (_22003_, _22002_, _22001_);
  nor _54399_ (_22004_, _20811_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _54400_ (_22005_, _20811_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or _54401_ (_22006_, _22005_, _22004_);
  or _54402_ (_22007_, _22006_, _22003_);
  or _54403_ (_22008_, _22007_, _22000_);
  or _54404_ (_22009_, _22008_, _21997_);
  or _54405_ (_22010_, _22009_, _21973_);
  or _54406_ (_22011_, _22010_, _21972_);
  or _54407_ (_22012_, _22011_, _21969_);
  and _54408_ (_22013_, _22012_, _21957_);
  and _54409_ (_22014_, _21638_, _21594_);
  and _54410_ (_22015_, _22014_, _21724_);
  and _54411_ (_22016_, _21921_, _21812_);
  or _54412_ (_22017_, _22016_, _22015_);
  nor _54413_ (_22018_, _21766_, _21637_);
  nand _54414_ (_22019_, _22018_, _21723_);
  nand _54415_ (_22020_, _21812_, _21639_);
  and _54416_ (_22021_, _22020_, _22019_);
  nor _54417_ (_22022_, _22021_, _21857_);
  or _54418_ (_22023_, _22022_, _22017_);
  and _54419_ (_22024_, _22023_, _21934_);
  and _54420_ (_22025_, _21926_, _21949_);
  or _54421_ (_22026_, _21919_, _21767_);
  or _54422_ (_22027_, _21680_, _21916_);
  and _54423_ (_22028_, _22027_, _21908_);
  and _54424_ (_22029_, _22028_, _22026_);
  or _54425_ (_22030_, _22029_, _22025_);
  and _54426_ (_22031_, _22030_, _21857_);
  nor _54427_ (_22032_, _21856_, _21766_);
  not _54428_ (_22033_, _21856_);
  or _54429_ (_22034_, _21945_, _22033_);
  and _54430_ (_22035_, _22034_, _21901_);
  or _54431_ (_22036_, _22035_, _22032_);
  and _54432_ (_22037_, _22036_, _21681_);
  nor _54433_ (_22038_, _21908_, _21857_);
  or _54434_ (_22039_, _21942_, _21767_);
  nor _54435_ (_22040_, _22039_, _21681_);
  or _54436_ (_22041_, _22040_, _22038_);
  and _54437_ (_22042_, _22041_, _21910_);
  and _54438_ (_22043_, _21948_, _21908_);
  nor _54439_ (_22044_, _22027_, _22033_);
  and _54440_ (_22045_, _22044_, _21594_);
  or _54441_ (_22046_, _22045_, _21950_);
  and _54442_ (_22047_, _22046_, _21908_);
  or _54443_ (_22048_, _22047_, _22043_);
  or _54444_ (_22049_, _22048_, _22042_);
  or _54445_ (_22050_, _22049_, _22037_);
  or _54446_ (_22051_, _22050_, _22031_);
  or _54447_ (_22052_, _22051_, _22024_);
  and _54448_ (_22053_, _20780_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _54449_ (_22054_, _22053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and _54450_ (_22055_, _22054_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54451_ (_22056_, _22053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54452_ (_22057_, _22056_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or _54453_ (_22058_, _22057_, _22055_);
  and _54454_ (_22059_, _22058_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _54455_ (_22060_, _20791_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _54456_ (_22061_, _22890_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54457_ (_22062_, _22061_, _22060_);
  nor _54458_ (_22063_, _22062_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _54459_ (_22064_, _22062_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not _54460_ (_22065_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _54461_ (_22066_, _20657_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54462_ (_22067_, _22066_, _20660_);
  and _54463_ (_22068_, _22067_, _20664_);
  and _54464_ (_22069_, _22068_, _22065_);
  nor _54465_ (_22070_, _22068_, _22065_);
  or _54466_ (_22071_, _22070_, _22069_);
  and _54467_ (_22072_, _22071_, _22827_);
  or _54468_ (_22073_, _22072_, _22064_);
  or _54469_ (_22074_, _22073_, _22063_);
  and _54470_ (_22075_, _22067_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _54471_ (_22076_, _22075_, _22882_);
  nor _54472_ (_22077_, _22075_, _22882_);
  nor _54473_ (_22078_, _22077_, _22076_);
  and _54474_ (_22079_, _22078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _54475_ (_22080_, _20678_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _54476_ (_22081_, _20678_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _54477_ (_22082_, _22081_, _22080_);
  and _54478_ (_22083_, _20808_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _54479_ (_22084_, _22083_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _54480_ (_22085_, _22084_, _22067_);
  nor _54481_ (_22086_, _22085_, _22806_);
  and _54482_ (_22087_, _22085_, _22806_);
  or _54483_ (_22088_, _22087_, _22086_);
  or _54484_ (_22089_, _22088_, _22082_);
  nor _54485_ (_22090_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _54486_ (_22091_, _22090_, _22083_);
  nor _54487_ (_22092_, _22091_, _20816_);
  and _54488_ (_22093_, _22092_, _22802_);
  nor _54489_ (_22094_, _20685_, _22783_);
  and _54490_ (_22095_, _20685_, _22783_);
  or _54491_ (_22096_, _22095_, _22094_);
  nand _54492_ (_22097_, _21988_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _54493_ (_22098_, _21988_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54494_ (_22099_, _22098_, _22097_);
  nor _54495_ (_22100_, _22066_, _21981_);
  and _54496_ (_22101_, _22066_, _21981_);
  or _54497_ (_22102_, _22101_, _21233_);
  or _54498_ (_22103_, _22102_, _22100_);
  or _54499_ (_22104_, _22103_, _22099_);
  or _54500_ (_22105_, _22104_, _22096_);
  or _54501_ (_22106_, _22105_, _22093_);
  or _54502_ (_22107_, _22106_, _22089_);
  or _54503_ (_22108_, _22864_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand _54504_ (_22109_, _20862_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54505_ (_22110_, _22109_, _22108_);
  and _54506_ (_22111_, _22110_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _54507_ (_22112_, _22110_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or _54508_ (_22113_, _22112_, _22111_);
  or _54509_ (_22114_, _22113_, _22107_);
  or _54510_ (_22115_, _22114_, _22079_);
  nor _54511_ (_22116_, _22071_, _22827_);
  nor _54512_ (_22117_, _22078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  or _54513_ (_22118_, _22117_, _22116_);
  or _54514_ (_22119_, _22118_, _22115_);
  or _54515_ (_22120_, _22119_, _22074_);
  or _54516_ (_22121_, _22120_, _22059_);
  nor _54517_ (_22122_, _22057_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _54518_ (_22123_, _22122_, _21152_);
  nor _54519_ (_22124_, _22123_, _22055_);
  or _54520_ (_22125_, _20782_, _22841_);
  or _54521_ (_22126_, _22897_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _54522_ (_22127_, _22126_, _22125_);
  and _54523_ (_22128_, _22127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _54524_ (_22129_, _22067_, _20662_);
  and _54525_ (_22130_, _22129_, _22886_);
  nor _54526_ (_22131_, _22129_, _22886_);
  or _54527_ (_22132_, _22131_, _22130_);
  nor _54528_ (_22133_, _22132_, _22819_);
  and _54529_ (_22134_, _22132_, _22819_);
  nor _54530_ (_22135_, _22067_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _54531_ (_22136_, _22135_, _22075_);
  and _54532_ (_22137_, _22136_, _22810_);
  nor _54533_ (_22138_, _22136_, _22810_);
  nor _54534_ (_22139_, _22092_, _22802_);
  or _54535_ (_22140_, _22139_, _22138_);
  or _54536_ (_22141_, _22140_, _22137_);
  or _54537_ (_22142_, _22141_, _22134_);
  or _54538_ (_22143_, _22142_, _22133_);
  or _54539_ (_22144_, _22143_, _22128_);
  nor _54540_ (_22145_, _22127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _54541_ (_22146_, _22055_, _21153_);
  or _54542_ (_22147_, _22146_, _22145_);
  or _54543_ (_22148_, _22147_, _22144_);
  or _54544_ (_22149_, _22148_, _22124_);
  or _54545_ (_22150_, _22149_, _22121_);
  and _54546_ (_22151_, _22150_, _22052_);
  and _54547_ (_22152_, _21945_, _21725_);
  and _54548_ (_22153_, _21929_, _21942_);
  or _54549_ (_22154_, _22153_, _22152_);
  and _54550_ (_22155_, _22154_, _21902_);
  and _54551_ (_22156_, _21938_, _21811_);
  and _54552_ (_22157_, _21909_, _21908_);
  and _54553_ (_22158_, _22157_, _22015_);
  or _54554_ (_22159_, _22158_, _22156_);
  and _54555_ (_22160_, _22159_, _21907_);
  or _54556_ (_22161_, _22160_, _22155_);
  and _54557_ (_22162_, _21432_, _20660_);
  and _54558_ (_22163_, _22162_, _20663_);
  and _54559_ (_22164_, _22163_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _54560_ (_22165_, _22164_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _54561_ (_22166_, _22165_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _54562_ (_22167_, _22166_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _54563_ (_22168_, _22166_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _54564_ (_22169_, _22168_, _22167_);
  nor _54565_ (_22170_, _22169_, _22837_);
  nor _54566_ (_22171_, _22165_, _22897_);
  and _54567_ (_22172_, _22165_, _22897_);
  nor _54568_ (_22173_, _22172_, _22171_);
  nor _54569_ (_22174_, _22173_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _54570_ (_22175_, _22169_, _22837_);
  or _54571_ (_22176_, _22175_, _22174_);
  or _54572_ (_22177_, _22176_, _22170_);
  nor _54573_ (_22178_, _22164_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _54574_ (_22179_, _22178_, _22165_);
  and _54575_ (_22180_, _22179_, _22827_);
  nor _54576_ (_22181_, _22179_, _22827_);
  or _54577_ (_22182_, _22181_, _22180_);
  nor _54578_ (_22183_, _22167_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and _54579_ (_22184_, _22167_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _54580_ (_22185_, _22184_, _22183_);
  nor _54581_ (_22186_, _22185_, _14710_);
  or _54582_ (_22187_, _22186_, _22182_);
  and _54583_ (_22188_, _22162_, _20662_);
  nor _54584_ (_22189_, _22188_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _54585_ (_22190_, _22189_, _22163_);
  and _54586_ (_22191_, _22190_, _22819_);
  and _54587_ (_22192_, _22185_, _14710_);
  or _54588_ (_22193_, _22192_, _22191_);
  and _54589_ (_22194_, _22173_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _54590_ (_22195_, _21432_, _20659_);
  and _54591_ (_22196_, _21432_, _20658_);
  nor _54592_ (_22197_, _22196_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _54593_ (_22198_, _22197_, _22195_);
  and _54594_ (_22199_, _22198_, _22802_);
  nor _54595_ (_22200_, _22163_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _54596_ (_22201_, _22200_, _22164_);
  nor _54597_ (_22202_, _22201_, _22823_);
  and _54598_ (_22203_, _22162_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _54599_ (_22204_, _22162_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _54600_ (_22205_, _22204_, _22203_);
  nor _54601_ (_22206_, _22205_, _22810_);
  and _54602_ (_22207_, _22205_, _22810_);
  or _54603_ (_22208_, _22207_, _22206_);
  or _54604_ (_22209_, _22208_, _22202_);
  or _54605_ (_22210_, _22209_, _22199_);
  or _54606_ (_22211_, _22210_, _22194_);
  and _54607_ (_22212_, _22201_, _22823_);
  nor _54608_ (_22213_, _22203_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _54609_ (_22214_, _22213_, _22188_);
  nor _54610_ (_22215_, _22214_, _22814_);
  and _54611_ (_22216_, _22214_, _22814_);
  or _54612_ (_22217_, _22216_, _22215_);
  nor _54613_ (_22218_, _22195_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _54614_ (_22219_, _22218_, _22162_);
  and _54615_ (_22220_, _22219_, _22806_);
  nor _54616_ (_22221_, _22190_, _22819_);
  or _54617_ (_22222_, _22221_, _22220_);
  or _54618_ (_22223_, _22222_, _22217_);
  or _54619_ (_22224_, _21980_, _21432_);
  nand _54620_ (_22225_, _21980_, _21432_);
  and _54621_ (_22226_, _22225_, _22224_);
  nand _54622_ (_22227_, _21430_, _22783_);
  nand _54623_ (_22228_, _22227_, _22099_);
  or _54624_ (_22229_, _22228_, _22226_);
  and _54625_ (_22230_, _21432_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _54626_ (_22231_, _22230_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _54627_ (_22232_, _22231_, _22196_);
  and _54628_ (_22233_, _22232_, _22798_);
  nor _54629_ (_22234_, _22198_, _22802_);
  or _54630_ (_22235_, _22234_, _22233_);
  nor _54631_ (_22236_, _22232_, _22798_);
  nor _54632_ (_22237_, _21430_, _22783_);
  or _54633_ (_22238_, _22237_, _21233_);
  or _54634_ (_22239_, _22238_, _22236_);
  or _54635_ (_22240_, _22239_, _22235_);
  nor _54636_ (_22241_, _22219_, _22806_);
  or _54637_ (_22242_, _21434_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _54638_ (_22243_, _21434_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _54639_ (_22244_, _22243_, _22242_);
  or _54640_ (_22245_, _22244_, _22241_);
  or _54641_ (_22246_, _22245_, _22240_);
  or _54642_ (_22247_, _22246_, _22229_);
  or _54643_ (_22248_, _22247_, _22223_);
  or _54644_ (_22249_, _22248_, _22212_);
  or _54645_ (_22250_, _22249_, _22211_);
  or _54646_ (_22251_, _22250_, _22193_);
  or _54647_ (_22252_, _22251_, _22187_);
  or _54648_ (_22253_, _22252_, _22177_);
  and _54649_ (_22254_, _22253_, _22161_);
  or _54650_ (_22255_, _22254_, _22151_);
  or _54651_ (_22256_, _22255_, _22013_);
  and _54652_ (_22257_, _22256_, _21550_);
  or _54653_ (_22258_, _20984_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _54654_ (_22259_, _20984_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _54655_ (_22260_, _22259_, _22258_);
  or _54656_ (_22261_, _20900_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _54657_ (_22262_, _20900_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _54658_ (_22263_, _22262_, _22261_);
  or _54659_ (_22264_, _22263_, _22260_);
  or _54660_ (_22265_, _21066_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _54661_ (_22266_, _21066_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _54662_ (_22267_, _22266_, _22265_);
  and _54663_ (_22268_, _21105_, _22772_);
  nor _54664_ (_22269_, _21027_, _22783_);
  or _54665_ (_22270_, _22269_, _22268_);
  or _54666_ (_22271_, _22270_, _22267_);
  and _54667_ (_22272_, _21767_, _22810_);
  nor _54668_ (_22273_, _21767_, _22810_);
  or _54669_ (_22274_, _22273_, _22272_);
  nor _54670_ (_22275_, _21908_, _22814_);
  and _54671_ (_22276_, _21908_, _22814_);
  or _54672_ (_22277_, _22276_, _22275_);
  or _54673_ (_22278_, _22277_, _22274_);
  nor _54674_ (_22279_, _21857_, _22819_);
  and _54675_ (_22280_, _21857_, _22819_);
  or _54676_ (_22281_, _22280_, _22279_);
  or _54677_ (_22282_, _22281_, _21182_);
  or _54678_ (_22283_, _22282_, _22278_);
  nor _54679_ (_22284_, _21105_, _22772_);
  or _54680_ (_22285_, _22284_, _21969_);
  or _54681_ (_22286_, _22285_, _22283_);
  or _54682_ (_22287_, _22286_, _22271_);
  or _54683_ (_22288_, _20775_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand _54684_ (_22289_, _20775_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _54685_ (_22290_, _22289_, _22288_);
  and _54686_ (_22291_, _20855_, _22802_);
  or _54687_ (_22292_, _22291_, _22290_);
  nor _54688_ (_22293_, _20855_, _22802_);
  and _54689_ (_22294_, _20942_, _22794_);
  or _54690_ (_22295_, _22294_, _22293_);
  nor _54691_ (_22296_, _20942_, _22794_);
  and _54692_ (_22297_, _21027_, _22783_);
  or _54693_ (_22298_, _22297_, _22296_);
  or _54694_ (_22299_, _22298_, _22295_);
  or _54695_ (_22300_, _22299_, _22292_);
  or _54696_ (_22301_, _22300_, _22287_);
  or _54697_ (_22302_, _22301_, _22264_);
  and _54698_ (_22303_, _21638_, _21917_);
  and _54699_ (_22304_, _22303_, _21724_);
  and _54700_ (_22305_, _22304_, _22302_);
  and _54701_ (_22306_, _21886_, _20681_);
  or _54702_ (_22307_, _22306_, _20676_);
  and _54703_ (_22308_, _21881_, _20656_);
  and _54704_ (_22309_, _21891_, _21527_);
  and _54705_ (_22310_, _21895_, _20682_);
  or _54706_ (_22311_, _22310_, _22309_);
  or _54707_ (_22312_, _22311_, _22308_);
  or _54708_ (_22313_, _22312_, _22307_);
  and _54709_ (_22314_, _21865_, _20681_);
  or _54710_ (_22315_, _22314_, _20946_);
  and _54711_ (_22316_, _21860_, _20656_);
  and _54712_ (_22317_, _21870_, _21527_);
  and _54713_ (_22318_, _21874_, _20682_);
  or _54714_ (_22319_, _22318_, _22317_);
  or _54715_ (_22320_, _22319_, _22316_);
  or _54716_ (_22321_, _22320_, _22315_);
  nand _54717_ (_22322_, _22321_, _22313_);
  nor _54718_ (_22323_, _22322_, _21523_);
  nand _54719_ (_22324_, _22323_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or _54720_ (_22325_, _22323_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _54721_ (_22326_, _22325_, _22324_);
  not _54722_ (_22327_, _21523_);
  and _54723_ (_22328_, _21842_, _20681_);
  and _54724_ (_22329_, _21851_, _20682_);
  nor _54725_ (_22330_, _22329_, _22328_);
  and _54726_ (_22331_, _21837_, _20656_);
  and _54727_ (_22332_, _21847_, _21527_);
  nor _54728_ (_22333_, _22332_, _22331_);
  and _54729_ (_22334_, _22333_, _22330_);
  and _54730_ (_22335_, _22334_, _20946_);
  and _54731_ (_22336_, _21830_, _20682_);
  and _54732_ (_22337_, _21815_, _20656_);
  and _54733_ (_22338_, _21821_, _20681_);
  or _54734_ (_22339_, _22338_, _22337_);
  nor _54735_ (_22340_, _22339_, _22336_);
  and _54736_ (_22341_, _21826_, _21527_);
  nor _54737_ (_22342_, _22341_, _20946_);
  and _54738_ (_22343_, _22342_, _22340_);
  nor _54739_ (_22344_, _22343_, _22335_);
  and _54740_ (_22345_, _22344_, _22327_);
  nor _54741_ (_22346_, _22345_, _22806_);
  and _54742_ (_22347_, _22345_, _22806_);
  or _54743_ (_22348_, _22347_, _22346_);
  or _54744_ (_22349_, _22348_, _22326_);
  and _54745_ (_22350_, _21732_, _20681_);
  or _54746_ (_22351_, _22350_, _20946_);
  and _54747_ (_22352_, _21736_, _20656_);
  and _54748_ (_22353_, _21728_, _21527_);
  and _54749_ (_22354_, _21740_, _20682_);
  or _54750_ (_22355_, _22354_, _22353_);
  or _54751_ (_22356_, _22355_, _22352_);
  or _54752_ (_22357_, _22356_, _22351_);
  and _54753_ (_22358_, _21752_, _20681_);
  or _54754_ (_22359_, _22358_, _20676_);
  and _54755_ (_22360_, _21756_, _20656_);
  and _54756_ (_22361_, _21748_, _21527_);
  and _54757_ (_22362_, _21760_, _20682_);
  or _54758_ (_22363_, _22362_, _22361_);
  or _54759_ (_22364_, _22363_, _22360_);
  or _54760_ (_22365_, _22364_, _22359_);
  nand _54761_ (_22366_, _22365_, _22357_);
  nor _54762_ (_22367_, _22366_, _21523_);
  nand _54763_ (_22368_, _22367_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or _54764_ (_22369_, _22367_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _54765_ (_22370_, _22369_, _22368_);
  and _54766_ (_22371_, _21775_, _20681_);
  and _54767_ (_22372_, _21784_, _20682_);
  and _54768_ (_22373_, _21770_, _20656_);
  or _54769_ (_22374_, _22373_, _22372_);
  or _54770_ (_22375_, _22374_, _22371_);
  and _54771_ (_22376_, _21780_, _21527_);
  or _54772_ (_22377_, _22376_, _20946_);
  or _54773_ (_22378_, _22377_, _22375_);
  and _54774_ (_22379_, _21796_, _20681_);
  or _54775_ (_22380_, _22379_, _20676_);
  and _54776_ (_22381_, _21791_, _20656_);
  and _54777_ (_22382_, _21801_, _21527_);
  and _54778_ (_22383_, _21805_, _20682_);
  or _54779_ (_22384_, _22383_, _22382_);
  or _54780_ (_22385_, _22384_, _22381_);
  or _54781_ (_22386_, _22385_, _22380_);
  nand _54782_ (_22387_, _22386_, _22378_);
  nor _54783_ (_22388_, _22387_, _21523_);
  nand _54784_ (_22389_, _22388_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or _54785_ (_22390_, _22388_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _54786_ (_22391_, _22390_, _22389_);
  or _54787_ (_22392_, _22391_, _22370_);
  or _54788_ (_22393_, _22392_, _22349_);
  and _54789_ (_22394_, _21646_, _20681_);
  or _54790_ (_22395_, _22394_, _20946_);
  and _54791_ (_22396_, _21650_, _20656_);
  and _54792_ (_22397_, _21642_, _21527_);
  and _54793_ (_22398_, _21654_, _20682_);
  or _54794_ (_22399_, _22398_, _22397_);
  or _54795_ (_22400_, _22399_, _22396_);
  or _54796_ (_22401_, _22400_, _22395_);
  and _54797_ (_22402_, _21666_, _20681_);
  or _54798_ (_22403_, _22402_, _20676_);
  and _54799_ (_22404_, _21670_, _20656_);
  and _54800_ (_22405_, _21662_, _21527_);
  and _54801_ (_22406_, _21674_, _20682_);
  or _54802_ (_22407_, _22406_, _22405_);
  or _54803_ (_22408_, _22407_, _22404_);
  or _54804_ (_22409_, _22408_, _22403_);
  nand _54805_ (_22410_, _22409_, _22401_);
  nor _54806_ (_22411_, _22410_, _21523_);
  nand _54807_ (_22412_, _22411_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _54808_ (_22413_, _22411_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _54809_ (_22414_, _22413_, _22412_);
  and _54810_ (_22415_, _21704_, _21527_);
  and _54811_ (_22416_, _21716_, _20682_);
  and _54812_ (_22417_, _21712_, _20656_);
  and _54813_ (_22418_, _21708_, _20681_);
  or _54814_ (_22419_, _22418_, _22417_);
  or _54815_ (_22420_, _22419_, _22416_);
  or _54816_ (_22421_, _22420_, _22415_);
  and _54817_ (_22422_, _22421_, _20946_);
  and _54818_ (_22423_, _21684_, _21527_);
  and _54819_ (_22424_, _21696_, _20682_);
  and _54820_ (_22425_, _21692_, _20656_);
  and _54821_ (_22426_, _21688_, _20681_);
  or _54822_ (_22427_, _22426_, _22425_);
  or _54823_ (_22428_, _22427_, _22424_);
  or _54824_ (_22429_, _22428_, _22423_);
  and _54825_ (_22430_, _22429_, _20676_);
  or _54826_ (_22431_, _22430_, _22422_);
  and _54827_ (_22432_, _22431_, _22327_);
  and _54828_ (_22433_, _22432_, _22783_);
  nor _54829_ (_22434_, _22432_, _22783_);
  or _54830_ (_22435_, _22434_, _22433_);
  or _54831_ (_22436_, _22435_, _22414_);
  and _54832_ (_22437_, _21588_, _20682_);
  and _54833_ (_22438_, _21579_, _20681_);
  nor _54834_ (_22439_, _22438_, _22437_);
  and _54835_ (_22440_, _21584_, _21527_);
  and _54836_ (_22441_, _21574_, _20656_);
  nor _54837_ (_22442_, _22441_, _22440_);
  and _54838_ (_22443_, _22442_, _22439_);
  nor _54839_ (_22444_, _22443_, _20676_);
  and _54840_ (_22445_, _21567_, _20682_);
  and _54841_ (_22446_, _21558_, _20681_);
  nor _54842_ (_22447_, _22446_, _22445_);
  and _54843_ (_22448_, _21563_, _21527_);
  and _54844_ (_22449_, _21553_, _20656_);
  nor _54845_ (_22450_, _22449_, _22448_);
  and _54846_ (_22451_, _22450_, _22447_);
  nor _54847_ (_22452_, _22451_, _20946_);
  nor _54848_ (_22453_, _22452_, _22444_);
  nor _54849_ (_22454_, _22453_, _21523_);
  and _54850_ (_22455_, _22454_, _22778_);
  nor _54851_ (_22456_, _22454_, _22778_);
  or _54852_ (_22457_, _22456_, _22455_);
  and _54853_ (_22458_, _21607_, _20681_);
  or _54854_ (_22459_, _22458_, _20946_);
  and _54855_ (_22460_, _21611_, _20656_);
  and _54856_ (_22461_, _21602_, _21527_);
  and _54857_ (_22462_, _21597_, _20682_);
  or _54858_ (_22463_, _22462_, _22461_);
  or _54859_ (_22464_, _22463_, _22460_);
  or _54860_ (_22465_, _22464_, _22459_);
  and _54861_ (_22466_, _21628_, _20681_);
  or _54862_ (_22467_, _22466_, _20676_);
  and _54863_ (_22468_, _21632_, _20656_);
  and _54864_ (_22469_, _21623_, _21527_);
  and _54865_ (_22470_, _21618_, _20682_);
  or _54866_ (_22471_, _22470_, _22469_);
  or _54867_ (_22472_, _22471_, _22468_);
  or _54868_ (_22473_, _22472_, _22467_);
  nand _54869_ (_22474_, _22473_, _22465_);
  nor _54870_ (_22475_, _22474_, _21523_);
  and _54871_ (_22476_, _22475_, _22772_);
  nor _54872_ (_22477_, _22475_, _22772_);
  or _54873_ (_22478_, _22477_, _22476_);
  or _54874_ (_22479_, _22478_, _22457_);
  or _54875_ (_22480_, _22479_, _22436_);
  or _54876_ (_22481_, _22480_, _22393_);
  or _54877_ (_22482_, _21066_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _54878_ (_22483_, _21066_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _54879_ (_22484_, _22483_, _22482_);
  and _54880_ (_22485_, _21105_, _22810_);
  nor _54881_ (_22486_, _21105_, _22810_);
  or _54882_ (_22487_, _22486_, _22485_);
  or _54883_ (_22488_, _22487_, _22484_);
  or _54884_ (_22489_, _20984_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _54885_ (_22490_, _20984_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _54886_ (_22491_, _22490_, _22489_);
  nor _54887_ (_22492_, _21027_, _22819_);
  and _54888_ (_22493_, _21027_, _22819_);
  or _54889_ (_22494_, _22493_, _22492_);
  or _54890_ (_22495_, _22494_, _22491_);
  or _54891_ (_22496_, _22495_, _22488_);
  and _54892_ (_22497_, _20942_, _22827_);
  nor _54893_ (_22498_, _20942_, _22827_);
  or _54894_ (_22499_, _22498_, _22497_);
  or _54895_ (_22500_, _20900_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _54896_ (_22501_, _20900_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _54897_ (_22502_, _22501_, _22500_);
  or _54898_ (_22503_, _22502_, _22499_);
  and _54899_ (_22504_, _20775_, _14710_);
  nor _54900_ (_22505_, _20775_, _14710_);
  or _54901_ (_22506_, _22505_, _22504_);
  and _54902_ (_22507_, _20855_, _22837_);
  nor _54903_ (_22508_, _20855_, _22837_);
  or _54904_ (_22509_, _22508_, _22507_);
  or _54905_ (_22510_, _22509_, _22506_);
  or _54906_ (_22511_, _22510_, _22503_);
  or _54907_ (_22512_, _22511_, _22496_);
  or _54908_ (_22513_, _22512_, _22481_);
  and _54909_ (_22514_, _22038_, _21933_);
  and _54910_ (_22515_, _22514_, _22513_);
  or _54911_ (_22516_, _22515_, _22305_);
  and _54912_ (_22517_, _22516_, _21550_);
  or _54913_ (_22518_, _22517_, _22257_);
  or _54914_ (property_invalid, _22518_, _21906_);
  and _54915_ (_22519_, _24121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  not _54916_ (_22520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _54917_ (_22521_, _25687_, _25024_);
  nor _54918_ (_22522_, _22521_, _22520_);
  and _54919_ (_22523_, _22521_, _22520_);
  nor _54920_ (_22524_, _22523_, _22522_);
  nor _54921_ (_22525_, _22524_, _24127_);
  and _54922_ (_22526_, _24127_, _23642_);
  or _54923_ (_22527_, _22526_, _22525_);
  and _54924_ (_22528_, _22527_, _24166_);
  or _54925_ (_12540_, _22528_, _22519_);
  and _54926_ (_22529_, _03300_, _23707_);
  and _54927_ (_22530_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or _54928_ (_12543_, _22530_, _22529_);
  and _54929_ (_22531_, _18217_, _23946_);
  and _54930_ (_22532_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or _54931_ (_12545_, _22532_, _22531_);
  and _54932_ (_22533_, _21544_, first_instr);
  or _54933_ (_00000_, _22533_, rst);
  and _54934_ (_22534_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  and _54935_ (_22535_, _16331_, _23707_);
  or _54936_ (_12565_, _22535_, _22534_);
  and _54937_ (_22536_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  and _54938_ (_22537_, _16331_, _24050_);
  or _54939_ (_12569_, _22537_, _22536_);
  and _54940_ (_22538_, _18217_, _23649_);
  and _54941_ (_22539_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or _54942_ (_12586_, _22539_, _22538_);
  and _54943_ (_22540_, _25739_, _24050_);
  and _54944_ (_22541_, _25741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  or _54945_ (_12613_, _22541_, _22540_);
  and _54946_ (_22543_, _03300_, _24050_);
  and _54947_ (_22544_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or _54948_ (_12615_, _22544_, _22543_);
  and _54949_ (_22545_, _16326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and _54950_ (_22546_, _16325_, _23778_);
  or _54951_ (_12617_, _22546_, _22545_);
  and _54952_ (_22547_, _18217_, _23747_);
  and _54953_ (_22548_, _18219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or _54954_ (_27215_, _22548_, _22547_);
  and _54955_ (_22549_, _10347_, _23824_);
  and _54956_ (_22550_, _10350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  or _54957_ (_12632_, _22550_, _22549_);
  and _54958_ (_22551_, _08548_, _23778_);
  and _54959_ (_22552_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  or _54960_ (_27136_, _22552_, _22551_);
  and _54961_ (_22553_, _06508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and _54962_ (_22554_, _06507_, _23649_);
  or _54963_ (_12672_, _22554_, _22553_);
  and _54964_ (_22555_, _03300_, _23946_);
  and _54965_ (_22556_, _03302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or _54966_ (_12674_, _22556_, _22555_);
  and _54967_ (_22557_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  and _54968_ (_22558_, _16331_, _23898_);
  or _54969_ (_12679_, _22558_, _22557_);
  and _54970_ (_22559_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  and _54971_ (_22560_, _16331_, _23778_);
  or _54972_ (_12681_, _22560_, _22559_);
  and _54973_ (_22561_, _08548_, _23824_);
  and _54974_ (_22562_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  or _54975_ (_12704_, _22562_, _22561_);
  and _54976_ (_22563_, _08548_, _23898_);
  and _54977_ (_22564_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  or _54978_ (_12706_, _22564_, _22563_);
  and _54979_ (_22565_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  and _54980_ (_22566_, _16331_, _23649_);
  or _54981_ (_12711_, _22566_, _22565_);
  or _54982_ (_22567_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _54983_ (_22568_, _22567_, _22762_);
  or _54984_ (_22569_, _24079_, _23892_);
  and _54985_ (_12717_, _22569_, _22568_);
  nand _54986_ (_22570_, _24073_, _23772_);
  or _54987_ (_22571_, _24073_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _54988_ (_22572_, _22571_, _22762_);
  and _54989_ (_12720_, _22572_, _22570_);
  and _54990_ (_22573_, _16332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  and _54991_ (_22574_, _16331_, _23747_);
  or _54992_ (_26966_, _22574_, _22573_);
  and _54993_ (_22575_, _25748_, _23707_);
  and _54994_ (_22576_, _25750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or _54995_ (_27070_, _22576_, _22575_);
  or _54996_ (_22577_, _04891_, _23892_);
  and _54997_ (_22578_, _26115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _54998_ (_22579_, _22578_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _54999_ (_22580_, _04880_, _26098_);
  and _55000_ (_22581_, _22580_, _22579_);
  and _55001_ (_22582_, _24300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _55002_ (_22583_, _22582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not _55003_ (_22584_, _14815_);
  and _55004_ (_22585_, _22584_, _24302_);
  and _55005_ (_22586_, _22585_, _22583_);
  not _55006_ (_22587_, _14810_);
  and _55007_ (_22588_, _22587_, _04860_);
  or _55008_ (_22589_, _22588_, _26100_);
  and _55009_ (_22590_, _26110_, _26099_);
  and _55010_ (_22591_, _22590_, _15862_);
  or _55011_ (_22592_, _22591_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _55012_ (_22593_, _22592_, _22589_);
  or _55013_ (_22594_, _22593_, _22586_);
  or _55014_ (_22595_, _22594_, _22581_);
  or _55015_ (_22596_, _22595_, _24299_);
  and _55016_ (_22597_, _22596_, _24294_);
  and _55017_ (_22598_, _22597_, _22577_);
  and _55018_ (_22599_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _55019_ (_22600_, _22599_, _22598_);
  and _55020_ (_12731_, _22600_, _22762_);
  not _55021_ (_22601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _55022_ (_22602_, _26115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _55023_ (_22603_, _22602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _55024_ (_22604_, _22603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  nand _55025_ (_22605_, _22604_, _26099_);
  nand _55026_ (_22606_, _22605_, _22601_);
  or _55027_ (_22607_, _22605_, _22601_);
  and _55028_ (_22608_, _22607_, _22606_);
  and _55029_ (_22609_, _22608_, _04861_);
  or _55030_ (_22610_, _24300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not _55031_ (_22611_, _22582_);
  and _55032_ (_22612_, _22611_, _24302_);
  and _55033_ (_22613_, _22612_, _22610_);
  or _55034_ (_22614_, _26115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _55035_ (_22615_, _22578_, _26098_);
  and _55036_ (_22616_, _22615_, _22614_);
  or _55037_ (_22617_, _22616_, _22613_);
  or _55038_ (_22618_, _22617_, _22609_);
  or _55039_ (_22619_, _22618_, _24299_);
  nand _55040_ (_22620_, _24299_, _23772_);
  and _55041_ (_22621_, _22620_, _24294_);
  and _55042_ (_22622_, _22621_, _22619_);
  and _55043_ (_22623_, _24293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _55044_ (_22624_, _22623_, _22622_);
  and _55045_ (_12736_, _22624_, _22762_);
  and _55046_ (_22625_, _05042_, _23649_);
  and _55047_ (_22626_, _05045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or _55048_ (_12741_, _22626_, _22625_);
  dff _55049_ (first_instr, _00000_, clk);
  dff _55050_ (\oc8051_symbolic_cxrom1.regarray[0] [0], _26843_[0], clk);
  dff _55051_ (\oc8051_symbolic_cxrom1.regarray[0] [1], _26843_[1], clk);
  dff _55052_ (\oc8051_symbolic_cxrom1.regarray[0] [2], _26843_[2], clk);
  dff _55053_ (\oc8051_symbolic_cxrom1.regarray[0] [3], _26843_[3], clk);
  dff _55054_ (\oc8051_symbolic_cxrom1.regarray[0] [4], _26843_[4], clk);
  dff _55055_ (\oc8051_symbolic_cxrom1.regarray[0] [5], _26843_[5], clk);
  dff _55056_ (\oc8051_symbolic_cxrom1.regarray[0] [6], _26843_[6], clk);
  dff _55057_ (\oc8051_symbolic_cxrom1.regarray[0] [7], _26843_[7], clk);
  dff _55058_ (\oc8051_symbolic_cxrom1.regvalid [0], _26859_, clk);
  dff _55059_ (\oc8051_symbolic_cxrom1.regvalid [1], _26842_[1], clk);
  dff _55060_ (\oc8051_symbolic_cxrom1.regvalid [2], _26842_[2], clk);
  dff _55061_ (\oc8051_symbolic_cxrom1.regvalid [3], _26842_[3], clk);
  dff _55062_ (\oc8051_symbolic_cxrom1.regvalid [4], _26842_[4], clk);
  dff _55063_ (\oc8051_symbolic_cxrom1.regvalid [5], _26842_[5], clk);
  dff _55064_ (\oc8051_symbolic_cxrom1.regvalid [6], _26842_[6], clk);
  dff _55065_ (\oc8051_symbolic_cxrom1.regvalid [7], _26842_[7], clk);
  dff _55066_ (\oc8051_symbolic_cxrom1.regvalid [8], _26842_[8], clk);
  dff _55067_ (\oc8051_symbolic_cxrom1.regvalid [9], _26842_[9], clk);
  dff _55068_ (\oc8051_symbolic_cxrom1.regvalid [10], _26842_[10], clk);
  dff _55069_ (\oc8051_symbolic_cxrom1.regvalid [11], _26842_[11], clk);
  dff _55070_ (\oc8051_symbolic_cxrom1.regvalid [12], _26842_[12], clk);
  dff _55071_ (\oc8051_symbolic_cxrom1.regvalid [13], _26842_[13], clk);
  dff _55072_ (\oc8051_symbolic_cxrom1.regvalid [14], _26842_[14], clk);
  dff _55073_ (\oc8051_symbolic_cxrom1.regvalid [15], _26842_[15], clk);
  dff _55074_ (\oc8051_symbolic_cxrom1.regarray[1] [0], _26850_[0], clk);
  dff _55075_ (\oc8051_symbolic_cxrom1.regarray[1] [1], _26850_[1], clk);
  dff _55076_ (\oc8051_symbolic_cxrom1.regarray[1] [2], _26850_[2], clk);
  dff _55077_ (\oc8051_symbolic_cxrom1.regarray[1] [3], _26850_[3], clk);
  dff _55078_ (\oc8051_symbolic_cxrom1.regarray[1] [4], _26850_[4], clk);
  dff _55079_ (\oc8051_symbolic_cxrom1.regarray[1] [5], _26850_[5], clk);
  dff _55080_ (\oc8051_symbolic_cxrom1.regarray[1] [6], _26850_[6], clk);
  dff _55081_ (\oc8051_symbolic_cxrom1.regarray[1] [7], _26850_[7], clk);
  dff _55082_ (\oc8051_symbolic_cxrom1.regarray[2] [0], _26851_[0], clk);
  dff _55083_ (\oc8051_symbolic_cxrom1.regarray[2] [1], _26851_[1], clk);
  dff _55084_ (\oc8051_symbolic_cxrom1.regarray[2] [2], _26851_[2], clk);
  dff _55085_ (\oc8051_symbolic_cxrom1.regarray[2] [3], _26851_[3], clk);
  dff _55086_ (\oc8051_symbolic_cxrom1.regarray[2] [4], _26851_[4], clk);
  dff _55087_ (\oc8051_symbolic_cxrom1.regarray[2] [5], _26851_[5], clk);
  dff _55088_ (\oc8051_symbolic_cxrom1.regarray[2] [6], _26851_[6], clk);
  dff _55089_ (\oc8051_symbolic_cxrom1.regarray[2] [7], _26851_[7], clk);
  dff _55090_ (\oc8051_symbolic_cxrom1.regarray[3] [0], _26852_[0], clk);
  dff _55091_ (\oc8051_symbolic_cxrom1.regarray[3] [1], _26852_[1], clk);
  dff _55092_ (\oc8051_symbolic_cxrom1.regarray[3] [2], _26852_[2], clk);
  dff _55093_ (\oc8051_symbolic_cxrom1.regarray[3] [3], _26852_[3], clk);
  dff _55094_ (\oc8051_symbolic_cxrom1.regarray[3] [4], _26852_[4], clk);
  dff _55095_ (\oc8051_symbolic_cxrom1.regarray[3] [5], _26852_[5], clk);
  dff _55096_ (\oc8051_symbolic_cxrom1.regarray[3] [6], _26852_[6], clk);
  dff _55097_ (\oc8051_symbolic_cxrom1.regarray[3] [7], _26852_[7], clk);
  dff _55098_ (\oc8051_symbolic_cxrom1.regarray[4] [0], _26853_[0], clk);
  dff _55099_ (\oc8051_symbolic_cxrom1.regarray[4] [1], _26853_[1], clk);
  dff _55100_ (\oc8051_symbolic_cxrom1.regarray[4] [2], _26853_[2], clk);
  dff _55101_ (\oc8051_symbolic_cxrom1.regarray[4] [3], _26853_[3], clk);
  dff _55102_ (\oc8051_symbolic_cxrom1.regarray[4] [4], _26853_[4], clk);
  dff _55103_ (\oc8051_symbolic_cxrom1.regarray[4] [5], _26853_[5], clk);
  dff _55104_ (\oc8051_symbolic_cxrom1.regarray[4] [6], _26853_[6], clk);
  dff _55105_ (\oc8051_symbolic_cxrom1.regarray[4] [7], _26853_[7], clk);
  dff _55106_ (\oc8051_symbolic_cxrom1.regarray[5] [0], _26854_[0], clk);
  dff _55107_ (\oc8051_symbolic_cxrom1.regarray[5] [1], _26854_[1], clk);
  dff _55108_ (\oc8051_symbolic_cxrom1.regarray[5] [2], _26854_[2], clk);
  dff _55109_ (\oc8051_symbolic_cxrom1.regarray[5] [3], _26854_[3], clk);
  dff _55110_ (\oc8051_symbolic_cxrom1.regarray[5] [4], _26854_[4], clk);
  dff _55111_ (\oc8051_symbolic_cxrom1.regarray[5] [5], _26854_[5], clk);
  dff _55112_ (\oc8051_symbolic_cxrom1.regarray[5] [6], _26854_[6], clk);
  dff _55113_ (\oc8051_symbolic_cxrom1.regarray[5] [7], _26854_[7], clk);
  dff _55114_ (\oc8051_symbolic_cxrom1.regarray[6] [0], _26855_[0], clk);
  dff _55115_ (\oc8051_symbolic_cxrom1.regarray[6] [1], _26855_[1], clk);
  dff _55116_ (\oc8051_symbolic_cxrom1.regarray[6] [2], _26855_[2], clk);
  dff _55117_ (\oc8051_symbolic_cxrom1.regarray[6] [3], _26855_[3], clk);
  dff _55118_ (\oc8051_symbolic_cxrom1.regarray[6] [4], _26855_[4], clk);
  dff _55119_ (\oc8051_symbolic_cxrom1.regarray[6] [5], _26855_[5], clk);
  dff _55120_ (\oc8051_symbolic_cxrom1.regarray[6] [6], _26855_[6], clk);
  dff _55121_ (\oc8051_symbolic_cxrom1.regarray[6] [7], _26855_[7], clk);
  dff _55122_ (\oc8051_symbolic_cxrom1.regarray[7] [0], _26856_[0], clk);
  dff _55123_ (\oc8051_symbolic_cxrom1.regarray[7] [1], _26856_[1], clk);
  dff _55124_ (\oc8051_symbolic_cxrom1.regarray[7] [2], _26856_[2], clk);
  dff _55125_ (\oc8051_symbolic_cxrom1.regarray[7] [3], _26856_[3], clk);
  dff _55126_ (\oc8051_symbolic_cxrom1.regarray[7] [4], _26856_[4], clk);
  dff _55127_ (\oc8051_symbolic_cxrom1.regarray[7] [5], _26856_[5], clk);
  dff _55128_ (\oc8051_symbolic_cxrom1.regarray[7] [6], _26856_[6], clk);
  dff _55129_ (\oc8051_symbolic_cxrom1.regarray[7] [7], _26856_[7], clk);
  dff _55130_ (\oc8051_symbolic_cxrom1.regarray[8] [0], _26857_[0], clk);
  dff _55131_ (\oc8051_symbolic_cxrom1.regarray[8] [1], _26857_[1], clk);
  dff _55132_ (\oc8051_symbolic_cxrom1.regarray[8] [2], _26857_[2], clk);
  dff _55133_ (\oc8051_symbolic_cxrom1.regarray[8] [3], _26857_[3], clk);
  dff _55134_ (\oc8051_symbolic_cxrom1.regarray[8] [4], _26857_[4], clk);
  dff _55135_ (\oc8051_symbolic_cxrom1.regarray[8] [5], _26857_[5], clk);
  dff _55136_ (\oc8051_symbolic_cxrom1.regarray[8] [6], _26857_[6], clk);
  dff _55137_ (\oc8051_symbolic_cxrom1.regarray[8] [7], _26857_[7], clk);
  dff _55138_ (\oc8051_symbolic_cxrom1.regarray[9] [0], _26858_[0], clk);
  dff _55139_ (\oc8051_symbolic_cxrom1.regarray[9] [1], _26858_[1], clk);
  dff _55140_ (\oc8051_symbolic_cxrom1.regarray[9] [2], _26858_[2], clk);
  dff _55141_ (\oc8051_symbolic_cxrom1.regarray[9] [3], _26858_[3], clk);
  dff _55142_ (\oc8051_symbolic_cxrom1.regarray[9] [4], _26858_[4], clk);
  dff _55143_ (\oc8051_symbolic_cxrom1.regarray[9] [5], _26858_[5], clk);
  dff _55144_ (\oc8051_symbolic_cxrom1.regarray[9] [6], _26858_[6], clk);
  dff _55145_ (\oc8051_symbolic_cxrom1.regarray[9] [7], _26858_[7], clk);
  dff _55146_ (\oc8051_symbolic_cxrom1.regarray[10] [0], _26844_[0], clk);
  dff _55147_ (\oc8051_symbolic_cxrom1.regarray[10] [1], _26844_[1], clk);
  dff _55148_ (\oc8051_symbolic_cxrom1.regarray[10] [2], _26844_[2], clk);
  dff _55149_ (\oc8051_symbolic_cxrom1.regarray[10] [3], _26844_[3], clk);
  dff _55150_ (\oc8051_symbolic_cxrom1.regarray[10] [4], _26844_[4], clk);
  dff _55151_ (\oc8051_symbolic_cxrom1.regarray[10] [5], _26844_[5], clk);
  dff _55152_ (\oc8051_symbolic_cxrom1.regarray[10] [6], _26844_[6], clk);
  dff _55153_ (\oc8051_symbolic_cxrom1.regarray[10] [7], _26844_[7], clk);
  dff _55154_ (\oc8051_symbolic_cxrom1.regarray[11] [0], _26845_[0], clk);
  dff _55155_ (\oc8051_symbolic_cxrom1.regarray[11] [1], _26845_[1], clk);
  dff _55156_ (\oc8051_symbolic_cxrom1.regarray[11] [2], _26845_[2], clk);
  dff _55157_ (\oc8051_symbolic_cxrom1.regarray[11] [3], _26845_[3], clk);
  dff _55158_ (\oc8051_symbolic_cxrom1.regarray[11] [4], _26845_[4], clk);
  dff _55159_ (\oc8051_symbolic_cxrom1.regarray[11] [5], _26845_[5], clk);
  dff _55160_ (\oc8051_symbolic_cxrom1.regarray[11] [6], _26845_[6], clk);
  dff _55161_ (\oc8051_symbolic_cxrom1.regarray[11] [7], _26845_[7], clk);
  dff _55162_ (\oc8051_symbolic_cxrom1.regarray[12] [0], _26846_[0], clk);
  dff _55163_ (\oc8051_symbolic_cxrom1.regarray[12] [1], _26846_[1], clk);
  dff _55164_ (\oc8051_symbolic_cxrom1.regarray[12] [2], _26846_[2], clk);
  dff _55165_ (\oc8051_symbolic_cxrom1.regarray[12] [3], _26846_[3], clk);
  dff _55166_ (\oc8051_symbolic_cxrom1.regarray[12] [4], _26846_[4], clk);
  dff _55167_ (\oc8051_symbolic_cxrom1.regarray[12] [5], _26846_[5], clk);
  dff _55168_ (\oc8051_symbolic_cxrom1.regarray[12] [6], _26846_[6], clk);
  dff _55169_ (\oc8051_symbolic_cxrom1.regarray[12] [7], _26846_[7], clk);
  dff _55170_ (\oc8051_symbolic_cxrom1.regarray[13] [0], _26847_[0], clk);
  dff _55171_ (\oc8051_symbolic_cxrom1.regarray[13] [1], _26847_[1], clk);
  dff _55172_ (\oc8051_symbolic_cxrom1.regarray[13] [2], _26847_[2], clk);
  dff _55173_ (\oc8051_symbolic_cxrom1.regarray[13] [3], _26847_[3], clk);
  dff _55174_ (\oc8051_symbolic_cxrom1.regarray[13] [4], _26847_[4], clk);
  dff _55175_ (\oc8051_symbolic_cxrom1.regarray[13] [5], _26847_[5], clk);
  dff _55176_ (\oc8051_symbolic_cxrom1.regarray[13] [6], _26847_[6], clk);
  dff _55177_ (\oc8051_symbolic_cxrom1.regarray[13] [7], _26847_[7], clk);
  dff _55178_ (\oc8051_symbolic_cxrom1.regarray[14] [0], _26848_[0], clk);
  dff _55179_ (\oc8051_symbolic_cxrom1.regarray[14] [1], _26848_[1], clk);
  dff _55180_ (\oc8051_symbolic_cxrom1.regarray[14] [2], _26848_[2], clk);
  dff _55181_ (\oc8051_symbolic_cxrom1.regarray[14] [3], _26848_[3], clk);
  dff _55182_ (\oc8051_symbolic_cxrom1.regarray[14] [4], _26848_[4], clk);
  dff _55183_ (\oc8051_symbolic_cxrom1.regarray[14] [5], _26848_[5], clk);
  dff _55184_ (\oc8051_symbolic_cxrom1.regarray[14] [6], _26848_[6], clk);
  dff _55185_ (\oc8051_symbolic_cxrom1.regarray[14] [7], _26848_[7], clk);
  dff _55186_ (\oc8051_symbolic_cxrom1.regarray[15] [0], _26849_[0], clk);
  dff _55187_ (\oc8051_symbolic_cxrom1.regarray[15] [1], _26849_[1], clk);
  dff _55188_ (\oc8051_symbolic_cxrom1.regarray[15] [2], _26849_[2], clk);
  dff _55189_ (\oc8051_symbolic_cxrom1.regarray[15] [3], _26849_[3], clk);
  dff _55190_ (\oc8051_symbolic_cxrom1.regarray[15] [4], _26849_[4], clk);
  dff _55191_ (\oc8051_symbolic_cxrom1.regarray[15] [5], _26849_[5], clk);
  dff _55192_ (\oc8051_symbolic_cxrom1.regarray[15] [6], _26849_[6], clk);
  dff _55193_ (\oc8051_symbolic_cxrom1.regarray[15] [7], _26849_[7], clk);
  dff _55194_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _11665_, clk);
  dff _55195_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _11643_, clk);
  dff _55196_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _09312_, clk);
  dff _55197_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _11604_, clk);
  dff _55198_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _11662_, clk);
  dff _55199_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _09317_, clk);
  dff _55200_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _09321_, clk);
  dff _55201_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _09302_, clk);
  dff _55202_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _11859_, clk);
  dff _55203_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _11759_, clk);
  dff _55204_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _11830_, clk);
  dff _55205_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _11817_, clk);
  dff _55206_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _11872_, clk);
  dff _55207_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _11857_, clk);
  dff _55208_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _11758_, clk);
  dff _55209_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _09315_, clk);
  dff _55210_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _12022_, clk);
  dff _55211_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22706_, clk);
  dff _55212_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _12035_, clk);
  dff _55213_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _12290_, clk);
  dff _55214_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _12040_, clk);
  dff _55215_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _12052_, clk);
  dff _55216_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _12026_, clk);
  dff _55217_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _12042_, clk);
  dff _55218_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _12048_, clk);
  dff _55219_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _12054_, clk);
  dff _55220_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _12050_, clk);
  dff _55221_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _12044_, clk);
  dff _55222_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _12037_, clk);
  dff _55223_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _12060_, clk);
  dff _55224_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _12056_, clk);
  dff _55225_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _12086_, clk);
  dff _55226_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _26860_[0], clk);
  dff _55227_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _26860_[1], clk);
  dff _55228_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _26860_[2], clk);
  dff _55229_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _26860_[3], clk);
  dff _55230_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _26860_[4], clk);
  dff _55231_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _26860_[5], clk);
  dff _55232_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _26860_[6], clk);
  dff _55233_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _26860_[7], clk);
  dff _55234_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _26887_[0], clk);
  dff _55235_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _26887_[1], clk);
  dff _55236_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _26887_[2], clk);
  dff _55237_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _26887_[3], clk);
  dff _55238_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _26887_[4], clk);
  dff _55239_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _26887_[5], clk);
  dff _55240_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _26887_[6], clk);
  dff _55241_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _26887_[7], clk);
  dff _55242_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _26897_[0], clk);
  dff _55243_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _26897_[1], clk);
  dff _55244_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _26897_[2], clk);
  dff _55245_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _26897_[3], clk);
  dff _55246_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _26897_[4], clk);
  dff _55247_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _26897_[5], clk);
  dff _55248_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _26897_[6], clk);
  dff _55249_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _26897_[7], clk);
  dff _55250_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _26867_[0], clk);
  dff _55251_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _26867_[1], clk);
  dff _55252_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _26868_[0], clk);
  dff _55253_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _26868_[1], clk);
  dff _55254_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _26868_[2], clk);
  dff _55255_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _26869_[0], clk);
  dff _55256_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _26869_[1], clk);
  dff _55257_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _26869_[2], clk);
  dff _55258_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _26870_[0], clk);
  dff _55259_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _26870_[1], clk);
  dff _55260_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _26871_[0], clk);
  dff _55261_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _26871_[1], clk);
  dff _55262_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _26871_[2], clk);
  dff _55263_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _26871_[3], clk);
  dff _55264_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _26872_[0], clk);
  dff _55265_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _26872_[1], clk);
  dff _55266_ (\oc8051_top_1.oc8051_decoder1.wr , _26873_, clk);
  dff _55267_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _26861_[0], clk);
  dff _55268_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _26861_[1], clk);
  dff _55269_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _26861_[2], clk);
  dff _55270_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _26862_[0], clk);
  dff _55271_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _26862_[1], clk);
  dff _55272_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _26862_[2], clk);
  dff _55273_ (\oc8051_top_1.oc8051_decoder1.state [0], _26863_[0], clk);
  dff _55274_ (\oc8051_top_1.oc8051_decoder1.state [1], _26863_[1], clk);
  dff _55275_ (\oc8051_top_1.oc8051_decoder1.op [0], _26864_[0], clk);
  dff _55276_ (\oc8051_top_1.oc8051_decoder1.op [1], _26864_[1], clk);
  dff _55277_ (\oc8051_top_1.oc8051_decoder1.op [2], _26864_[2], clk);
  dff _55278_ (\oc8051_top_1.oc8051_decoder1.op [3], _26864_[3], clk);
  dff _55279_ (\oc8051_top_1.oc8051_decoder1.op [4], _26864_[4], clk);
  dff _55280_ (\oc8051_top_1.oc8051_decoder1.op [5], _26864_[5], clk);
  dff _55281_ (\oc8051_top_1.oc8051_decoder1.op [6], _26864_[6], clk);
  dff _55282_ (\oc8051_top_1.oc8051_decoder1.op [7], _26864_[7], clk);
  dff _55283_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _26865_, clk);
  dff _55284_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _26866_[0], clk);
  dff _55285_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _26866_[1], clk);
  dff _55286_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _26912_, clk);
  dff _55287_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _26874_[0], clk);
  dff _55288_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _26874_[1], clk);
  dff _55289_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _26874_[2], clk);
  dff _55290_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _26874_[3], clk);
  dff _55291_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _26874_[4], clk);
  dff _55292_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _26874_[5], clk);
  dff _55293_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _26874_[6], clk);
  dff _55294_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _26874_[7], clk);
  dff _55295_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _26875_[0], clk);
  dff _55296_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _26875_[1], clk);
  dff _55297_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _26875_[2], clk);
  dff _55298_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _26875_[3], clk);
  dff _55299_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _26875_[4], clk);
  dff _55300_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _26875_[5], clk);
  dff _55301_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _26875_[6], clk);
  dff _55302_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _26875_[7], clk);
  dff _55303_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _26876_[0], clk);
  dff _55304_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _26876_[1], clk);
  dff _55305_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _26876_[2], clk);
  dff _55306_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _26876_[3], clk);
  dff _55307_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _26876_[4], clk);
  dff _55308_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _26876_[5], clk);
  dff _55309_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _26876_[6], clk);
  dff _55310_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _26876_[7], clk);
  dff _55311_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _26877_[0], clk);
  dff _55312_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _26877_[1], clk);
  dff _55313_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _26877_[2], clk);
  dff _55314_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _26877_[3], clk);
  dff _55315_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _26877_[4], clk);
  dff _55316_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _26877_[5], clk);
  dff _55317_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _26877_[6], clk);
  dff _55318_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _26877_[7], clk);
  dff _55319_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _26878_[0], clk);
  dff _55320_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _26878_[1], clk);
  dff _55321_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _26878_[2], clk);
  dff _55322_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _26878_[3], clk);
  dff _55323_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _26878_[4], clk);
  dff _55324_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _26878_[5], clk);
  dff _55325_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _26878_[6], clk);
  dff _55326_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _26878_[7], clk);
  dff _55327_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _26879_[0], clk);
  dff _55328_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _26879_[1], clk);
  dff _55329_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _26879_[2], clk);
  dff _55330_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _26879_[3], clk);
  dff _55331_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _26879_[4], clk);
  dff _55332_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _26879_[5], clk);
  dff _55333_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _26879_[6], clk);
  dff _55334_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _26879_[7], clk);
  dff _55335_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _26880_[0], clk);
  dff _55336_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _26880_[1], clk);
  dff _55337_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _26880_[2], clk);
  dff _55338_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _26880_[3], clk);
  dff _55339_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _26880_[4], clk);
  dff _55340_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _26880_[5], clk);
  dff _55341_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _26880_[6], clk);
  dff _55342_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _26880_[7], clk);
  dff _55343_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _26881_[0], clk);
  dff _55344_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _26881_[1], clk);
  dff _55345_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _26881_[2], clk);
  dff _55346_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _26881_[3], clk);
  dff _55347_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _26881_[4], clk);
  dff _55348_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _26881_[5], clk);
  dff _55349_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _26881_[6], clk);
  dff _55350_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _26881_[7], clk);
  dff _55351_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _26885_[0], clk);
  dff _55352_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _26885_[1], clk);
  dff _55353_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _26885_[2], clk);
  dff _55354_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _26885_[3], clk);
  dff _55355_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _26885_[4], clk);
  dff _55356_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _26882_[0], clk);
  dff _55357_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _26882_[1], clk);
  dff _55358_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _26882_[2], clk);
  dff _55359_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _26882_[3], clk);
  dff _55360_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _26882_[4], clk);
  dff _55361_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _26882_[5], clk);
  dff _55362_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _26882_[6], clk);
  dff _55363_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _26882_[7], clk);
  dff _55364_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _26882_[8], clk);
  dff _55365_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _26882_[9], clk);
  dff _55366_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _26882_[10], clk);
  dff _55367_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _26882_[11], clk);
  dff _55368_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _26882_[12], clk);
  dff _55369_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _26882_[13], clk);
  dff _55370_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _26882_[14], clk);
  dff _55371_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _26882_[15], clk);
  dff _55372_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _26883_[0], clk);
  dff _55373_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _26883_[1], clk);
  dff _55374_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _26883_[2], clk);
  dff _55375_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _26883_[3], clk);
  dff _55376_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _26883_[4], clk);
  dff _55377_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _26883_[5], clk);
  dff _55378_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _26883_[6], clk);
  dff _55379_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _26883_[7], clk);
  dff _55380_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _26883_[8], clk);
  dff _55381_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _26883_[9], clk);
  dff _55382_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _26883_[10], clk);
  dff _55383_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _26883_[11], clk);
  dff _55384_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _26883_[12], clk);
  dff _55385_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _26883_[13], clk);
  dff _55386_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _26883_[14], clk);
  dff _55387_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _26883_[15], clk);
  dff _55388_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _26903_[0], clk);
  dff _55389_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _26903_[1], clk);
  dff _55390_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _26903_[2], clk);
  dff _55391_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _26903_[3], clk);
  dff _55392_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _26903_[4], clk);
  dff _55393_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _26903_[5], clk);
  dff _55394_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _26903_[6], clk);
  dff _55395_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _26903_[7], clk);
  dff _55396_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _26903_[8], clk);
  dff _55397_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _26903_[9], clk);
  dff _55398_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _26903_[10], clk);
  dff _55399_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _26903_[11], clk);
  dff _55400_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _26903_[12], clk);
  dff _55401_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _26903_[13], clk);
  dff _55402_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _26903_[14], clk);
  dff _55403_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _26903_[15], clk);
  dff _55404_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _26903_[16], clk);
  dff _55405_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _26903_[17], clk);
  dff _55406_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _26903_[18], clk);
  dff _55407_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _26903_[19], clk);
  dff _55408_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _26903_[20], clk);
  dff _55409_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _26903_[21], clk);
  dff _55410_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _26903_[22], clk);
  dff _55411_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _26903_[23], clk);
  dff _55412_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _26903_[24], clk);
  dff _55413_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _26903_[25], clk);
  dff _55414_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _26903_[26], clk);
  dff _55415_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _26903_[27], clk);
  dff _55416_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _26903_[28], clk);
  dff _55417_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _26903_[29], clk);
  dff _55418_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _26903_[30], clk);
  dff _55419_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _26903_[31], clk);
  dff _55420_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _26884_, clk);
  dff _55421_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _26886_[0], clk);
  dff _55422_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _26886_[1], clk);
  dff _55423_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _26886_[2], clk);
  dff _55424_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _26886_[3], clk);
  dff _55425_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _26886_[4], clk);
  dff _55426_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _26886_[5], clk);
  dff _55427_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _26886_[6], clk);
  dff _55428_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _26886_[7], clk);
  dff _55429_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _26888_, clk);
  dff _55430_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _26889_, clk);
  dff _55431_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _26890_[0], clk);
  dff _55432_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _26890_[1], clk);
  dff _55433_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _26890_[2], clk);
  dff _55434_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _26890_[3], clk);
  dff _55435_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _26890_[4], clk);
  dff _55436_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _26890_[5], clk);
  dff _55437_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _26890_[6], clk);
  dff _55438_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _26890_[7], clk);
  dff _55439_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _26890_[8], clk);
  dff _55440_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _26890_[9], clk);
  dff _55441_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _26890_[10], clk);
  dff _55442_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _26890_[11], clk);
  dff _55443_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _26890_[12], clk);
  dff _55444_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _26890_[13], clk);
  dff _55445_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _26890_[14], clk);
  dff _55446_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _26890_[15], clk);
  dff _55447_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _26891_[0], clk);
  dff _55448_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _26891_[1], clk);
  dff _55449_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _26891_[2], clk);
  dff _55450_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _26891_[3], clk);
  dff _55451_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _26891_[4], clk);
  dff _55452_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _26891_[5], clk);
  dff _55453_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _26891_[6], clk);
  dff _55454_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _26891_[7], clk);
  dff _55455_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _26891_[8], clk);
  dff _55456_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _26891_[9], clk);
  dff _55457_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _26891_[10], clk);
  dff _55458_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _26891_[11], clk);
  dff _55459_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _26891_[12], clk);
  dff _55460_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _26891_[13], clk);
  dff _55461_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _26891_[14], clk);
  dff _55462_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _26891_[15], clk);
  dff _55463_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _26892_, clk);
  dff _55464_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _26894_, clk);
  dff _55465_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _26893_, clk);
  dff _55466_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _26895_[0], clk);
  dff _55467_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _26895_[1], clk);
  dff _55468_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _26895_[2], clk);
  dff _55469_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _26895_[3], clk);
  dff _55470_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _26895_[4], clk);
  dff _55471_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _26895_[5], clk);
  dff _55472_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _26895_[6], clk);
  dff _55473_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _26895_[7], clk);
  dff _55474_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _26896_[0], clk);
  dff _55475_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _26896_[1], clk);
  dff _55476_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _26896_[2], clk);
  dff _55477_ (\oc8051_top_1.oc8051_memory_interface1.reti , _26898_, clk);
  dff _55478_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _26899_[0], clk);
  dff _55479_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _26899_[1], clk);
  dff _55480_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _26899_[2], clk);
  dff _55481_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _26899_[3], clk);
  dff _55482_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _26899_[4], clk);
  dff _55483_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _26899_[5], clk);
  dff _55484_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _26899_[6], clk);
  dff _55485_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _26899_[7], clk);
  dff _55486_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _26900_, clk);
  dff _55487_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _26901_, clk);
  dff _55488_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _26902_[0], clk);
  dff _55489_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _26902_[1], clk);
  dff _55490_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _26902_[2], clk);
  dff _55491_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _26902_[3], clk);
  dff _55492_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _26904_[0], clk);
  dff _55493_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _26904_[1], clk);
  dff _55494_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _26904_[2], clk);
  dff _55495_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _26904_[3], clk);
  dff _55496_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _26904_[4], clk);
  dff _55497_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _26904_[5], clk);
  dff _55498_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _26904_[6], clk);
  dff _55499_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _26904_[7], clk);
  dff _55500_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _26904_[8], clk);
  dff _55501_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _26904_[9], clk);
  dff _55502_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _26904_[10], clk);
  dff _55503_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _26904_[11], clk);
  dff _55504_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _26904_[12], clk);
  dff _55505_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _26904_[13], clk);
  dff _55506_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _26904_[14], clk);
  dff _55507_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _26904_[15], clk);
  dff _55508_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _26904_[16], clk);
  dff _55509_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _26904_[17], clk);
  dff _55510_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _26904_[18], clk);
  dff _55511_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _26904_[19], clk);
  dff _55512_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _26904_[20], clk);
  dff _55513_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _26904_[21], clk);
  dff _55514_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _26904_[22], clk);
  dff _55515_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _26904_[23], clk);
  dff _55516_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _26904_[24], clk);
  dff _55517_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _26904_[25], clk);
  dff _55518_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _26904_[26], clk);
  dff _55519_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _26904_[27], clk);
  dff _55520_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _26904_[28], clk);
  dff _55521_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _26904_[29], clk);
  dff _55522_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _26904_[30], clk);
  dff _55523_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _26904_[31], clk);
  dff _55524_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _26905_, clk);
  dff _55525_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _26906_, clk);
  dff _55526_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _26907_, clk);
  dff _55527_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _26908_[0], clk);
  dff _55528_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _26908_[1], clk);
  dff _55529_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _26908_[2], clk);
  dff _55530_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _26908_[3], clk);
  dff _55531_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _26909_, clk);
  dff _55532_ (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _26910_, clk);
  dff _55533_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _26911_[0], clk);
  dff _55534_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _26911_[1], clk);
  dff _55535_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _26911_[2], clk);
  dff _55536_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _26911_[3], clk);
  dff _55537_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _26911_[4], clk);
  dff _55538_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _26911_[5], clk);
  dff _55539_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _26911_[6], clk);
  dff _55540_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _26911_[7], clk);
  dff _55541_ (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _26913_[0], clk);
  dff _55542_ (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _26913_[1], clk);
  dff _55543_ (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _26913_[2], clk);
  dff _55544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _22681_, clk);
  dff _55545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _22683_, clk);
  dff _55546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _22682_, clk);
  dff _55547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _22703_, clk);
  dff _55548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _22701_, clk);
  dff _55549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _26992_, clk);
  dff _55550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _11711_, clk);
  dff _55551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _22673_, clk);
  dff _55552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _22880_, clk);
  dff _55553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _22863_, clk);
  dff _55554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _11715_, clk);
  dff _55555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _26978_, clk);
  dff _55556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _22705_, clk);
  dff _55557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _22740_, clk);
  dff _55558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _22727_, clk);
  dff _55559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _22726_, clk);
  dff _55560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _22959_, clk);
  dff _55561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _12237_, clk);
  dff _55562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _23125_, clk);
  dff _55563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _23119_, clk);
  dff _55564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _12234_, clk);
  dff _55565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _11791_, clk);
  dff _55566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _22759_, clk);
  dff _55567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _22758_, clk);
  dff _55568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _12226_, clk);
  dff _55569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _11793_, clk);
  dff _55570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _26942_, clk);
  dff _55571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _23210_, clk);
  dff _55572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _12232_, clk);
  dff _55573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _23297_, clk);
  dff _55574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _12228_, clk);
  dff _55575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _22993_, clk);
  dff _55576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _27008_, clk);
  dff _55577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _22675_, clk);
  dff _55578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _22677_, clk);
  dff _55579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _22676_, clk);
  dff _55580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _12241_, clk);
  dff _55581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _27009_, clk);
  dff _55582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _11867_, clk);
  dff _55583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _22656_, clk);
  dff _55584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _23507_, clk);
  dff _55585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _23513_, clk);
  dff _55586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _12224_, clk);
  dff _55587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _23566_, clk);
  dff _55588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _27301_, clk);
  dff _55589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _23406_, clk);
  dff _55590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _27302_, clk);
  dff _55591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _23388_, clk);
  dff _55592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _04653_, clk);
  dff _55593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _04647_, clk);
  dff _55594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _04638_, clk);
  dff _55595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _27156_, clk);
  dff _55596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _04733_, clk);
  dff _55597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _04716_, clk);
  dff _55598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _22694_, clk);
  dff _55599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _04697_, clk);
  dff _55600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _23723_, clk);
  dff _55601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _27138_, clk);
  dff _55602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _04779_, clk);
  dff _55603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _27139_, clk);
  dff _55604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _22697_, clk);
  dff _55605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _04818_, clk);
  dff _55606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _04847_, clk);
  dff _55607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _27140_, clk);
  dff _55608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _05321_, clk);
  dff _55609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _23410_, clk);
  dff _55610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _05465_, clk);
  dff _55611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _05456_, clk);
  dff _55612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _05451_, clk);
  dff _55613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _05503_, clk);
  dff _55614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _05498_, clk);
  dff _55615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _23650_, clk);
  dff _55616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _27199_, clk);
  dff _55617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _27200_, clk);
  dff _55618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _23685_, clk);
  dff _55619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _10452_, clk);
  dff _55620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _26771_, clk);
  dff _55621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _22715_, clk);
  dff _55622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _23162_, clk);
  dff _55623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _27201_, clk);
  dff _55624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _27196_, clk);
  dff _55625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _27197_, clk);
  dff _55626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _10416_, clk);
  dff _55627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _02571_, clk);
  dff _55628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _03365_, clk);
  dff _55629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _27198_, clk);
  dff _55630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _08203_, clk);
  dff _55631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _06170_, clk);
  dff _55632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _10399_, clk);
  dff _55633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _10737_, clk);
  dff _55634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _10390_, clk);
  dff _55635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _08205_, clk);
  dff _55636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _05707_, clk);
  dff _55637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _10406_, clk);
  dff _55638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _07531_, clk);
  dff _55639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _27195_, clk);
  dff _55640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _12185_, clk);
  dff _55641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _08175_, clk);
  dff _55642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _08442_, clk);
  dff _55643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _11698_, clk);
  dff _55644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _11783_, clk);
  dff _55645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _23426_, clk);
  dff _55646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _10377_, clk);
  dff _55647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _09523_, clk);
  dff _55648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _27193_, clk);
  dff _55649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _10342_, clk);
  dff _55650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _08208_, clk);
  dff _55651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _08909_, clk);
  dff _55652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _27194_, clk);
  dff _55653_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _10355_, clk);
  dff _55654_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _12101_, clk);
  dff _55655_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _12292_, clk);
  dff _55656_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _08210_, clk);
  dff _55657_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _22714_, clk);
  dff _55658_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _22723_, clk);
  dff _55659_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _10336_, clk);
  dff _55660_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _27192_, clk);
  dff _55661_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _18519_, clk);
  dff _55662_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _08749_, clk);
  dff _55663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _08765_, clk);
  dff _55664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _22704_, clk);
  dff _55665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _10310_, clk);
  dff _55666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _27191_, clk);
  dff _55667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _10770_, clk);
  dff _55668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _08179_, clk);
  dff _55669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _01784_, clk);
  dff _55670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _07708_, clk);
  dff _55671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _02210_, clk);
  dff _55672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _27189_, clk);
  dff _55673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _10280_, clk);
  dff _55674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _07185_, clk);
  dff _55675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _27190_, clk);
  dff _55676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _22925_, clk);
  dff _55677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _10297_, clk);
  dff _55678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _07402_, clk);
  dff _55679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _08181_, clk);
  dff _55680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _11617_, clk);
  dff _55681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _10015_, clk);
  dff _55682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _10138_, clk);
  dff _55683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _11458_, clk);
  dff _55684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _10291_, clk);
  dff _55685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _11456_, clk);
  dff _55686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _27188_, clk);
  dff _55687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _11615_, clk);
  dff _55688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _11539_, clk);
  dff _55689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _27186_, clk);
  dff _55690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _09680_, clk);
  dff _55691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _27187_, clk);
  dff _55692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _11463_, clk);
  dff _55693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _09958_, clk);
  dff _55694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _11460_, clk);
  dff _55695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _09981_, clk);
  dff _55696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _09490_, clk);
  dff _55697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _11543_, clk);
  dff _55698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _09519_, clk);
  dff _55699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _11471_, clk);
  dff _55700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _27185_, clk);
  dff _55701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _11541_, clk);
  dff _55702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _09609_, clk);
  dff _55703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _09650_, clk);
  dff _55704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _10349_, clk);
  dff _55705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _10368_, clk);
  dff _55706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _09368_, clk);
  dff _55707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _10100_, clk);
  dff _55708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _10379_, clk);
  dff _55709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _09366_, clk);
  dff _55710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _27297_, clk);
  dff _55711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _10403_, clk);
  dff _55712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _09375_, clk);
  dff _55713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _10287_, clk);
  dff _55714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _10301_, clk);
  dff _55715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _27295_, clk);
  dff _55716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _09373_, clk);
  dff _55717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _27296_, clk);
  dff _55718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _10345_, clk);
  dff _55719_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _09370_, clk);
  dff _55720_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _11258_, clk);
  dff _55721_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _11246_, clk);
  dff _55722_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _27292_, clk);
  dff _55723_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _27293_, clk);
  dff _55724_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _27294_, clk);
  dff _55725_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _11307_, clk);
  dff _55726_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _11331_, clk);
  dff _55727_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _11312_, clk);
  dff _55728_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _27289_, clk);
  dff _55729_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _11134_, clk);
  dff _55730_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _09094_, clk);
  dff _55731_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _27290_, clk);
  dff _55732_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _27291_, clk);
  dff _55733_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _11408_, clk);
  dff _55734_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _11364_, clk);
  dff _55735_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _11388_, clk);
  dff _55736_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _11071_, clk);
  dff _55737_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _08963_, clk);
  dff _55738_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _11077_, clk);
  dff _55739_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _27287_, clk);
  dff _55740_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _08959_, clk);
  dff _55741_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _09202_, clk);
  dff _55742_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _11106_, clk);
  dff _55743_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _27288_, clk);
  dff _55744_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _27282_, clk);
  dff _55745_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _27283_, clk);
  dff _55746_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _08971_, clk);
  dff _55747_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _27284_, clk);
  dff _55748_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _08969_, clk);
  dff _55749_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _27285_, clk);
  dff _55750_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _09110_, clk);
  dff _55751_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _27286_, clk);
  dff _55752_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _09270_, clk);
  dff _55753_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _10973_, clk);
  dff _55754_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _27279_, clk);
  dff _55755_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _08977_, clk);
  dff _55756_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _27280_, clk);
  dff _55757_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _08975_, clk);
  dff _55758_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _27281_, clk);
  dff _55759_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _09114_, clk);
  dff _55760_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _09206_, clk);
  dff _55761_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _10892_, clk);
  dff _55762_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _10915_, clk);
  dff _55763_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _08983_, clk);
  dff _55764_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _10945_, clk);
  dff _55765_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _08981_, clk);
  dff _55766_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _10955_, clk);
  dff _55767_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _09118_, clk);
  dff _55768_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _10055_, clk);
  dff _55769_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _11092_, clk);
  dff _55770_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _12266_, clk);
  dff _55771_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _11193_, clk);
  dff _55772_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _11080_, clk);
  dff _55773_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _12256_, clk);
  dff _55774_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _12243_, clk);
  dff _55775_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _12239_, clk);
  dff _55776_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _10830_, clk);
  dff _55777_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _09014_, clk);
  dff _55778_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _10834_, clk);
  dff _55779_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _10864_, clk);
  dff _55780_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _09011_, clk);
  dff _55781_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _27277_, clk);
  dff _55782_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _09010_, clk);
  dff _55783_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _10876_, clk);
  dff _55784_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _11104_, clk);
  dff _55785_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _11124_, clk);
  dff _55786_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _09945_, clk);
  dff _55787_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _11127_, clk);
  dff _55788_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _11139_, clk);
  dff _55789_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _09274_, clk);
  dff _55790_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _26934_, clk);
  dff _55791_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _26935_, clk);
  dff _55792_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _09954_, clk);
  dff _55793_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _26930_, clk);
  dff _55794_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _09282_, clk);
  dff _55795_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _11057_, clk);
  dff _55796_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _09950_, clk);
  dff _55797_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _26931_, clk);
  dff _55798_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _26932_, clk);
  dff _55799_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _26933_, clk);
  dff _55800_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _09966_, clk);
  dff _55801_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _26924_, clk);
  dff _55802_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _26925_, clk);
  dff _55803_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _09956_, clk);
  dff _55804_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _26926_, clk);
  dff _55805_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _26927_, clk);
  dff _55806_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _26928_, clk);
  dff _55807_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _26929_, clk);
  dff _55808_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _26922_, clk);
  dff _55809_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _09974_, clk);
  dff _55810_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _10928_, clk);
  dff _55811_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _10960_, clk);
  dff _55812_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _09305_, clk);
  dff _55813_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _10083_, clk);
  dff _55814_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _26923_, clk);
  dff _55815_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _09299_, clk);
  dff _55816_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _09022_, clk);
  dff _55817_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _07507_, clk);
  dff _55818_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _07705_, clk);
  dff _55819_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _05661_, clk);
  dff _55820_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _05784_, clk);
  dff _55821_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _07564_, clk);
  dff _55822_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _05659_, clk);
  dff _55823_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _07569_, clk);
  dff _55824_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _07529_, clk);
  dff _55825_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _08162_, clk);
  dff _55826_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _08170_, clk);
  dff _55827_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _07635_, clk);
  dff _55828_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _08172_, clk);
  dff _55829_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _26945_, clk);
  dff _55830_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _07520_, clk);
  dff _55831_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _08965_, clk);
  dff _55832_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _06543_, clk);
  dff _55833_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _06913_, clk);
  dff _55834_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _07644_, clk);
  dff _55835_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _06926_, clk);
  dff _55836_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _07567_, clk);
  dff _55837_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _07532_, clk);
  dff _55838_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _07712_, clk);
  dff _55839_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _07625_, clk);
  dff _55840_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _06562_, clk);
  dff _55841_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _02062_, clk);
  dff _55842_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _06664_, clk);
  dff _55843_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _27161_, clk);
  dff _55844_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _27162_, clk);
  dff _55845_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _27163_, clk);
  dff _55846_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _06368_, clk);
  dff _55847_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _06342_, clk);
  dff _55848_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _25152_, clk);
  dff _55849_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _06784_, clk);
  dff _55850_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _27159_, clk);
  dff _55851_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _06915_, clk);
  dff _55852_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _06891_, clk);
  dff _55853_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _25147_, clk);
  dff _55854_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _25673_, clk);
  dff _55855_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _27160_, clk);
  dff _55856_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _07278_, clk);
  dff _55857_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _07253_, clk);
  dff _55858_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _02013_, clk);
  dff _55859_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _25575_, clk);
  dff _55860_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _06986_, clk);
  dff _55861_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _02033_, clk);
  dff _55862_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _07092_, clk);
  dff _55863_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _07089_, clk);
  dff _55864_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _25747_, clk);
  dff _55865_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _07359_, clk);
  dff _55866_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _07338_, clk);
  dff _55867_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _02008_, clk);
  dff _55868_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _07435_, clk);
  dff _55869_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _02003_, clk);
  dff _55870_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _07191_, clk);
  dff _55871_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _27158_, clk);
  dff _55872_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _01104_, clk);
  dff _55873_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _25458_, clk);
  dff _55874_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _12284_, clk);
  dff _55875_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _01833_, clk);
  dff _55876_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _25457_, clk);
  dff _55877_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _11117_, clk);
  dff _55878_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _27157_, clk);
  dff _55879_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _01837_, clk);
  dff _55880_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _27154_, clk);
  dff _55881_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _01750_, clk);
  dff _55882_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _25758_, clk);
  dff _55883_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _01806_, clk);
  dff _55884_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _06103_, clk);
  dff _55885_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _01789_, clk);
  dff _55886_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _27155_, clk);
  dff _55887_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _01344_, clk);
  dff _55888_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _22698_, clk);
  dff _55889_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _01761_, clk);
  dff _55890_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _10856_, clk);
  dff _55891_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _11267_, clk);
  dff _55892_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _01780_, clk);
  dff _55893_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _27153_, clk);
  dff _55894_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _25492_, clk);
  dff _55895_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _23328_, clk);
  dff _55896_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _27152_, clk);
  dff _55897_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _07658_, clk);
  dff _55898_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _07633_, clk);
  dff _55899_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _07611_, clk);
  dff _55900_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _01991_, clk);
  dff _55901_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _25578_, clk);
  dff _55902_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _25771_, clk);
  dff _55903_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _11834_, clk);
  dff _55904_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _25589_, clk);
  dff _55905_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _07729_, clk);
  dff _55906_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _07719_, clk);
  dff _55907_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _07777_, clk);
  dff _55908_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _07797_, clk);
  dff _55909_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _07781_, clk);
  dff _55910_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _25288_, clk);
  dff _55911_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _07523_, clk);
  dff _55912_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _09038_, clk);
  dff _55913_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _27150_, clk);
  dff _55914_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _27151_, clk);
  dff _55915_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _08103_, clk);
  dff _55916_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _08092_, clk);
  dff _55917_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _01976_, clk);
  dff _55918_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _08429_, clk);
  dff _55919_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _08118_, clk);
  dff _55920_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _09191_, clk);
  dff _55921_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _27149_, clk);
  dff _55922_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _09952_, clk);
  dff _55923_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _09387_, clk);
  dff _55924_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _25295_, clk);
  dff _55925_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _08882_, clk);
  dff _55926_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _08463_, clk);
  dff _55927_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _08458_, clk);
  dff _55928_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _10623_, clk);
  dff _55929_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _25298_, clk);
  dff _55930_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _10147_, clk);
  dff _55931_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _27146_, clk);
  dff _55932_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _27147_, clk);
  dff _55933_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _01946_, clk);
  dff _55934_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _27148_, clk);
  dff _55935_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _09225_, clk);
  dff _55936_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _27239_, clk);
  dff _55937_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _08538_, clk);
  dff _55938_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _27240_, clk);
  dff _55939_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _08931_, clk);
  dff _55940_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _11074_, clk);
  dff _55941_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _26828_, clk);
  dff _55942_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _26769_, clk);
  dff _55943_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _07775_, clk);
  dff _55944_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _25366_, clk);
  dff _55945_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _10982_, clk);
  dff _55946_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _10952_, clk);
  dff _55947_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _01933_, clk);
  dff _55948_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _27145_, clk);
  dff _55949_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _25357_, clk);
  dff _55950_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _10397_, clk);
  dff _55951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _01943_, clk);
  dff _55952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _11863_, clk);
  dff _55953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _27143_, clk);
  dff _55954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _11454_, clk);
  dff _55955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _27144_, clk);
  dff _55956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _11595_, clk);
  dff _55957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _11216_, clk);
  dff _55958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _11207_, clk);
  dff _55959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _11265_, clk);
  dff _55960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _27141_, clk);
  dff _55961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _11964_, clk);
  dff _55962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _12002_, clk);
  dff _55963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _12230_, clk);
  dff _55964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _27142_, clk);
  dff _55965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _01885_, clk);
  dff _55966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _11733_, clk);
  dff _55967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _11724_, clk);
  dff _55968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _27136_, clk);
  dff _55969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _12706_, clk);
  dff _55970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _12704_, clk);
  dff _55971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _01866_, clk);
  dff _55972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _12282_, clk);
  dff _55973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _01881_, clk);
  dff _55974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _27137_, clk);
  dff _55975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _01878_, clk);
  dff _55976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _23300_, clk);
  dff _55977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _27134_, clk);
  dff _55978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _27135_, clk);
  dff _55979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _25440_, clk);
  dff _55980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _12741_, clk);
  dff _55981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _09327_, clk);
  dff _55982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _01860_, clk);
  dff _55983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _25632_, clk);
  dff _55984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _27130_, clk);
  dff _55985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _05849_, clk);
  dff _55986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _03160_, clk);
  dff _55987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _27131_, clk);
  dff _55988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _23620_, clk);
  dff _55989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _27132_, clk);
  dff _55990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _27133_, clk);
  dff _55991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _03439_, clk);
  dff _55992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _06601_, clk);
  dff _55993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _27128_, clk);
  dff _55994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _06642_, clk);
  dff _55995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _03164_, clk);
  dff _55996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _07408_, clk);
  dff _55997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _00995_, clk);
  dff _55998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _27129_, clk);
  dff _55999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _03333_, clk);
  dff _56000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _03346_, clk);
  dff _56001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _27125_, clk);
  dff _56002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _12632_, clk);
  dff _56003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _27126_, clk);
  dff _56004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _04117_, clk);
  dff _56005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _27127_, clk);
  dff _56006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _07203_, clk);
  dff _56007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _03168_, clk);
  dff _56008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _03357_, clk);
  dff _56009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _03441_, clk);
  dff _56010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _22902_, clk);
  dff _56011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _24357_, clk);
  dff _56012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _27123_, clk);
  dff _56013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _23234_, clk);
  dff _56014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _27124_, clk);
  dff _56015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _10574_, clk);
  dff _56016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _27120_, clk);
  dff _56017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _03362_, clk);
  dff _56018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _07744_, clk);
  dff _56019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _22633_, clk);
  dff _56020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _27121_, clk);
  dff _56021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _22756_, clk);
  dff _56022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _27122_, clk);
  dff _56023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _06787_, clk);
  dff _56024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _22691_, clk);
  dff _56025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _07800_, clk);
  dff _56026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _08427_, clk);
  dff _56027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _26642_, clk);
  dff _56028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _26649_, clk);
  dff _56029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _26667_, clk);
  dff _56030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _27237_, clk);
  dff _56031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _27238_, clk);
  dff _56032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _27115_, clk);
  dff _56033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _27116_, clk);
  dff _56034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _27117_, clk);
  dff _56035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _22689_, clk);
  dff _56036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _22688_, clk);
  dff _56037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _27118_, clk);
  dff _56038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _22687_, clk);
  dff _56039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _27119_, clk);
  dff _56040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _02876_, clk);
  dff _56041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _22699_, clk);
  dff _56042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _03222_, clk);
  dff _56043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _22696_, clk);
  dff _56044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _02874_, clk);
  dff _56045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _22695_, clk);
  dff _56046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _03211_, clk);
  dff _56047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _22692_, clk);
  dff _56048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _07282_, clk);
  dff _56049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _27233_, clk);
  dff _56050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _09860_, clk);
  dff _56051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _07820_, clk);
  dff _56052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _11538_, clk);
  dff _56053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _04364_, clk);
  dff _56054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _22641_, clk);
  dff _56055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _23255_, clk);
  dff _56056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _07250_, clk);
  dff _56057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _07011_, clk);
  dff _56058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _07805_, clk);
  dff _56059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _22709_, clk);
  dff _56060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _27235_, clk);
  dff _56061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _22707_, clk);
  dff _56062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _22690_, clk);
  dff _56063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _27236_, clk);
  dff _56064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _03114_, clk);
  dff _56065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _08487_, clk);
  dff _56066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _03294_, clk);
  dff _56067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _03433_, clk);
  dff _56068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _22713_, clk);
  dff _56069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _02882_, clk);
  dff _56070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _22711_, clk);
  dff _56071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _03225_, clk);
  dff _56072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _00203_, clk);
  dff _56073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _03129_, clk);
  dff _56074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _09638_, clk);
  dff _56075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _03139_, clk);
  dff _56076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _10966_, clk);
  dff _56077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _03125_, clk);
  dff _56078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _27114_, clk);
  dff _56079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _03310_, clk);
  dff _56080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _22725_, clk);
  dff _56081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _27111_, clk);
  dff _56082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _27112_, clk);
  dff _56083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _27113_, clk);
  dff _56084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _22720_, clk);
  dff _56085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _03227_, clk);
  dff _56086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _03418_, clk);
  dff _56087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _11998_, clk);
  dff _56088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _01296_, clk);
  dff _56089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _01285_, clk);
  dff _56090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _27227_, clk);
  dff _56091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _01393_, clk);
  dff _56092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _27228_, clk);
  dff _56093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _27229_, clk);
  dff _56094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _08195_, clk);
  dff _56095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _23698_, clk);
  dff _56096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _27230_, clk);
  dff _56097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _23703_, clk);
  dff _56098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _00874_, clk);
  dff _56099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _01020_, clk);
  dff _56100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _00921_, clk);
  dff _56101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _27231_, clk);
  dff _56102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _27232_, clk);
  dff _56103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _10013_, clk);
  dff _56104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _27222_, clk);
  dff _56105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _09002_, clk);
  dff _56106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _09059_, clk);
  dff _56107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _08090_, clk);
  dff _56108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _08432_, clk);
  dff _56109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _08476_, clk);
  dff _56110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _05389_, clk);
  dff _56111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _05306_, clk);
  dff _56112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _27223_, clk);
  dff _56113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _27224_, clk);
  dff _56114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _05639_, clk);
  dff _56115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _10980_, clk);
  dff _56116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _03995_, clk);
  dff _56117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _03969_, clk);
  dff _56118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _03676_, clk);
  dff _56119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _05179_, clk);
  dff _56120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _25585_, clk);
  dff _56121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _12028_, clk);
  dff _56122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _11803_, clk);
  dff _56123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _25487_, clk);
  dff _56124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _25478_, clk);
  dff _56125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _25535_, clk);
  dff _56126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _27082_, clk);
  dff _56127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _11738_, clk);
  dff _56128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _10920_, clk);
  dff _56129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _10895_, clk);
  dff _56130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _08094_, clk);
  dff _56131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _09919_, clk);
  dff _56132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _09906_, clk);
  dff _56133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _09900_, clk);
  dff _56134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _10360_, clk);
  dff _56135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _10938_, clk);
  dff _56136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _26914_, clk);
  dff _56137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _25617_, clk);
  dff _56138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _25614_, clk);
  dff _56139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _12024_, clk);
  dff _56140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _25658_, clk);
  dff _56141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _25648_, clk);
  dff _56142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _11754_, clk);
  dff _56143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _26915_, clk);
  dff _56144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _27203_, clk);
  dff _56145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _24502_, clk);
  dff _56146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _24499_, clk);
  dff _56147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _24496_, clk);
  dff _56148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _12072_, clk);
  dff _56149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _24395_, clk);
  dff _56150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _27204_, clk);
  dff _56151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _24387_, clk);
  dff _56152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _25347_, clk);
  dff _56153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _11734_, clk);
  dff _56154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _24547_, clk);
  dff _56155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _24557_, clk);
  dff _56156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _24551_, clk);
  dff _56157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _12070_, clk);
  dff _56158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _24590_, clk);
  dff _56159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _12068_, clk);
  dff _56160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _25392_, clk);
  dff _56161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _25452_, clk);
  dff _56162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _25436_, clk);
  dff _56163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _12063_, clk);
  dff _56164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _24681_, clk);
  dff _56165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _27172_, clk);
  dff _56166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _24638_, clk);
  dff _56167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _12066_, clk);
  dff _56168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _24205_, clk);
  dff _56169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _11726_, clk);
  dff _56170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _23996_, clk);
  dff _56171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _24002_, clk);
  dff _56172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _23999_, clk);
  dff _56173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _12111_, clk);
  dff _56174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _24099_, clk);
  dff _56175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _24097_, clk);
  dff _56176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _24321_, clk);
  dff _56177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _24314_, clk);
  dff _56178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _12105_, clk);
  dff _56179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _24133_, clk);
  dff _56180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _24183_, clk);
  dff _56181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _27234_, clk);
  dff _56182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _12109_, clk);
  dff _56183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _24202_, clk);
  dff _56184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _24423_, clk);
  dff _56185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _24419_, clk);
  dff _56186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _24413_, clk);
  dff _56187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _24410_, clk);
  dff _56188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _11728_, clk);
  dff _56189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _11849_, clk);
  dff _56190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _24281_, clk);
  dff _56191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _12107_, clk);
  dff _56192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _23826_, clk);
  dff _56193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _23815_, clk);
  dff _56194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _23763_, clk);
  dff _56195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _23931_, clk);
  dff _56196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _23928_, clk);
  dff _56197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _27278_, clk);
  dff _56198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _12116_, clk);
  dff _56199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _11795_, clk);
  dff _56200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _26664_, clk);
  dff _56201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _27108_, clk);
  dff _56202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _02906_, clk);
  dff _56203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _25180_, clk);
  dff _56204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _27109_, clk);
  dff _56205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _25177_, clk);
  dff _56206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _27110_, clk);
  dff _56207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _23176_, clk);
  dff _56208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _26731_, clk);
  dff _56209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _02972_, clk);
  dff _56210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _26726_, clk);
  dff _56211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _03270_, clk);
  dff _56212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _26720_, clk);
  dff _56213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _27107_, clk);
  dff _56214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _02923_, clk);
  dff _56215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _03391_, clk);
  dff _56216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _27106_, clk);
  dff _56217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _26834_, clk);
  dff _56218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _03108_, clk);
  dff _56219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _26805_, clk);
  dff _56220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _03287_, clk);
  dff _56221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _26764_, clk);
  dff _56222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _26748_, clk);
  dff _56223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _03046_, clk);
  dff _56224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _24330_, clk);
  dff _56225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _24580_, clk);
  dff _56226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _05568_, clk);
  dff _56227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _24583_, clk);
  dff _56228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _05573_, clk);
  dff _56229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _05842_, clk);
  dff _56230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _24603_, clk);
  dff _56231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _24609_, clk);
  dff _56232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _05557_, clk);
  dff _56233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _27105_, clk);
  dff _56234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _05625_, clk);
  dff _56235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _05584_, clk);
  dff _56236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _05643_, clk);
  dff _56237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _24571_, clk);
  dff _56238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _24311_, clk);
  dff _56239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _24327_, clk);
  dff _56240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _27103_, clk);
  dff _56241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _05108_, clk);
  dff _56242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _27104_, clk);
  dff _56243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _03936_, clk);
  dff _56244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _05788_, clk);
  dff _56245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _05804_, clk);
  dff _56246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _05754_, clk);
  dff _56247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _05543_, clk);
  dff _56248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _04238_, clk);
  dff _56249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _05010_, clk);
  dff _56250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _05046_, clk);
  dff _56251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _05059_, clk);
  dff _56252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _27102_, clk);
  dff _56253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _05071_, clk);
  dff _56254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _04140_, clk);
  dff _56255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _05078_, clk);
  dff _56256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _04932_, clk);
  dff _56257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _27100_, clk);
  dff _56258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _04954_, clk);
  dff _56259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _27101_, clk);
  dff _56260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _03987_, clk);
  dff _56261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _04990_, clk);
  dff _56262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _03984_, clk);
  dff _56263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _04997_, clk);
  dff _56264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _27097_, clk);
  dff _56265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _27098_, clk);
  dff _56266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _04889_, clk);
  dff _56267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _04174_, clk);
  dff _56268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _04906_, clk);
  dff _56269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _04921_, clk);
  dff _56270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _04171_, clk);
  dff _56271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _04923_, clk);
  dff _56272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _04784_, clk);
  dff _56273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _04195_, clk);
  dff _56274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _04796_, clk);
  dff _56275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _04824_, clk);
  dff _56276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _27096_, clk);
  dff _56277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _04258_, clk);
  dff _56278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _04837_, clk);
  dff _56279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _04868_, clk);
  dff _56280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _04203_, clk);
  dff _56281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _04722_, clk);
  dff _56282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _04731_, clk);
  dff _56283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _04750_, clk);
  dff _56284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _04031_, clk);
  dff _56285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _04755_, clk);
  dff _56286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _04199_, clk);
  dff _56287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _27095_, clk);
  dff _56288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _04422_, clk);
  dff _56289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _04456_, clk);
  dff _56290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _04120_, clk);
  dff _56291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _04664_, clk);
  dff _56292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _04672_, clk);
  dff _56293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _04045_, clk);
  dff _56294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _04692_, clk);
  dff _56295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _04713_, clk);
  dff _56296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _04209_, clk);
  dff _56297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _04345_, clk);
  dff _56298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _04359_, clk);
  dff _56299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _04332_, clk);
  dff _56300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _04133_, clk);
  dff _56301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _04385_, clk);
  dff _56302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _04412_, clk);
  dff _56303_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _04125_, clk);
  dff _56304_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _04217_, clk);
  dff _56305_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _04580_, clk);
  dff _56306_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _04614_, clk);
  dff _56307_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _04214_, clk);
  dff _56308_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _04620_, clk);
  dff _56309_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _27093_, clk);
  dff _56310_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _27094_, clk);
  dff _56311_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _04655_, clk);
  dff _56312_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _04534_, clk);
  dff _56313_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _04098_, clk);
  dff _56314_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _04548_, clk);
  dff _56315_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _27091_, clk);
  dff _56316_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _04553_, clk);
  dff _56317_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _04275_, clk);
  dff _56318_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _27092_, clk);
  dff _56319_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _04573_, clk);
  dff _56320_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _05577_, clk);
  dff _56321_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _04468_, clk);
  dff _56322_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _04114_, clk);
  dff _56323_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _04472_, clk);
  dff _56324_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _04225_, clk);
  dff _56325_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _04489_, clk);
  dff _56326_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _04502_, clk);
  dff _56327_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _27090_, clk);
  dff _56328_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _25522_, clk);
  dff _56329_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _05622_, clk);
  dff _56330_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _25351_, clk);
  dff _56331_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _25344_, clk);
  dff _56332_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _25124_, clk);
  dff _56333_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _25428_, clk);
  dff _56334_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _25424_, clk);
  dff _56335_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _25413_, clk);
  dff _56336_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _24306_, clk);
  dff _56337_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _25567_, clk);
  dff _56338_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _05598_, clk);
  dff _56339_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _25463_, clk);
  dff _56340_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _25471_, clk);
  dff _56341_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _25465_, clk);
  dff _56342_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _05633_, clk);
  dff _56343_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _25513_, clk);
  dff _56344_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _24468_, clk);
  dff _56345_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _05542_, clk);
  dff _56346_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _24278_, clk);
  dff _56347_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _24233_, clk);
  dff _56348_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _24227_, clk);
  dff _56349_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _24398_, clk);
  dff _56350_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _24390_, clk);
  dff _56351_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _24355_, clk);
  dff _56352_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _05769_, clk);
  dff _56353_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _25951_, clk);
  dff _56354_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _25944_, clk);
  dff _56355_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _25999_, clk);
  dff _56356_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _24416_, clk);
  dff _56357_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _24433_, clk);
  dff _56358_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _05549_, clk);
  dff _56359_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _24465_, clk);
  dff _56360_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _25606_, clk);
  dff _56361_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _25600_, clk);
  dff _56362_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _27088_, clk);
  dff _56363_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _25655_, clk);
  dff _56364_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _25643_, clk);
  dff _56365_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _25637_, clk);
  dff _56366_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _27089_, clk);
  dff _56367_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _25819_, clk);
  dff _56368_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _25149_, clk);
  dff _56369_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _25107_, clk);
  dff _56370_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _05115_, clk);
  dff _56371_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _03724_, clk);
  dff _56372_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _25670_, clk);
  dff _56373_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _27087_, clk);
  dff _56374_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _25768_, clk);
  dff _56375_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _25767_, clk);
  dff _56376_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _01277_, clk);
  dff _56377_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _01130_, clk);
  dff _56378_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _05112_, clk);
  dff _56379_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _01396_, clk);
  dff _56380_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _01348_, clk);
  dff _56381_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _03453_, clk);
  dff _56382_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _11483_, clk);
  dff _56383_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _11156_, clk);
  dff _56384_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _05570_, clk);
  dff _56385_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _27086_, clk);
  dff _56386_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _01542_, clk);
  dff _56387_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _01538_, clk);
  dff _56388_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _05106_, clk);
  dff _56389_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _03524_, clk);
  dff _56390_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _03448_, clk);
  dff _56391_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _05103_, clk);
  dff _56392_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _05854_, clk);
  dff _56393_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _05076_, clk);
  dff _56394_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _09331_, clk);
  dff _56395_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _09061_, clk);
  dff _56396_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _27085_, clk);
  dff _56397_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _05225_, clk);
  dff _56398_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _04419_, clk);
  dff _56399_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _04379_, clk);
  dff _56400_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _05043_, clk);
  dff _56401_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _10021_, clk);
  dff _56402_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _05062_, clk);
  dff _56403_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _10606_, clk);
  dff _56404_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _27084_, clk);
  dff _56405_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _05056_, clk);
  dff _56406_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _06131_, clk);
  dff _56407_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _05905_, clk);
  dff _56408_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _11568_, clk);
  dff _56409_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _11755_, clk);
  dff _56410_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _05015_, clk);
  dff _56411_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _10975_, clk);
  dff _56412_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _27083_, clk);
  dff _56413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _10930_, clk);
  dff _56414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _05051_, clk);
  dff _56415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _11100_, clk);
  dff _56416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _22642_, clk);
  dff _56417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _22708_, clk);
  dff _56418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _22898_, clk);
  dff _56419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _05004_, clk);
  dff _56420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _03742_, clk);
  dff _56421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _11396_, clk);
  dff _56422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _11358_, clk);
  dff _56423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _11280_, clk);
  dff _56424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _03605_, clk);
  dff _56425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _23207_, clk);
  dff _56426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _22998_, clk);
  dff _56427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _22719_, clk);
  dff _56428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _04988_, clk);
  dff _56429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _12674_, clk);
  dff _56430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _12615_, clk);
  dff _56431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _12543_, clk);
  dff _56432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _25454_, clk);
  dff _56433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _25732_, clk);
  dff _56434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _04975_, clk);
  dff _56435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _27078_, clk);
  dff _56436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _01521_, clk);
  dff _56437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _04971_, clk);
  dff _56438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _03748_, clk);
  dff _56439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _27079_, clk);
  dff _56440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _03505_, clk);
  dff _56441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _27077_, clk);
  dff _56442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _02348_, clk);
  dff _56443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _02338_, clk);
  dff _56444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _04963_, clk);
  dff _56445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _04687_, clk);
  dff _56446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _04592_, clk);
  dff _56447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _03894_, clk);
  dff _56448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _09258_, clk);
  dff _56449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _27076_, clk);
  dff _56450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _03509_, clk);
  dff _56451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _07086_, clk);
  dff _56452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _05964_, clk);
  dff _56453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _04951_, clk);
  dff _56454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _08939_, clk);
  dff _56455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _07688_, clk);
  dff _56456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _09652_, clk);
  dff _56457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _09626_, clk);
  dff _56458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _09737_, clk);
  dff _56459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _09731_, clk);
  dff _56460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _04916_, clk);
  dff _56461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _09049_, clk);
  dff _56462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _09047_, clk);
  dff _56463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _04930_, clk);
  dff _56464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _03846_, clk);
  dff _56465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _27075_, clk);
  dff _56466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _09839_, clk);
  dff _56467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _09818_, clk);
  dff _56468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _10947_, clk);
  dff _56469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _10810_, clk);
  dff _56470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _10710_, clk);
  dff _56471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _03518_, clk);
  dff _56472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _27071_, clk);
  dff _56473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _27072_, clk);
  dff _56474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _04875_, clk);
  dff _56475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _11515_, clk);
  dff _56476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _11400_, clk);
  dff _56477_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _11270_, clk);
  dff _56478_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _27073_, clk);
  dff _56479_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _27074_, clk);
  dff _56480_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _04841_, clk);
  dff _56481_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _27069_, clk);
  dff _56482_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _22702_, clk);
  dff _56483_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _04870_, clk);
  dff _56484_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _02098_, clk);
  dff _56485_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _04865_, clk);
  dff _56486_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _03763_, clk);
  dff _56487_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _27070_, clk);
  dff _56488_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _09823_, clk);
  dff _56489_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _03557_, clk);
  dff _56490_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _03849_, clk);
  dff _56491_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _02539_, clk);
  dff _56492_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _04912_, clk);
  dff _56493_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _03304_, clk);
  dff _56494_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _04844_, clk);
  dff _56495_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _05479_, clk);
  dff _56496_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _11659_, clk);
  dff _56497_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _23189_, clk);
  dff _56498_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _04798_, clk);
  dff _56499_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _08215_, clk);
  dff _56500_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _08951_, clk);
  dff _56501_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _08947_, clk);
  dff _56502_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _04827_, clk);
  dff _56503_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _10206_, clk);
  dff _56504_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _27068_, clk);
  dff _56505_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _08826_, clk);
  dff _56506_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _08828_, clk);
  dff _56507_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _03574_, clk);
  dff _56508_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _12509_, clk);
  dff _56509_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _19972_, clk);
  dff _56510_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _12613_, clk);
  dff _56511_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _04803_, clk);
  dff _56512_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _08771_, clk);
  dff _56513_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _22710_, clk);
  dff _56514_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _22761_, clk);
  dff _56515_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _08522_, clk);
  dff _56516_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _08526_, clk);
  dff _56517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _03577_, clk);
  dff _56518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _09140_, clk);
  dff _56519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _27067_, clk);
  dff _56520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _09681_, clk);
  dff _56521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _07741_, clk);
  dff _56522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _00562_, clk);
  dff _56523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _23819_, clk);
  dff _56524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _04759_, clk);
  dff _56525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _03768_, clk);
  dff _56526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _08773_, clk);
  dff _56527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _08740_, clk);
  dff _56528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _27066_, clk);
  dff _56529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _03209_, clk);
  dff _56530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _26068_, clk);
  dff _56531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _05423_, clk);
  dff _56532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _04753_, clk);
  dff _56533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _22916_, clk);
  dff _56534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _04747_, clk);
  dff _56535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _26706_, clk);
  dff _56536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _04902_, clk);
  dff _56537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _03539_, clk);
  dff _56538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _07818_, clk);
  dff _56539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _06925_, clk);
  dff _56540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _07244_, clk);
  dff _56541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _27065_, clk);
  dff _56542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _09421_, clk);
  dff _56543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _24298_, clk);
  dff _56544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _27275_, clk);
  dff _56545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _10679_, clk);
  dff _56546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _27276_, clk);
  dff _56547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _09025_, clk);
  dff _56548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _10735_, clk);
  dff _56549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _10750_, clk);
  dff _56550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _10791_, clk);
  dff _56551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _09018_, clk);
  dff _56552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _10157_, clk);
  dff _56553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _09219_, clk);
  dff _56554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _10201_, clk);
  dff _56555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _10225_, clk);
  dff _56556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _10253_, clk);
  dff _56557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _09086_, clk);
  dff _56558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _10260_, clk);
  dff _56559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _09179_, clk);
  dff _56560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _10436_, clk);
  dff _56561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _27271_, clk);
  dff _56562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _09172_, clk);
  dff _56563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _10559_, clk);
  dff _56564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _27272_, clk);
  dff _56565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _10179_, clk);
  dff _56566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _27273_, clk);
  dff _56567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _27274_, clk);
  dff _56568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _09071_, clk);
  dff _56569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _09215_, clk);
  dff _56570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _10375_, clk);
  dff _56571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _10395_, clk);
  dff _56572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _09174_, clk);
  dff _56573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _10401_, clk);
  dff _56574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _10413_, clk);
  dff _56575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _09035_, clk);
  dff _56576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _10308_, clk);
  dff _56577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _09079_, clk);
  dff _56578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _10314_, clk);
  dff _56579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _27269_, clk);
  dff _56580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _10346_, clk);
  dff _56581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _09075_, clk);
  dff _56582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _27270_, clk);
  dff _56583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _09074_, clk);
  dff _56584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _11341_, clk);
  dff _56585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _27265_, clk);
  dff _56586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _27266_, clk);
  dff _56587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _27267_, clk);
  dff _56588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _11299_, clk);
  dff _56589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _22757_, clk);
  dff _56590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _27268_, clk);
  dff _56591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _10293_, clk);
  dff _56592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _27258_, clk);
  dff _56593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _27259_, clk);
  dff _56594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _27260_, clk);
  dff _56595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _27261_, clk);
  dff _56596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _27262_, clk);
  dff _56597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _11322_, clk);
  dff _56598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _27263_, clk);
  dff _56599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _27264_, clk);
  dff _56600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _27254_, clk);
  dff _56601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _03117_, clk);
  dff _56602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _12009_, clk);
  dff _56603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _11273_, clk);
  dff _56604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _07690_, clk);
  dff _56605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _27255_, clk);
  dff _56606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _27256_, clk);
  dff _56607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _27257_, clk);
  dff _56608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _27252_, clk);
  dff _56609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _11262_, clk);
  dff _56610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _16236_, clk);
  dff _56611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _22627_, clk);
  dff _56612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _16455_, clk);
  dff _56613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _11244_, clk);
  dff _56614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _27253_, clk);
  dff _56615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _22660_, clk);
  dff _56616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _11356_, clk);
  dff _56617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _03855_, clk);
  dff _56618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _03788_, clk);
  dff _56619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _11394_, clk);
  dff _56620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _04742_, clk);
  dff _56621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _04519_, clk);
  dff _56622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _27251_, clk);
  dff _56623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _05258_, clk);
  dff _56624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _02903_, clk);
  dff _56625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _11353_, clk);
  dff _56626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _27247_, clk);
  dff _56627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _27248_, clk);
  dff _56628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _11418_, clk);
  dff _56629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _27249_, clk);
  dff _56630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _27250_, clk);
  dff _56631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _01716_, clk);
  dff _56632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _11189_, clk);
  dff _56633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _11183_, clk);
  dff _56634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _11136_, clk);
  dff _56635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _08190_, clk);
  dff _56636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _27246_, clk);
  dff _56637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _02437_, clk);
  dff _56638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _11404_, clk);
  dff _56639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _03083_, clk);
  dff _56640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _11255_, clk);
  dff _56641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _27243_, clk);
  dff _56642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _11132_, clk);
  dff _56643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _11368_, clk);
  dff _56644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _27244_, clk);
  dff _56645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _07746_, clk);
  dff _56646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _27245_, clk);
  dff _56647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _04080_, clk);
  dff _56648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _27241_, clk);
  dff _56649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _07752_, clk);
  dff _56650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _11489_, clk);
  dff _56651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _11473_, clk);
  dff _56652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _27242_, clk);
  dff _56653_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _11591_, clk);
  dff _56654_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _11534_, clk);
  dff _56655_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _07750_, clk);
  dff _56656_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _11102_, clk);
  dff _56657_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _22724_, clk);
  dff _56658_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _22693_, clk);
  dff _56659_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _07771_, clk);
  dff _56660_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _11721_, clk);
  dff _56661_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _11718_, clk);
  dff _56662_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _11696_, clk);
  dff _56663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _11853_, clk);
  dff _56664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _04610_, clk);
  dff _56665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _23554_, clk);
  dff _56666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _09433_, clk);
  dff _56667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _27205_, clk);
  dff _56668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _08496_, clk);
  dff _56669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _04849_, clk);
  dff _56670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _10227_, clk);
  dff _56671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _22679_, clk);
  dff _56672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _09156_, clk);
  dff _56673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _11548_, clk);
  dff _56674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _27182_, clk);
  dff _56675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _27183_, clk);
  dff _56676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _27184_, clk);
  dff _56677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _09277_, clk);
  dff _56678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _11545_, clk);
  dff _56679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _09338_, clk);
  dff _56680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _10196_, clk);
  dff _56681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _07300_, clk);
  dff _56682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _08188_, clk);
  dff _56683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _22716_, clk);
  dff _56684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _18188_, clk);
  dff _56685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _10165_, clk);
  dff _56686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _09887_, clk);
  dff _56687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _10163_, clk);
  dff _56688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _27179_, clk);
  dff _56689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _08852_, clk);
  dff _56690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _27180_, clk);
  dff _56691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _08908_, clk);
  dff _56692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _11478_, clk);
  dff _56693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _09009_, clk);
  dff _56694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _27181_, clk);
  dff _56695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _09081_, clk);
  dff _56696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _10646_, clk);
  dff _56697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _11694_, clk);
  dff _56698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _11526_, clk);
  dff _56699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _11425_, clk);
  dff _56700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _08115_, clk);
  dff _56701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _10182_, clk);
  dff _56702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _09184_, clk);
  dff _56703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _27202_, clk);
  dff _56704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _08572_, clk);
  dff _56705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _27177_, clk);
  dff _56706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _11487_, clk);
  dff _56707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _11621_, clk);
  dff _56708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _27178_, clk);
  dff _56709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _11485_, clk);
  dff _56710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _08777_, clk);
  dff _56711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _11562_, clk);
  dff _56712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _08202_, clk);
  dff _56713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _11924_, clk);
  dff _56714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _11911_, clk);
  dff _56715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _12273_, clk);
  dff _56716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _12294_, clk);
  dff _56717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _12277_, clk);
  dff _56718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _11230_, clk);
  dff _56719_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _11153_, clk);
  dff _56720_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _11569_, clk);
  dff _56721_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _08365_, clk);
  dff _56722_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _08416_, clk);
  dff _56723_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _11493_, clk);
  dff _56724_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _11622_, clk);
  dff _56725_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _08466_, clk);
  dff _56726_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _08544_, clk);
  dff _56727_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _11491_, clk);
  dff _56728_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _06542_, clk);
  dff _56729_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _11613_, clk);
  dff _56730_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _06585_, clk);
  dff _56731_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _27175_, clk);
  dff _56732_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _11532_, clk);
  dff _56733_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _11628_, clk);
  dff _56734_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _08161_, clk);
  dff _56735_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _27176_, clk);
  dff _56736_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _07925_, clk);
  dff _56737_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _11505_, clk);
  dff _56738_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _11625_, clk);
  dff _56739_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _07944_, clk);
  dff _56740_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _08032_, clk);
  dff _56741_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _11502_, clk);
  dff _56742_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _08086_, clk);
  dff _56743_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _08131_, clk);
  dff _56744_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _27173_, clk);
  dff _56745_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _07490_, clk);
  dff _56746_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _11510_, clk);
  dff _56747_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _27174_, clk);
  dff _56748_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _07528_, clk);
  dff _56749_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _07737_, clk);
  dff _56750_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _11506_, clk);
  dff _56751_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _07894_, clk);
  dff _56752_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _11524_, clk);
  dff _56753_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _06977_, clk);
  dff _56754_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _11522_, clk);
  dff _56755_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _07034_, clk);
  dff _56756_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _11609_, clk);
  dff _56757_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _07208_, clk);
  dff _56758_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _11519_, clk);
  dff _56759_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _27171_, clk);
  dff _56760_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _06777_, clk);
  dff _56761_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _04899_, clk);
  dff _56762_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _04933_, clk);
  dff _56763_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _04960_, clk);
  dff _56764_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _23319_, clk);
  dff _56765_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _27169_, clk);
  dff _56766_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _27170_, clk);
  dff _56767_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _11528_, clk);
  dff _56768_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _22774_, clk);
  dff _56769_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _22671_, clk);
  dff _56770_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _00828_, clk);
  dff _56771_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _04699_, clk);
  dff _56772_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _27166_, clk);
  dff _56773_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _27167_, clk);
  dff _56774_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _04910_, clk);
  dff _56775_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _27168_, clk);
  dff _56776_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _27165_, clk);
  dff _56777_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _12113_, clk);
  dff _56778_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _04999_, clk);
  dff _56779_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _04986_, clk);
  dff _56780_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _22659_, clk);
  dff _56781_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _05082_, clk);
  dff _56782_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _05069_, clk);
  dff _56783_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _05048_, clk);
  dff _56784_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _27164_, clk);
  dff _56785_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _05232_, clk);
  dff _56786_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _05155_, clk);
  dff _56787_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _05150_, clk);
  dff _56788_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _05136_, clk);
  dff _56789_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _05123_, clk);
  dff _56790_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _05202_, clk);
  dff _56791_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _05198_, clk);
  dff _56792_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _27033_, clk);
  dff _56793_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _21247_, clk);
  dff _56794_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _21419_, clk);
  dff _56795_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _21348_, clk);
  dff _56796_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _27034_, clk);
  dff _56797_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _22629_, clk);
  dff _56798_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _22542_, clk);
  dff _56799_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _12247_, clk);
  dff _56800_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _05418_, clk);
  dff _56801_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _05408_, clk);
  dff _56802_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _23659_, clk);
  dff _56803_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _05287_, clk);
  dff _56804_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _05280_, clk);
  dff _56805_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _05274_, clk);
  dff _56806_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _27099_, clk);
  dff _56807_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _05341_, clk);
  dff _56808_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _27300_, clk);
  dff _56809_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _10110_, clk);
  dff _56810_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _10197_, clk);
  dff _56811_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _10231_, clk);
  dff _56812_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _09384_, clk);
  dff _56813_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _10240_, clk);
  dff _56814_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _09379_, clk);
  dff _56815_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _10258_, clk);
  dff _56816_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _22640_, clk);
  dff _56817_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _22637_, clk);
  dff _56818_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _22658_, clk);
  dff _56819_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _04530_, clk);
  dff _56820_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _27041_, clk);
  dff _56821_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _21820_, clk);
  dff _56822_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _04550_, clk);
  dff _56823_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _04542_, clk);
  dff _56824_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _27042_, clk);
  dff _56825_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _04562_, clk);
  dff _56826_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _20570_, clk);
  dff _56827_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _03664_, clk);
  dff _56828_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _03871_, clk);
  dff _56829_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _12920_, clk);
  dff _56830_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _12950_, clk);
  dff _56831_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _15784_, clk);
  dff _56832_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _06171_, clk);
  dff _56833_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _27020_, clk);
  dff _56834_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _26054_, clk);
  dff _56835_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _26057_, clk);
  dff _56836_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _27021_, clk);
  dff _56837_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _26059_, clk);
  dff _56838_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _26066_, clk);
  dff _56839_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _06100_, clk);
  dff _56840_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _26981_, clk);
  dff _56841_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _26982_, clk);
  dff _56842_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _06660_, clk);
  dff _56843_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _26983_, clk);
  dff _56844_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _10194_, clk);
  dff _56845_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _26984_, clk);
  dff _56846_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _10304_, clk);
  dff _56847_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _10289_, clk);
  dff _56848_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _09382_, clk);
  dff _56849_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _09309_, clk);
  dff _56850_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _09296_, clk);
  dff _56851_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _10104_, clk);
  dff _56852_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _10036_, clk);
  dff _56853_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _09991_, clk);
  dff _56854_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _06864_, clk);
  dff _56855_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _09101_, clk);
  dff _56856_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _11164_, clk);
  dff _56857_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _05546_, clk);
  dff _56858_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _09837_, clk);
  dff _56859_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _09359_, clk);
  dff _56860_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _06705_, clk);
  dff _56861_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _06611_, clk);
  dff _56862_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _01901_, clk);
  dff _56863_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _26980_, clk);
  dff _56864_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _11161_, clk);
  dff _56865_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _01372_, clk);
  dff _56866_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _06709_, clk);
  dff _56867_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _06528_, clk);
  dff _56868_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _22835_, clk);
  dff _56869_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _06714_, clk);
  dff _56870_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _06711_, clk);
  dff _56871_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _26962_, clk);
  dff _56872_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _27298_, clk);
  dff _56873_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _10454_, clk);
  dff _56874_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _10511_, clk);
  dff _56875_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _10569_, clk);
  dff _56876_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _10625_, clk);
  dff _56877_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _09357_, clk);
  dff _56878_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _10172_, clk);
  dff _56879_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _27299_, clk);
  dff _56880_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _04409_, clk);
  dff _56881_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _07854_, clk);
  dff _56882_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _01524_, clk);
  dff _56883_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _01495_, clk);
  dff _56884_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _27225_, clk);
  dff _56885_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _02826_, clk);
  dff _56886_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _02446_, clk);
  dff _56887_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _27226_, clk);
  dff _56888_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _27219_, clk);
  dff _56889_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _27220_, clk);
  dff _56890_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _27221_, clk);
  dff _56891_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _11203_, clk);
  dff _56892_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _11200_, clk);
  dff _56893_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _10897_, clk);
  dff _56894_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _10784_, clk);
  dff _56895_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _10799_, clk);
  dff _56896_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _11236_, clk);
  dff _56897_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _11228_, clk);
  dff _56898_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _27217_, clk);
  dff _56899_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _11497_, clk);
  dff _56900_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _11468_, clk);
  dff _56901_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _08107_, clk);
  dff _56902_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _08435_, clk);
  dff _56903_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _27218_, clk);
  dff _56904_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _10813_, clk);
  dff _56905_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _04851_, clk);
  dff _56906_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _27214_, clk);
  dff _56907_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _09923_, clk);
  dff _56908_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _02714_, clk);
  dff _56909_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _22685_, clk);
  dff _56910_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _22684_, clk);
  dff _56911_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _22670_, clk);
  dff _56912_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _12477_, clk);
  dff _56913_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _12288_, clk);
  dff _56914_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _11882_, clk);
  dff _56915_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _27215_, clk);
  dff _56916_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _12586_, clk);
  dff _56917_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _12545_, clk);
  dff _56918_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _27216_, clk);
  dff _56919_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _11222_, clk);
  dff _56920_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _10838_, clk);
  dff _56921_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _25628_, clk);
  dff _56922_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _26780_, clk);
  dff _56923_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _22639_, clk);
  dff _56924_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _19920_, clk);
  dff _56925_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _22636_, clk);
  dff _56926_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _22638_, clk);
  dff _56927_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _08110_, clk);
  dff _56928_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _27209_, clk);
  dff _56929_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _08439_, clk);
  dff _56930_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _05185_, clk);
  dff _56931_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _05689_, clk);
  dff _56932_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _05300_, clk);
  dff _56933_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _07535_, clk);
  dff _56934_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _07290_, clk);
  dff _56935_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _10755_, clk);
  dff _56936_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _27213_, clk);
  dff _56937_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _01820_, clk);
  dff _56938_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _01566_, clk);
  dff _56939_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _24697_, clk);
  dff _56940_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _24449_, clk);
  dff _56941_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _10832_, clk);
  dff _56942_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _25792_, clk);
  dff _56943_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _25972_, clk);
  dff _56944_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _27210_, clk);
  dff _56945_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _02362_, clk);
  dff _56946_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _10797_, clk);
  dff _56947_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _27211_, clk);
  dff _56948_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _04640_, clk);
  dff _56949_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _10780_, clk);
  dff _56950_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _27212_, clk);
  dff _56951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _00764_, clk);
  dff _56952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _10748_, clk);
  dff _56953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _10650_, clk);
  dff _56954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _27206_, clk);
  dff _56955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _09668_, clk);
  dff _56956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _10706_, clk);
  dff _56957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _09753_, clk);
  dff _56958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _09733_, clk);
  dff _56959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _27207_, clk);
  dff _56960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _09254_, clk);
  dff _56961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _10731_, clk);
  dff _56962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _09612_, clk);
  dff _56963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _09600_, clk);
  dff _56964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _27208_, clk);
  dff _56965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _08995_, clk);
  dff _56966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _08943_, clk);
  dff _56967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _10745_, clk);
  dff _56968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _05902_, clk);
  dff _56969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _05673_, clk);
  dff _56970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _05587_, clk);
  dff _56971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _10652_, clk);
  dff _56972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _10604_, clk);
  dff _56973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _12268_, clk);
  dff _56974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _05386_, clk);
  dff _56975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _05370_, clk);
  dff _56976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _27080_, clk);
  dff _56977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _12258_, clk);
  dff _56978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _11091_, clk);
  dff _56979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _11051_, clk);
  dff _56980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _27081_, clk);
  dff _56981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _12264_, clk);
  dff _56982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _11792_, clk);
  dff _56983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _11681_, clk);
  dff _56984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _17981_, clk);
  dff _56985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _18303_, clk);
  dff _56986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _12252_, clk);
  dff _56987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _19421_, clk);
  dff _56988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _20043_, clk);
  dff _56989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _27058_, clk);
  dff _56990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _11787_, clk);
  dff _56991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _14938_, clk);
  dff _56992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _14601_, clk);
  dff _56993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _14450_, clk);
  dff _56994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _17417_, clk);
  dff _56995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _17267_, clk);
  dff _56996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _12254_, clk);
  dff _56997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _12344_, clk);
  dff _56998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _12223_, clk);
  dff _56999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _12805_, clk);
  dff _57000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _22661_, clk);
  dff _57001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _22669_, clk);
  dff _57002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _22662_, clk);
  dff _57003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _11707_, clk);
  dff _57004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _22632_, clk);
  dff _57005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _22631_, clk);
  dff _57006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _12245_, clk);
  dff _57007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _22635_, clk);
  dff _57008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _04802_, clk);
  dff _57009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _04719_, clk);
  dff _57010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _08089_, clk);
  dff _57011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _04710_, clk);
  dff _57012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _03792_, clk);
  dff _57013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _05383_, clk);
  dff _57014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _22787_, clk);
  dff _57015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _22678_, clk);
  dff _57016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _03880_, clk);
  dff _57017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _22722_, clk);
  dff _57018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _22643_, clk);
  dff _57019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _27063_, clk);
  dff _57020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _27064_, clk);
  dff _57021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _07342_, clk);
  dff _57022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _05815_, clk);
  dff _57023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _04689_, clk);
  dff _57024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _13798_, clk);
  dff _57025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _04670_, clk);
  dff _57026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _22628_, clk);
  dff _57027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _17600_, clk);
  dff _57028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _24247_, clk);
  dff _57029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _19941_, clk);
  dff _57030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _10888_, clk);
  dff _57031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _03613_, clk);
  dff _57032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _23504_, clk);
  dff _57033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _03703_, clk);
  dff _57034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _27060_, clk);
  dff _57035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _04446_, clk);
  dff _57036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _03701_, clk);
  dff _57037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _23248_, clk);
  dff _57038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _27061_, clk);
  dff _57039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _27062_, clk);
  dff _57040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _27050_, clk);
  dff _57041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _27051_, clk);
  dff _57042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _27052_, clk);
  dff _57043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _27053_, clk);
  dff _57044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _27054_, clk);
  dff _57045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _27055_, clk);
  dff _57046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _04651_, clk);
  dff _57047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _03802_, clk);
  dff _57048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _24200_, clk);
  dff _57049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _04330_, clk);
  dff _57050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _03883_, clk);
  dff _57051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _04400_, clk);
  dff _57052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _23586_, clk);
  dff _57053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _27059_, clk);
  dff _57054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _23477_, clk);
  dff _57055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _23517_, clk);
  dff _57056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _04352_, clk);
  dff _57057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _24091_, clk);
  dff _57058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _27056_, clk);
  dff _57059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _04382_, clk);
  dff _57060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _23891_, clk);
  dff _57061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _03713_, clk);
  dff _57062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _27057_, clk);
  dff _57063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _24106_, clk);
  dff _57064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _03542_, clk);
  dff _57065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _27046_, clk);
  dff _57066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _27047_, clk);
  dff _57067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _27048_, clk);
  dff _57068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _27049_, clk);
  dff _57069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _04645_, clk);
  dff _57070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _02060_, clk);
  dff _57071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _01953_, clk);
  dff _57072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _04361_, clk);
  dff _57073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _04416_, clk);
  dff _57074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _04626_, clk);
  dff _57075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _27045_, clk);
  dff _57076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _05825_, clk);
  dff _57077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _03638_, clk);
  dff _57078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _02867_, clk);
  dff _57079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _02582_, clk);
  dff _57080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _04583_, clk);
  dff _57081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _08380_, clk);
  dff _57082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _08049_, clk);
  dff _57083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _07629_, clk);
  dff _57084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _04617_, clk);
  dff _57085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _09056_, clk);
  dff _57086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _09393_, clk);
  dff _57087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _04597_, clk);
  dff _57088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _22700_, clk);
  dff _57089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _04503_, clk);
  dff _57090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _27038_, clk);
  dff _57091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _22672_, clk);
  dff _57092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _27039_, clk);
  dff _57093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _27040_, clk);
  dff _57094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _22674_, clk);
  dff _57095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _04512_, clk);
  dff _57096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _03656_, clk);
  dff _57097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _11987_, clk);
  dff _57098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _04577_, clk);
  dff _57099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _27043_, clk);
  dff _57100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _27044_, clk);
  dff _57101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _03809_, clk);
  dff _57102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _10628_, clk);
  dff _57103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _04587_, clk);
  dff _57104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _03341_, clk);
  dff _57105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _06116_, clk);
  dff _57106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _25580_, clk);
  dff _57107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _23037_, clk);
  dff _57108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _23136_, clk);
  dff _57109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _27031_, clk);
  dff _57110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _27032_, clk);
  dff _57111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _22818_, clk);
  dff _57112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _22936_, clk);
  dff _57113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _27035_, clk);
  dff _57114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _22718_, clk);
  dff _57115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _22717_, clk);
  dff _57116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _27036_, clk);
  dff _57117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _22754_, clk);
  dff _57118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _04492_, clk);
  dff _57119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _27037_, clk);
  dff _57120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _03282_, clk);
  dff _57121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _03289_, clk);
  dff _57122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _27027_, clk);
  dff _57123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _27028_, clk);
  dff _57124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _03291_, clk);
  dff _57125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _03326_, clk);
  dff _57126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _27029_, clk);
  dff _57127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _27030_, clk);
  dff _57128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _03231_, clk);
  dff _57129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _05915_, clk);
  dff _57130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _03233_, clk);
  dff _57131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _06123_, clk);
  dff _57132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _06289_, clk);
  dff _57133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _03244_, clk);
  dff _57134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _27026_, clk);
  dff _57135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _05907_, clk);
  dff _57136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _05968_, clk);
  dff _57137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _03175_, clk);
  dff _57138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _05956_, clk);
  dff _57139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _03177_, clk);
  dff _57140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _06134_, clk);
  dff _57141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _03194_, clk);
  dff _57142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _05949_, clk);
  dff _57143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _03199_, clk);
  dff _57144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _02893_, clk);
  dff _57145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _02908_, clk);
  dff _57146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _05995_, clk);
  dff _57147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _02911_, clk);
  dff _57148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _27024_, clk);
  dff _57149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _05987_, clk);
  dff _57150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _06257_, clk);
  dff _57151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _02996_, clk);
  dff _57152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _03052_, clk);
  dff _57153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _06151_, clk);
  dff _57154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _03069_, clk);
  dff _57155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _03123_, clk);
  dff _57156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _27025_, clk);
  dff _57157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _06254_, clk);
  dff _57158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _03144_, clk);
  dff _57159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _05974_, clk);
  dff _57160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _06163_, clk);
  dff _57161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _01694_, clk);
  dff _57162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _06016_, clk);
  dff _57163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _01696_, clk);
  dff _57164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _27023_, clk);
  dff _57165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _02844_, clk);
  dff _57166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _02880_, clk);
  dff _57167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _06009_, clk);
  dff _57168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _00090_, clk);
  dff _57169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _00200_, clk);
  dff _57170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _27018_, clk);
  dff _57171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _06273_, clk);
  dff _57172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _00206_, clk);
  dff _57173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _00269_, clk);
  dff _57174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _06051_, clk);
  dff _57175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _00275_, clk);
  dff _57176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _26050_, clk);
  dff _57177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _06112_, clk);
  dff _57178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _00617_, clk);
  dff _57179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _06023_, clk);
  dff _57180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _00626_, clk);
  dff _57181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _06168_, clk);
  dff _57182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _27022_, clk);
  dff _57183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _01690_, clk);
  dff _57184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _00279_, clk);
  dff _57185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _06184_, clk);
  dff _57186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _00296_, clk);
  dff _57187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _27019_, clk);
  dff _57188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _00299_, clk);
  dff _57189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _06180_, clk);
  dff _57190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _00309_, clk);
  dff _57191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _00385_, clk);
  dff _57192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _06205_, clk);
  dff _57193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _26081_, clk);
  dff _57194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _26087_, clk);
  dff _57195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _06085_, clk);
  dff _57196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _06276_, clk);
  dff _57197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _26093_, clk);
  dff _57198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _26132_, clk);
  dff _57199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _06077_, clk);
  dff _57200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _27015_, clk);
  dff _57201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _04025_, clk);
  dff _57202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _27016_, clk);
  dff _57203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _07425_, clk);
  dff _57204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _03751_, clk);
  dff _57205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _07416_, clk);
  dff _57206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _26071_, clk);
  dff _57207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _27017_, clk);
  dff _57208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _03436_, clk);
  dff _57209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _03608_, clk);
  dff _57210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _27013_, clk);
  dff _57211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _07055_, clk);
  dff _57212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _26025_, clk);
  dff _57213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _27014_, clk);
  dff _57214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _03398_, clk);
  dff _57215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _03371_, clk);
  dff _57216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _03710_, clk);
  dff _57217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _03683_, clk);
  dff _57218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _03680_, clk);
  dff _57219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _07053_, clk);
  dff _57220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _03775_, clk);
  dff _57221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _03765_, clk);
  dff _57222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _06332_, clk);
  dff _57223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _03463_, clk);
  dff _57224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _06446_, clk);
  dff _57225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _06470_, clk);
  dff _57226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _02068_, clk);
  dff _57227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _25569_, clk);
  dff _57228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _06141_, clk);
  dff _57229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _06178_, clk);
  dff _57230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _06160_, clk);
  dff _57231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _02085_, clk);
  dff _57232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _04193_, clk);
  dff _57233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _04212_, clk);
  dff _57234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _06338_, clk);
  dff _57235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _03878_, clk);
  dff _57236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _03865_, clk);
  dff _57237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _04007_, clk);
  dff _57238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _04003_, clk);
  dff _57239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _03980_, clk);
  dff _57240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _04270_, clk);
  dff _57241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _27012_, clk);
  dff _57242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _04371_, clk);
  dff _57243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _04355_, clk);
  dff _57244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _06360_, clk);
  dff _57245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _04049_, clk);
  dff _57246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _04111_, clk);
  dff _57247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _04090_, clk);
  dff _57248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _04662_, clk);
  dff _57249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _04649_, clk);
  dff _57250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _04635_, clk);
  dff _57251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _04777_, clk);
  dff _57252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _04765_, clk);
  dff _57253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _04739_, clk);
  dff _57254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _07018_, clk);
  dff _57255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _04482_, clk);
  dff _57256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _27010_, clk);
  dff _57257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _04450_, clk);
  dff _57258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _04566_, clk);
  dff _57259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _27011_, clk);
  dff _57260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _04539_, clk);
  dff _57261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _07022_, clk);
  dff _57262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _06546_, clk);
  dff _57263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _04246_, clk);
  dff _57264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _05094_, clk);
  dff _57265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _06370_, clk);
  dff _57266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _04815_, clk);
  dff _57267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _04808_, clk);
  dff _57268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _04884_, clk);
  dff _57269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _04904_, clk);
  dff _57270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _04893_, clk);
  dff _57271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _06364_, clk);
  dff _57272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _27007_, clk);
  dff _57273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _06999_, clk);
  dff _57274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _06549_, clk);
  dff _57275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _05040_, clk);
  dff _57276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _05021_, clk);
  dff _57277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _05002_, clk);
  dff _57278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _05092_, clk);
  dff _57279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _05124_, clk);
  dff _57280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _06994_, clk);
  dff _57281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _05421_, clk);
  dff _57282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _05406_, clk);
  dff _57283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _27004_, clk);
  dff _57284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _27005_, clk);
  dff _57285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _05220_, clk);
  dff _57286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _27006_, clk);
  dff _57287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _05312_, clk);
  dff _57288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _06391_, clk);
  dff _57289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _05991_, clk);
  dff _57290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _05971_, clk);
  dff _57291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _05589_, clk);
  dff _57292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _26998_, clk);
  dff _57293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _06041_, clk);
  dff _57294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _06031_, clk);
  dff _57295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _06974_, clk);
  dff _57296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _05476_, clk);
  dff _57297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _05473_, clk);
  dff _57298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _26999_, clk);
  dff _57299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _27000_, clk);
  dff _57300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _27001_, clk);
  dff _57301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _27002_, clk);
  dff _57302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _06631_, clk);
  dff _57303_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _27003_, clk);
  dff _57304_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _06264_, clk);
  dff _57305_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _06969_, clk);
  dff _57306_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _26997_, clk);
  dff _57307_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _06395_, clk);
  dff _57308_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _06109_, clk);
  dff _57309_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _06098_, clk);
  dff _57310_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _06972_, clk);
  dff _57311_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _06176_, clk);
  dff _57312_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _06403_, clk);
  dff _57313_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _06401_, clk);
  dff _57314_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _06386_, clk);
  dff _57315_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _06492_, clk);
  dff _57316_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _06473_, clk);
  dff _57317_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _06398_, clk);
  dff _57318_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _06633_, clk);
  dff _57319_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _06271_, clk);
  dff _57320_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _06938_, clk);
  dff _57321_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _06571_, clk);
  dff _57322_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _06556_, clk);
  dff _57323_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _06565_, clk);
  dff _57324_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _06560_, clk);
  dff _57325_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _06965_, clk);
  dff _57326_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _06617_, clk);
  dff _57327_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _06640_, clk);
  dff _57328_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _07061_, clk);
  dff _57329_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _26994_, clk);
  dff _57330_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _26995_, clk);
  dff _57331_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _06635_, clk);
  dff _57332_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _06869_, clk);
  dff _57333_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _06859_, clk);
  dff _57334_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _06837_, clk);
  dff _57335_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _06932_, clk);
  dff _57336_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _06917_, clk);
  dff _57337_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _06911_, clk);
  dff _57338_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _06415_, clk);
  dff _57339_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _06707_, clk);
  dff _57340_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _06695_, clk);
  dff _57341_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _26996_, clk);
  dff _57342_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _06758_, clk);
  dff _57343_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _06765_, clk);
  dff _57344_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _07195_, clk);
  dff _57345_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _26993_, clk);
  dff _57346_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _07173_, clk);
  dff _57347_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _07150_, clk);
  dff _57348_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _06430_, clk);
  dff _57349_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _07013_, clk);
  dff _57350_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _06929_, clk);
  dff _57351_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _07081_, clk);
  dff _57352_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _06923_, clk);
  dff _57353_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _07287_, clk);
  dff _57354_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _07310_, clk);
  dff _57355_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _07305_, clk);
  dff _57356_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _26991_, clk);
  dff _57357_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _07098_, clk);
  dff _57358_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _07110_, clk);
  dff _57359_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _07106_, clk);
  dff _57360_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _07396_, clk);
  dff _57361_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _07390_, clk);
  dff _57362_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _07363_, clk);
  dff _57363_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _26989_, clk);
  dff _57364_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _26990_, clk);
  dff _57365_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _07428_, clk);
  dff _57366_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _06440_, clk);
  dff _57367_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _07246_, clk);
  dff _57368_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _07739_, clk);
  dff _57369_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _07851_, clk);
  dff _57370_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _07823_, clk);
  dff _57371_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _06450_, clk);
  dff _57372_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _07640_, clk);
  dff _57373_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _07638_, clk);
  dff _57374_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _07617_, clk);
  dff _57375_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _06901_, clk);
  dff _57376_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _07694_, clk);
  dff _57377_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _26987_, clk);
  dff _57378_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _07495_, clk);
  dff _57379_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _07491_, clk);
  dff _57380_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _07485_, clk);
  dff _57381_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _26988_, clk);
  dff _57382_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _07561_, clk);
  dff _57383_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _07538_, clk);
  dff _57384_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _06457_, clk);
  dff _57385_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _06638_, clk);
  dff _57386_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _08100_, clk);
  dff _57387_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _06887_, clk);
  dff _57388_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _08424_, clk);
  dff _57389_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _08421_, clk);
  dff _57390_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _06885_, clk);
  dff _57391_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _07765_, clk);
  dff _57392_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _26985_, clk);
  dff _57393_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _09228_, clk);
  dff _57394_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _09194_, clk);
  dff _57395_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _06461_, clk);
  dff _57396_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _08454_, clk);
  dff _57397_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _08449_, clk);
  dff _57398_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _08988_, clk);
  dff _57399_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _26986_, clk);
  dff _57400_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _06684_, clk);
  dff _57401_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _25285_, clk);
  dff _57402_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _06679_, clk);
  dff _57403_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _11884_, clk);
  dff _57404_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _12672_, clk);
  dff _57405_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _06689_, clk);
  dff _57406_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _26979_, clk);
  dff _57407_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _06702_, clk);
  dff _57408_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _06824_, clk);
  dff _57409_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _26976_, clk);
  dff _57410_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _10370_, clk);
  dff _57411_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _06833_, clk);
  dff _57412_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _10599_, clk);
  dff _57413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _26977_, clk);
  dff _57414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _06468_, clk);
  dff _57415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _06645_, clk);
  dff _57416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _11195_, clk);
  dff _57417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _26972_, clk);
  dff _57418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _26973_, clk);
  dff _57419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _06591_, clk);
  dff _57420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _10701_, clk);
  dff _57421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _26974_, clk);
  dff _57422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _06831_, clk);
  dff _57423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _26975_, clk);
  dff _57424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _06782_, clk);
  dff _57425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _06595_, clk);
  dff _57426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _11723_, clk);
  dff _57427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _26969_, clk);
  dff _57428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _11855_, clk);
  dff _57429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _06793_, clk);
  dff _57430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _26970_, clk);
  dff _57431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _11499_, clk);
  dff _57432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _11645_, clk);
  dff _57433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _06802_, clk);
  dff _57434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _06648_, clk);
  dff _57435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _11286_, clk);
  dff _57436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _06812_, clk);
  dff _57437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _11414_, clk);
  dff _57438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _06484_, clk);
  dff _57439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _26971_, clk);
  dff _57440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _12617_, clk);
  dff _57441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _06512_, clk);
  dff _57442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _26967_, clk);
  dff _57443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _12260_, clk);
  dff _57444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _12280_, clk);
  dff _57445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _26968_, clk);
  dff _57446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _11962_, clk);
  dff _57447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _06790_, clk);
  dff _57448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _12681_, clk);
  dff _57449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _12679_, clk);
  dff _57450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _06770_, clk);
  dff _57451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _26966_, clk);
  dff _57452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _12711_, clk);
  dff _57453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _06516_, clk);
  dff _57454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _12569_, clk);
  dff _57455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _12565_, clk);
  dff _57456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _06721_, clk);
  dff _57457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _26963_, clk);
  dff _57458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _26964_, clk);
  dff _57459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _11335_, clk);
  dff _57460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _06748_, clk);
  dff _57461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _12249_, clk);
  dff _57462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _06523_, clk);
  dff _57463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _01928_, clk);
  dff _57464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _06754_, clk);
  dff _57465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _05700_, clk);
  dff _57466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _06121_, clk);
  dff _57467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _06521_, clk);
  dff _57468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _26965_, clk);
  dff _57469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _11684_, clk);
  dff _57470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _11410_, clk);
  dff _57471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _06519_, clk);
  dff _57472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _11119_, clk);
  dff _57473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _26961_, clk);
  dff _57474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _11141_, clk);
  dff _57475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _07445_, clk);
  dff _57476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _11147_, clk);
  dff _57477_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _07441_, clk);
  dff _57478_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _11149_, clk);
  dff _57479_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _11159_, clk);
  dff _57480_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _07587_, clk);
  dff _57481_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _11062_, clk);
  dff _57482_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _26959_, clk);
  dff _57483_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _11083_, clk);
  dff _57484_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _07453_, clk);
  dff _57485_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _11094_, clk);
  dff _57486_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _26960_, clk);
  dff _57487_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _11109_, clk);
  dff _57488_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _26952_, clk);
  dff _57489_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _07607_, clk);
  dff _57490_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _10958_, clk);
  dff _57491_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _07487_, clk);
  dff _57492_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _10968_, clk);
  dff _57493_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _07604_, clk);
  dff _57494_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _26953_, clk);
  dff _57495_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _26954_, clk);
  dff _57496_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _07602_, clk);
  dff _57497_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _07724_, clk);
  dff _57498_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _26955_, clk);
  dff _57499_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _07481_, clk);
  dff _57500_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _26956_, clk);
  dff _57501_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _07598_, clk);
  dff _57502_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _26957_, clk);
  dff _57503_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _26958_, clk);
  dff _57504_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _10192_, clk);
  dff _57505_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _26950_, clk);
  dff _57506_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _26951_, clk);
  dff _57507_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _10221_, clk);
  dff _57508_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _07498_, clk);
  dff _57509_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _10806_, clk);
  dff _57510_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _07614_, clk);
  dff _57511_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _10902_, clk);
  dff _57512_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _09167_, clk);
  dff _57513_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _07627_, clk);
  dff _57514_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _09291_, clk);
  dff _57515_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _10089_, clk);
  dff _57516_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _26948_, clk);
  dff _57517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _07702_, clk);
  dff _57518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _26949_, clk);
  dff _57519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _10188_, clk);
  dff _57520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _05862_, clk);
  dff _57521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _05899_, clk);
  dff _57522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _06088_, clk);
  dff _57523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _26946_, clk);
  dff _57524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _06093_, clk);
  dff _57525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _07680_, clk);
  dff _57526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _26947_, clk);
  dff _57527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _09112_, clk);
  dff _57528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _26943_, clk);
  dff _57529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _11349_, clk);
  dff _57530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _26944_, clk);
  dff _57531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _06526_, clk);
  dff _57532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _06535_, clk);
  dff _57533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _07540_, clk);
  dff _57534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _06537_, clk);
  dff _57535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _07654_, clk);
  dff _57536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _11289_, clk);
  dff _57537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _24175_, clk);
  dff _57538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _11296_, clk);
  dff _57539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _22746_, clk);
  dff _57540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _26939_, clk);
  dff _57541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _26940_, clk);
  dff _57542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _11346_, clk);
  dff _57543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _26941_, clk);
  dff _57544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _11315_, clk);
  dff _57545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _11329_, clk);
  dff _57546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _11317_, clk);
  dff _57547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _22866_, clk);
  dff _57548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _11242_, clk);
  dff _57549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _22680_, clk);
  dff _57550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _07579_, clk);
  dff _57551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _26938_, clk);
  dff _57552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _09340_, clk);
  dff _57553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _10844_, clk);
  dff _57554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _09988_, clk);
  dff _57555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _26920_, clk);
  dff _57556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _10880_, clk);
  dff _57557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _09334_, clk);
  dff _57558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _26921_, clk);
  dff _57559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _10886_, clk);
  dff _57560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _10239_, clk);
  dff _57561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _22686_, clk);
  dff _57562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _03822_, clk);
  dff _57563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _06233_, clk);
  dff _57564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _08183_, clk);
  dff _57565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _08451_, clk);
  dff _57566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _09854_, clk);
  dff _57567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _09821_, clk);
  dff _57568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _11406_, clk);
  dff _57569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _11374_, clk);
  dff _57570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _11376_, clk);
  dff _57571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _24383_, clk);
  dff _57572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _11252_, clk);
  dff _57573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _26936_, clk);
  dff _57574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _26937_, clk);
  dff _57575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _11319_, clk);
  dff _57576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _26917_, clk);
  dff _57577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _09347_, clk);
  dff _57578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _10775_, clk);
  dff _57579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _26918_, clk);
  dff _57580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _26919_, clk);
  dff _57581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _10826_, clk);
  dff _57582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _09343_, clk);
  dff _57583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _10114_, clk);
  dff _57584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _10108_, clk);
  dff _57585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _10660_, clk);
  dff _57586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _09354_, clk);
  dff _57587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _10677_, clk);
  dff _57588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _10007_, clk);
  dff _57589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _26916_, clk);
  dff _57590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _10742_, clk);
  dff _57591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _09350_, clk);
  dff _57592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _05084_, clk);
  dff _57593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _22712_, clk);
  dff _57594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _11797_, clk);
  dff _57595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _04499_, clk);
  dff _57596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _03400_, clk);
  dff _57597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _04033_, clk);
  dff _57598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _22721_, clk);
  dff _57599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _11175_, clk);
  dff _57600_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0], clk);
  dff _57601_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1], clk);
  dff _57602_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2], clk);
  dff _57603_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3], clk);
  dff _57604_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4], clk);
  dff _57605_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5], clk);
  dff _57606_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6], clk);
  dff _57607_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7], clk);
  dff _57608_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8], clk);
  dff _57609_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9], clk);
  dff _57610_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10], clk);
  dff _57611_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11], clk);
  dff _57612_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12], clk);
  dff _57613_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13], clk);
  dff _57614_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14], clk);
  dff _57615_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15], clk);
  dff _57616_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16], clk);
  dff _57617_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17], clk);
  dff _57618_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18], clk);
  dff _57619_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19], clk);
  dff _57620_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20], clk);
  dff _57621_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21], clk);
  dff _57622_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22], clk);
  dff _57623_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23], clk);
  dff _57624_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24], clk);
  dff _57625_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25], clk);
  dff _57626_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26], clk);
  dff _57627_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27], clk);
  dff _57628_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28], clk);
  dff _57629_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29], clk);
  dff _57630_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30], clk);
  dff _57631_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31], clk);
  dff _57632_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _27303_, clk);
  dff _57633_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _27304_[0], clk);
  dff _57634_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _27304_[1], clk);
  dff _57635_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _27304_[2], clk);
  dff _57636_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _27304_[3], clk);
  dff _57637_ (\oc8051_top_1.oc8051_sfr1.bit_out , _27305_, clk);
  dff _57638_ (\oc8051_top_1.oc8051_sfr1.wait_data , _27306_, clk);
  dff _57639_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _27307_[0], clk);
  dff _57640_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _27307_[1], clk);
  dff _57641_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _27307_[2], clk);
  dff _57642_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _27307_[3], clk);
  dff _57643_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _27307_[4], clk);
  dff _57644_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _27307_[5], clk);
  dff _57645_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _27307_[6], clk);
  dff _57646_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _27307_[7], clk);
  dff _57647_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _10657_, clk);
  dff _57648_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _10641_, clk);
  dff _57649_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _10471_, clk);
  dff _57650_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _10500_, clk);
  dff _57651_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _10550_, clk);
  dff _57652_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _10516_, clk);
  dff _57653_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _10431_, clk);
  dff _57654_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _10353_, clk);
  dff _57655_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _06742_, clk);
  dff _57656_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _06745_, clk);
  dff _57657_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _06744_, clk);
  dff _57658_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _06752_, clk);
  dff _57659_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _06762_, clk);
  dff _57660_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _06760_, clk);
  dff _57661_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _06767_, clk);
  dff _57662_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _05678_, clk);
  dff _57663_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _10133_, clk);
  dff _57664_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _10132_, clk);
  dff _57665_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _10097_, clk);
  dff _57666_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _10085_, clk);
  dff _57667_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _10074_, clk);
  dff _57668_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _09940_, clk);
  dff _57669_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _10169_, clk);
  dff _57670_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _09964_, clk);
  dff _57671_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _09976_, clk);
  dff _57672_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _10125_, clk);
  dff _57673_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _10050_, clk);
  dff _57674_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _10005_, clk);
  dff _57675_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _10130_, clk);
  dff _57676_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _10128_, clk);
  dff _57677_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _10048_, clk);
  dff _57678_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _10143_, clk);
  dff _57679_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _11762_, clk);
  dff _57680_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _22664_, clk);
  dff _57681_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _09728_, clk);
  dff _57682_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _09843_, clk);
  dff _57683_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _09791_, clk);
  dff _57684_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _09772_, clk);
  dff _57685_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _09750_, clk);
  dff _57686_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22663_, clk);
  dff _57687_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _11828_, clk);
  dff _57688_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _09190_, clk);
  dff _57689_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _11565_, clk);
  dff _57690_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _11704_, clk);
  dff _57691_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _09127_, clk);
  dff _57692_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _22666_, clk);
  dff _57693_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _11663_, clk);
  dff _57694_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _09413_, clk);
  dff _57695_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _22665_, clk);
  dff _57696_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _11656_, clk);
  dff _57697_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _08672_, clk);
  dff _57698_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _08926_, clk);
  dff _57699_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _11683_, clk);
  dff _57700_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _11577_, clk);
  dff _57701_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _11677_, clk);
  dff _57702_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _11637_, clk);
  dff _57703_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _08258_, clk);
  dff _57704_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _08240_, clk);
  dff _57705_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _08221_, clk);
  dff _57706_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _11651_, clk);
  dff _57707_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _07683_, clk);
  dff _57708_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _07512_, clk);
  dff _57709_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _07661_, clk);
  dff _57710_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _07595_, clk);
  dff _57711_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _07548_, clk);
  dff _57712_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _22667_, clk);
  dff _57713_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _07995_, clk);
  dff _57714_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _11710_, clk);
  dff _57715_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _06934_, clk);
  dff _57716_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _06909_, clk);
  dff _57717_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _06893_, clk);
  dff _57718_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _06844_, clk);
  dff _57719_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _22668_, clk);
  dff _57720_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _07281_, clk);
  dff _57721_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _07234_, clk);
  dff _57722_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _11687_, clk);
  dff _57723_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _12192_, clk);
  dff _57724_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _12170_, clk);
  dff _57725_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _12139_, clk);
  dff _57726_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _06267_, clk);
  dff _57727_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _12529_, clk);
  dff _57728_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _12395_, clk);
  dff _57729_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _12507_, clk);
  dff _57730_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _11111_, clk);
  dff _57731_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _11583_, clk);
  dff _57732_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _11558_, clk);
  dff _57733_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _11482_, clk);
  dff _57734_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _11413_, clk);
  dff _57735_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _06280_, clk);
  dff _57736_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _11954_, clk);
  dff _57737_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _11878_, clk);
  dff _57738_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _11086_, clk);
  dff _57739_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _10891_, clk);
  dff _57740_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _10718_, clk);
  dff _57741_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _10855_, clk);
  dff _57742_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _10829_, clk);
  dff _57743_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _10779_, clk);
  dff _57744_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _10757_, clk);
  dff _57745_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _06293_, clk);
  dff _57746_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _10940_, clk);
  dff _57747_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _10236_, clk);
  dff _57748_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _10212_, clk);
  dff _57749_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _10186_, clk);
  dff _57750_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _10161_, clk);
  dff _57751_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _06326_, clk);
  dff _57752_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _10540_, clk);
  dff _57753_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _10409_, clk);
  dff _57754_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _11053_, clk);
  dff _57755_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _10364_, clk);
  dff _57756_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _10338_, clk);
  dff _57757_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _10329_, clk);
  dff _57758_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _10317_, clk);
  dff _57759_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _10330_, clk);
  dff _57760_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _10341_, clk);
  dff _57761_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _10039_, clk);
  dff _57762_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _06939_, clk);
  dff _57763_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _07222_, clk);
  dff _57764_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _07218_, clk);
  dff _57765_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _07231_, clk);
  dff _57766_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _07226_, clk);
  dff _57767_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _07228_, clk);
  dff _57768_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _07241_, clk);
  dff _57769_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _07237_, clk);
  dff _57770_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _06960_, clk);
  dff _57771_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _22634_, clk);
  dff _57772_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _01412_, clk);
  dff _57773_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _04590_, clk);
  dff _57774_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _11690_, clk);
  dff _57775_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _11512_, clk);
  dff _57776_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _04585_, clk);
  dff _57777_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _00832_, clk);
  dff _57778_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _05875_, clk);
  dff _57779_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _03997_, clk);
  dff _57780_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _06794_, clk);
  dff _57781_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _04624_, clk);
  dff _57782_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _00740_, clk);
  dff _57783_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _09365_, clk);
  dff _57784_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _15153_, clk);
  dff _57785_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _12540_, clk);
  dff _57786_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _18600_, clk);
  dff _57787_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _26774_, clk);
  dff _57788_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _02663_, clk);
  dff _57789_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _22657_, clk);
  dff _57790_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _10382_, clk);
  dff _57791_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _05196_, clk);
  dff _57792_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _03628_, clk);
  dff _57793_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _02555_, clk);
  dff _57794_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _04642_, clk);
  dff _57795_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _10788_, clk);
  dff _57796_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _11085_, clk);
  dff _57797_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _10873_, clk);
  dff _57798_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _22630_, clk);
  dff _57799_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _12736_, clk);
  dff _57800_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _12731_, clk);
  dff _57801_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _04657_, clk);
  dff _57802_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _23032_, clk);
  dff _57803_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _26617_, clk);
  dff _57804_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _26690_, clk);
  dff _57805_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _09769_, clk);
  dff _57806_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _23573_, clk);
  dff _57807_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _04338_, clk);
  dff _57808_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _12720_, clk);
  dff _57809_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _12717_, clk);
  dff _57810_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _04659_, clk);
  dff _57811_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _26382_, clk);
  dff _57812_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _08395_, clk);
  dff _57813_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _15132_, clk);
  dff _57814_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _17294_, clk);
  dff _57815_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _06866_, clk);
  dff _57816_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _22655_, clk);
  dff _57817_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _22654_, clk);
  dff _57818_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _04546_, clk);
  dff _57819_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _22653_, clk);
  dff _57820_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _07802_, clk);
  dff _57821_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _03406_, clk);
  dff _57822_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _07838_, clk);
  dff _57823_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _07834_, clk);
  dff _57824_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _07832_, clk);
  dff _57825_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _07830_, clk);
  dff _57826_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _07828_, clk);
  dff _57827_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _11891_, clk);
  dff _57828_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _07779_, clk);
  dff _57829_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _07773_, clk);
  dff _57830_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _07769_, clk);
  dff _57831_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _07767_, clk);
  dff _57832_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _03409_, clk);
  dff _57833_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _10384_, clk);
  dff _57834_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _07716_, clk);
  dff _57835_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _22652_, clk);
  dff _57836_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _22648_, clk);
  dff _57837_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _03444_, clk);
  dff _57838_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _07656_, clk);
  dff _57839_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _07651_, clk);
  dff _57840_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _07646_, clk);
  dff _57841_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _03477_, clk);
  dff _57842_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _07699_, clk);
  dff _57843_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _07697_, clk);
  dff _57844_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _22647_, clk);
  dff _57845_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _07596_, clk);
  dff _57846_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _07593_, clk);
  dff _57847_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _03486_, clk);
  dff _57848_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _07630_, clk);
  dff _57849_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _07609_, clk);
  dff _57850_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _07622_, clk);
  dff _57851_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _07620_, clk);
  dff _57852_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _22645_, clk);
  dff _57853_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _22644_, clk);
  dff _57854_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _07549_, clk);
  dff _57855_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _07546_, clk);
  dff _57856_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _03500_, clk);
  dff _57857_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _07575_, clk);
  dff _57858_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _07565_, clk);
  dff _57859_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _07573_, clk);
  dff _57860_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _07571_, clk);
  dff _57861_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01438_, clk);
  dff _57862_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _23001_, clk);
  dff _57863_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _23013_, clk);
  dff _57864_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _23010_, clk);
  dff _57865_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _23007_, clk);
  dff _57866_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _22760_, clk);
  dff _57867_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _22873_, clk);
  dff _57868_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _22752_, clk);
  dff _57869_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _22753_, clk);
  dff _57870_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _22755_, clk);
  dff _57871_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _22776_, clk);
  dff _57872_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22790_, clk);
  dff _57873_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01419_, clk);
  dff _57874_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _01386_, clk);
  dff _57875_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _25815_, clk);
  dff _57876_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _25814_, clk);
  dff _57877_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _01455_, clk);
  dff _57878_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _25874_, clk);
  dff _57879_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _25872_, clk);
  dff _57880_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _22851_, clk);
  dff _57881_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _01452_, clk);
  dff _57882_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _22779_, clk);
  dff _57883_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _22792_, clk);
  dff _57884_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _22911_, clk);
  dff _57885_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _01384_, clk);
  dff _57886_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _22650_, clk);
  dff _57887_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _22651_, clk);
  dff _57888_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _22955_, clk);
  dff _57889_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _22649_, clk);
  dff _57890_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _22988_, clk);
  dff _57891_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _22933_, clk);
  dff _57892_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _22965_, clk);
  dff _57893_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _01407_, clk);
  dff _57894_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _25786_, clk);
  dff _57895_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _25778_, clk);
  dff _57896_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _25781_, clk);
  dff _57897_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _01466_, clk);
  dff _57898_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _22831_, clk);
  dff _57899_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _22856_, clk);
  dff _57900_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _22858_, clk);
  dff _57901_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _25800_, clk);
  dff _57902_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _22751_, clk);
  dff _57903_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _22750_, clk);
  dff _57904_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _22749_, clk);
  dff _57905_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _22748_, clk);
  dff _57906_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _22747_, clk);
  dff _57907_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _22745_, clk);
  dff _57908_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _22744_, clk);
  dff _57909_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _22743_, clk);
  dff _57910_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _22742_, clk);
  dff _57911_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _22741_, clk);
  dff _57912_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _25796_, clk);
  dff _57913_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _22739_, clk);
  dff _57914_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _22738_, clk);
  dff _57915_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _22646_, clk);
  dff _57916_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _22737_, clk);
  dff _57917_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _04622_, clk);
  dff _57918_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _22736_, clk);
  dff _57919_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _22735_, clk);
  dff _57920_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _01457_, clk);
  dff _57921_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _22734_, clk);
  dff _57922_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _22733_, clk);
  dff _57923_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _22732_, clk);
  dff _57924_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _22731_, clk);
  dff _57925_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _22730_, clk);
  dff _57926_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _22729_, clk);
  dff _57927_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _22728_, clk);
  dff _57928_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _01382_, clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
endmodule
