
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_inc_dir_iram, property_invalid_inc_acc, property_invalid_pcp1, property_invalid_pcp2, property_invalid_pcp3, property_invalid_sjmp, property_invalid_ljmp, property_invalid_ajmp, property_invalid_jc, property_invalid_jnc);
  wire [7:0] _00000_;
  wire _00001_;
  wire _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire [15:0] _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire [7:0] _36857_;
  wire _36858_;
  wire [1:0] _36859_;
  wire [5:0] _36860_;
  wire [7:0] _36861_;
  wire [1:0] _36862_;
  wire [15:0] _36863_;
  wire [7:0] _36864_;
  wire [7:0] _36865_;
  wire [7:0] _36866_;
  wire [2:0] _36867_;
  wire [2:0] _36868_;
  wire [1:0] _36869_;
  wire [7:0] _36870_;
  wire _36871_;
  wire [1:0] _36872_;
  wire [1:0] _36873_;
  wire [2:0] _36874_;
  wire [2:0] _36875_;
  wire [1:0] _36876_;
  wire [3:0] _36877_;
  wire [1:0] _36878_;
  wire _36879_;
  wire _36880_;
  wire [7:0] _36881_;
  wire [7:0] _36882_;
  wire [7:0] _36883_;
  wire [7:0] _36884_;
  wire [7:0] _36885_;
  wire [7:0] _36886_;
  wire [7:0] _36887_;
  wire [7:0] _36888_;
  wire [15:0] _36889_;
  wire [15:0] _36890_;
  wire _36891_;
  wire [4:0] _36892_;
  wire [7:0] _36893_;
  wire [7:0] _36894_;
  wire [7:0] _36895_;
  wire _36896_;
  wire _36897_;
  wire [7:0] _36898_;
  wire [15:0] _36899_;
  wire [15:0] _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire [7:0] _36904_;
  wire [2:0] _36905_;
  wire [7:0] _36906_;
  wire [7:0] _36907_;
  wire _36908_;
  wire [7:0] _36909_;
  wire _36910_;
  wire _36911_;
  wire [3:0] _36912_;
  wire [31:0] _36913_;
  wire [31:0] _36914_;
  wire [7:0] _36915_;
  wire _36916_;
  wire _36917_;
  wire [15:0] _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire [15:0] _36922_;
  wire _36923_;
  wire _36924_;
  wire [7:0] _36925_;
  wire _36926_;
  wire [2:0] _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire [7:0] _38984_;
  wire _38985_;
  wire [3:0] _38986_;
  wire _38987_;
  wire _38988_;
  wire [7:0] _38989_;
  wire _38990_;
  wire [7:0] _38991_;
  wire [7:0] _38992_;
  wire [7:0] _38993_;
  wire [7:0] _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire [7:0] _38998_;
  wire [1:0] _38999_;
  wire _39000_;
  wire [2:0] _39001_;
  wire [2:0] _39002_;
  wire [1:0] _39003_;
  wire [1:0] _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire [3:0] _39009_;
  wire [7:0] _39010_;
  wire [7:0] _39011_;
  wire [7:0] _39012_;
  wire [7:0] _39013_;
  wire [7:0] _39014_;
  wire [7:0] _39015_;
  wire [6:0] _39016_;
  wire _39017_;
  wire [7:0] _39018_;
  wire _39019_;
  wire _39020_;
  wire [7:0] _39021_;
  wire [7:0] _39022_;
  wire _39023_;
  wire _39024_;
  wire [7:0] _39025_;
  wire [7:0] _39026_;
  wire _39027_;
  wire [7:0] _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire [7:0] _39033_;
  wire [7:0] _39034_;
  wire _39035_;
  wire [7:0] _39036_;
  wire [7:0] _39037_;
  wire _39038_;
  wire [7:0] _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire [1:0] _39046_;
  wire [3:0] _39047_;
  wire [7:0] _39048_;
  wire [11:0] _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire [3:0] _39055_;
  wire [10:0] _39056_;
  wire [7:0] _39057_;
  wire [7:0] _39058_;
  wire [7:0] acc;
  wire [7:0] acc_reg;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire cy_reg;
  wire first_instr;
  wire [7:0] iram_op1;
  wire [7:0] iram_op1_reg;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire [7:0] op1_out_r;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  wire pc_change_r;
  wire pc_inc_acc_r;
  wire pc_inc_dir_r;
  output property_invalid_ajmp;
  output property_invalid_inc_acc;
  output property_invalid_inc_dir_iram;
  output property_invalid_jc;
  output property_invalid_jnc;
  output property_invalid_ljmp;
  output property_invalid_pcp1;
  output property_invalid_pcp2;
  output property_invalid_pcp3;
  output property_invalid_sjmp;
  wire [7:0] psw;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [31:0] word_in;
  and _39059_ (_33127_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _39060_ (_33128_, _33127_);
  not _39061_ (_33129_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _39062_ (_33130_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or _39063_ (_33131_, _33130_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _39064_ (_33132_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _39065_ (_33133_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _39066_ (_33134_, _33133_, _33132_);
  and _39067_ (_33135_, _33130_, _33129_);
  and _39068_ (_33136_, _33135_, _33134_);
  and _39069_ (_33137_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _39070_ (_33138_, _33137_);
  not _39071_ (_33139_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _39072_ (_33140_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _39073_ (_33141_, _33140_);
  not _39074_ (_33142_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  not _39075_ (_33143_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not _39076_ (_33144_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _39077_ (_33145_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _33144_);
  nand _39078_ (_33146_, _33145_, _33143_);
  or _39079_ (_33147_, _33146_, _33142_);
  not _39080_ (_33148_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _39081_ (_33149_, _33148_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _39082_ (_33150_, _33149_, _33143_);
  nand _39083_ (_33151_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _39084_ (_33152_, _33151_, _33147_);
  nor _39085_ (_33153_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _39086_ (_33154_, _33153_, _33143_);
  nand _39087_ (_33155_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _39088_ (_33156_, _33153_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _39089_ (_33157_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _39090_ (_33158_, _33157_, _33155_);
  and _39091_ (_33159_, _33153_, _33143_);
  nand _39092_ (_33160_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _39093_ (_33161_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _39094_ (_33162_, _33161_, _33143_);
  nand _39095_ (_33163_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and _39096_ (_33164_, _33163_, _33160_);
  and _39097_ (_33165_, _33164_, _33158_);
  nand _39098_ (_33166_, _33165_, _33152_);
  nand _39099_ (_33167_, _33166_, _33141_);
  nand _39100_ (_33168_, _33167_, _33139_);
  nor _39101_ (_33169_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _33139_);
  nor _39102_ (_33170_, _33169_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand _39103_ (_33171_, _33170_, _33168_);
  and _39104_ (_33172_, _33171_, _33138_);
  nand _39105_ (_33173_, _33172_, _33136_);
  not _39106_ (_33174_, _33134_);
  nor _39107_ (_33175_, _33135_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _39108_ (_33176_, _33175_, _33174_);
  and _39109_ (_33177_, _33176_, _33173_);
  and _39110_ (_33178_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _39111_ (_33179_, _33178_);
  nand _39112_ (_33180_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand _39113_ (_33181_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _39114_ (_33182_, _33181_, _33180_);
  nand _39115_ (_33183_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  not _39116_ (_33184_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _39117_ (_33185_, _33146_, _33184_);
  and _39118_ (_33186_, _33185_, _33183_);
  nand _39119_ (_33187_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand _39120_ (_33188_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _39121_ (_33189_, _33188_, _33187_);
  and _39122_ (_33190_, _33189_, _33186_);
  and _39123_ (_33191_, _33190_, _33182_);
  or _39124_ (_33192_, _33191_, _33140_);
  nand _39125_ (_33193_, _33192_, _33139_);
  nor _39126_ (_33194_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _33139_);
  nor _39127_ (_33195_, _33194_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand _39128_ (_33196_, _33195_, _33193_);
  and _39129_ (_33197_, _33196_, _33179_);
  nand _39130_ (_33198_, _33197_, _33136_);
  nor _39131_ (_33199_, _33135_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _39132_ (_33200_, _33199_, _33174_);
  and _39133_ (_33201_, _33200_, _33198_);
  nor _39134_ (_33202_, _33201_, _33177_);
  and _39135_ (_33203_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _39136_ (_33204_, _33203_);
  nand _39137_ (_33205_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not _39138_ (_33206_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _39139_ (_33207_, _33146_, _33206_);
  and _39140_ (_33208_, _33207_, _33205_);
  nand _39141_ (_33209_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand _39142_ (_33210_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _39143_ (_33211_, _33210_, _33209_);
  nand _39144_ (_33212_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nand _39145_ (_33213_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _39146_ (_33214_, _33213_, _33212_);
  and _39147_ (_33215_, _33214_, _33211_);
  nand _39148_ (_33216_, _33215_, _33208_);
  nand _39149_ (_33217_, _33216_, _33141_);
  nand _39150_ (_33218_, _33217_, _33139_);
  nor _39151_ (_33219_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _33139_);
  nor _39152_ (_33220_, _33219_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand _39153_ (_33221_, _33220_, _33218_);
  and _39154_ (_33222_, _33221_, _33204_);
  nand _39155_ (_33223_, _33222_, _33136_);
  nor _39156_ (_33224_, _33135_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _39157_ (_33225_, _33224_, _33174_);
  and _39158_ (_33226_, _33225_, _33223_);
  not _39159_ (_33227_, _33136_);
  and _39160_ (_33228_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _39161_ (_33229_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _39162_ (_33230_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _39163_ (_33231_, _33230_, _33229_);
  or _39164_ (_33232_, _33231_, _33228_);
  and _39165_ (_33233_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or _39166_ (_33234_, _33233_, _33140_);
  and _39167_ (_33235_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  not _39168_ (_33236_, _33146_);
  and _39169_ (_33237_, _33236_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _39170_ (_33238_, _33237_, _33235_);
  or _39171_ (_33239_, _33238_, _33234_);
  or _39172_ (_33240_, _33239_, _33232_);
  or _39173_ (_33241_, _33240_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _39174_ (_33242_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _33139_);
  nor _39175_ (_33243_, _33242_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _39176_ (_33244_, _33243_, _33241_);
  and _39177_ (_33245_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or _39178_ (_33246_, _33245_, _33244_);
  or _39179_ (_33247_, _33246_, _33227_);
  nor _39180_ (_33248_, _33135_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _39181_ (_33249_, _33248_, _33174_);
  and _39182_ (_33250_, _33249_, _33247_);
  nor _39183_ (_33251_, _33250_, _33226_);
  and _39184_ (_33252_, _33251_, _33202_);
  nand _39185_ (_33253_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nand _39186_ (_33254_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _39187_ (_33255_, _33254_, _33253_);
  not _39188_ (_33256_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _39189_ (_33257_, _33146_, _33256_);
  and _39190_ (_33258_, _33141_, _33257_);
  and _39191_ (_33259_, _33258_, _33255_);
  nand _39192_ (_33260_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nand _39193_ (_33261_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nand _39194_ (_33262_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _39195_ (_33263_, _33262_, _33261_);
  and _39196_ (_33264_, _33263_, _33260_);
  nand _39197_ (_33265_, _33264_, _33259_);
  or _39198_ (_33266_, _33265_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _39199_ (_33267_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _33139_);
  nor _39200_ (_33268_, _33267_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _39201_ (_33269_, _33268_, _33266_);
  and _39202_ (_33270_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or _39203_ (_33271_, _33270_, _33269_);
  or _39204_ (_33272_, _33271_, _33227_);
  nor _39205_ (_33273_, _33135_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _39206_ (_33274_, _33273_, _33174_);
  and _39207_ (_33275_, _33274_, _33272_);
  and _39208_ (_33276_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _39209_ (_33277_, _33276_);
  nand _39210_ (_33278_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nand _39211_ (_33279_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _39212_ (_33280_, _33279_, _33278_);
  nand _39213_ (_33281_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand _39214_ (_33282_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _39215_ (_33283_, _33282_, _33281_);
  nand _39216_ (_33284_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not _39217_ (_33285_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or _39218_ (_33286_, _33146_, _33285_);
  and _39219_ (_33287_, _33286_, _33284_);
  and _39220_ (_33288_, _33287_, _33283_);
  nand _39221_ (_33289_, _33288_, _33280_);
  and _39222_ (_33290_, _33289_, _33141_);
  or _39223_ (_33291_, _33290_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _39224_ (_33292_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _33139_);
  nor _39225_ (_33293_, _33292_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand _39226_ (_33294_, _33293_, _33291_);
  and _39227_ (_33295_, _33294_, _33277_);
  nand _39228_ (_33296_, _33295_, _33136_);
  nor _39229_ (_33297_, _33135_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _39230_ (_33298_, _33297_, _33174_);
  and _39231_ (_33299_, _33298_, _33296_);
  and _39232_ (_33300_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  not _39233_ (_33301_, _33300_);
  nand _39234_ (_33302_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not _39235_ (_33303_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _39236_ (_33304_, _33146_, _33303_);
  and _39237_ (_33305_, _33304_, _33302_);
  nand _39238_ (_33306_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand _39239_ (_33307_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _39240_ (_33308_, _33307_, _33306_);
  nand _39241_ (_33309_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand _39242_ (_33310_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and _39243_ (_33311_, _33310_, _33309_);
  and _39244_ (_33312_, _33311_, _33308_);
  and _39245_ (_33313_, _33312_, _33305_);
  or _39246_ (_33314_, _33313_, _33140_);
  nand _39247_ (_33315_, _33314_, _33139_);
  nor _39248_ (_33316_, _33139_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  nor _39249_ (_33317_, _33316_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand _39250_ (_33318_, _33317_, _33315_);
  and _39251_ (_33319_, _33318_, _33301_);
  nand _39252_ (_33320_, _33319_, _33136_);
  nor _39253_ (_33321_, _33135_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _39254_ (_33322_, _33321_, _33174_);
  and _39255_ (_33323_, _33322_, _33320_);
  not _39256_ (_33324_, _33323_);
  and _39257_ (_33325_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _39258_ (_33326_, _33325_);
  nand _39259_ (_33327_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand _39260_ (_33328_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _39261_ (_33329_, _33328_, _33327_);
  nand _39262_ (_33330_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  not _39263_ (_33331_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _39264_ (_33332_, _33146_, _33331_);
  and _39265_ (_33333_, _33332_, _33330_);
  nand _39266_ (_33334_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand _39267_ (_33335_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _39268_ (_33336_, _33335_, _33334_);
  and _39269_ (_33337_, _33336_, _33333_);
  and _39270_ (_33338_, _33337_, _33329_);
  or _39271_ (_33339_, _33338_, _33140_);
  nand _39272_ (_33340_, _33339_, _33139_);
  nor _39273_ (_33341_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _33139_);
  nor _39274_ (_33342_, _33341_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand _39275_ (_33343_, _33342_, _33340_);
  nand _39276_ (_33344_, _33343_, _33326_);
  or _39277_ (_33345_, _33344_, _33227_);
  nor _39278_ (_33346_, _33135_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _39279_ (_33347_, _33346_, _33174_);
  nand _39280_ (_33348_, _33347_, _33345_);
  and _39281_ (_33349_, _33348_, _33324_);
  and _39282_ (_33350_, _33349_, _33299_);
  and _39283_ (_33351_, _33350_, _33275_);
  and _39284_ (_33352_, _33351_, _33252_);
  not _39285_ (_33353_, _33352_);
  not _39286_ (_33354_, _33275_);
  and _39287_ (_33355_, _33350_, _33354_);
  nand _39288_ (_33356_, _33355_, _33252_);
  not _39289_ (_33357_, _33299_);
  and _39290_ (_33358_, _33349_, _33357_);
  and _39291_ (_33359_, _33358_, _33275_);
  nand _39292_ (_33360_, _33359_, _33252_);
  and _39293_ (_33361_, _33360_, _33356_);
  and _39294_ (_33362_, _33361_, _33353_);
  not _39295_ (_33363_, _33362_);
  not _39296_ (_33364_, _33201_);
  and _39297_ (_33365_, _33364_, _33177_);
  not _39298_ (_33366_, _33250_);
  and _39299_ (_33367_, _33366_, _33226_);
  and _39300_ (_33368_, _33367_, _33365_);
  not _39301_ (_33369_, _33348_);
  and _39302_ (_33370_, _33299_, _33369_);
  and _39303_ (_33371_, _33370_, _33323_);
  and _39304_ (_33372_, _33371_, _33354_);
  and _39305_ (_33373_, _33372_, _33368_);
  and _39306_ (_33374_, _33348_, _33323_);
  and _39307_ (_33375_, _33374_, _33299_);
  and _39308_ (_33376_, _33375_, _33275_);
  and _39309_ (_33377_, _33368_, _33376_);
  or _39310_ (_33378_, _33377_, _33373_);
  or _39311_ (_33379_, _33378_, _33363_);
  nor _39312_ (_33380_, _33299_, _33348_);
  and _39313_ (_33381_, _33380_, _33324_);
  and _39314_ (_33382_, _33381_, _33275_);
  or _39315_ (_33383_, _33350_, _33382_);
  and _39316_ (_33384_, _33383_, _33368_);
  and _39317_ (_33385_, _33202_, _33250_);
  and _39318_ (_33386_, _33382_, _33385_);
  and _39319_ (_33387_, _33374_, _33357_);
  and _39320_ (_33388_, _33387_, _33354_);
  nor _39321_ (_33389_, _33177_, _33366_);
  nor _39322_ (_33390_, _33201_, _33226_);
  and _39323_ (_33391_, _33390_, _33389_);
  and _39324_ (_33392_, _33391_, _33388_);
  or _39325_ (_33393_, _33392_, _33386_);
  or _39326_ (_33394_, _33393_, _33384_);
  and _39327_ (_33395_, _33358_, _33354_);
  and _39328_ (_33396_, _33395_, _33368_);
  and _39329_ (_33397_, _33375_, _33354_);
  and _39330_ (_33398_, _33365_, _33250_);
  and _39331_ (_33399_, _33398_, _33397_);
  or _39332_ (_33400_, _33399_, _33396_);
  or _39333_ (_33401_, _33400_, _33394_);
  or _39334_ (_33402_, _33401_, _33379_);
  and _39335_ (_33403_, _33381_, _33354_);
  and _39336_ (_33404_, _33368_, _33403_);
  and _39337_ (_33405_, _33397_, _33252_);
  or _39338_ (_33406_, _33405_, _33404_);
  and _39339_ (_33407_, _33370_, _33324_);
  and _39340_ (_33408_, _33407_, _33275_);
  and _39341_ (_33409_, _33391_, _33408_);
  and _39342_ (_33410_, _33385_, _33226_);
  and _39343_ (_33411_, _33403_, _33410_);
  and _39344_ (_33412_, _33391_, _33403_);
  or _39345_ (_33413_, _33412_, _33411_);
  or _39346_ (_33414_, _33413_, _33409_);
  nor _39347_ (_33415_, _33414_, _33406_);
  and _39348_ (_33416_, _33252_, _33376_);
  and _39349_ (_33417_, _33380_, _33323_);
  and _39350_ (_33418_, _33417_, _33275_);
  and _39351_ (_33419_, _33418_, _33368_);
  and _39352_ (_33420_, _33359_, _33368_);
  nor _39353_ (_33421_, _33420_, _33419_);
  nand _39354_ (_33422_, _33391_, _33376_);
  and _39355_ (_33423_, _33417_, _33354_);
  nand _39356_ (_33424_, _33391_, _33423_);
  and _39357_ (_33425_, _33424_, _33422_);
  nand _39358_ (_33426_, _33425_, _33421_);
  nor _39359_ (_33427_, _33426_, _33416_);
  and _39360_ (_33428_, _33427_, _33415_);
  and _39361_ (_33429_, _33407_, _33354_);
  and _39362_ (_33430_, _33429_, _33385_);
  and _39363_ (_33431_, _33252_, _33417_);
  or _39364_ (_33432_, _33431_, _33430_);
  and _39365_ (_33433_, _33429_, _33368_);
  and _39366_ (_33434_, _33368_, _33423_);
  or _39367_ (_33435_, _33434_, _33433_);
  and _39368_ (_33436_, _33388_, _33368_);
  and _39369_ (_33437_, _33387_, _33275_);
  and _39370_ (_33438_, _33437_, _33391_);
  or _39371_ (_33439_, _33438_, _33436_);
  nor _39372_ (_33440_, _33439_, _33435_);
  nand _39373_ (_33441_, _33437_, _33368_);
  nand _39374_ (_33442_, _33391_, _33350_);
  and _39375_ (_33443_, _33201_, _33354_);
  nand _39376_ (_33444_, _33443_, _33375_);
  and _39377_ (_33445_, _33444_, _33442_);
  and _39378_ (_33446_, _33445_, _33441_);
  nand _39379_ (_33447_, _33391_, _33418_);
  nand _39380_ (_33448_, _33391_, _33397_);
  and _39381_ (_33449_, _33448_, _33447_);
  and _39382_ (_33450_, _33449_, _33446_);
  nand _39383_ (_33451_, _33450_, _33440_);
  nor _39384_ (_33452_, _33451_, _33432_);
  nand _39385_ (_33453_, _33452_, _33428_);
  or _39386_ (_33454_, _33453_, _33402_);
  nand _39387_ (_33455_, _33454_, _33131_);
  not _39388_ (_33456_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _39389_ (_33457_, _33129_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _39390_ (_33458_, _33457_, _33456_);
  and _39391_ (_33459_, _33252_, _33407_);
  and _39392_ (_33460_, _33459_, _33458_);
  and _39393_ (_33461_, _33458_, _33252_);
  and _39394_ (_33462_, _33461_, _33381_);
  nor _39395_ (_33463_, _33462_, _33460_);
  not _39396_ (_33464_, _33226_);
  and _39397_ (_33465_, _33385_, _33464_);
  and _39398_ (_33466_, _33350_, _33465_);
  and _39399_ (_33467_, \oc8051_top_1.oc8051_decoder1.state [0], _33129_);
  and _39400_ (_33468_, _33467_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _39401_ (_33469_, _33468_, _33466_);
  not _39402_ (_33470_, _33469_);
  and _39403_ (_33471_, _33470_, _33463_);
  nand _39404_ (_33472_, _33471_, _33455_);
  nand _39405_ (_33473_, _33472_, _33129_);
  and _39406_ (_33474_, _33473_, _33128_);
  not _39407_ (_33475_, _33474_);
  and _39408_ (_33476_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _39409_ (_33477_, _33131_);
  and _39410_ (_33478_, _33251_, _33365_);
  and _39411_ (_33479_, _33478_, _33388_);
  and _39412_ (_33480_, _33478_, _33397_);
  nor _39413_ (_33481_, _33480_, _33479_);
  and _39414_ (_33482_, _33437_, _33410_);
  not _39415_ (_33483_, _33482_);
  nand _39416_ (_33484_, _33410_, _33408_);
  nand _39417_ (_33485_, _33397_, _33410_);
  and _39418_ (_33486_, _33485_, _33484_);
  and _39419_ (_33487_, _33486_, _33483_);
  and _39420_ (_33488_, _33487_, _33481_);
  nor _39421_ (_33489_, _33488_, _33477_);
  not _39422_ (_33490_, _33130_);
  and _39423_ (_33491_, _33480_, _33129_);
  and _39424_ (_33492_, _33491_, _33490_);
  and _39425_ (_33493_, _33479_, _33477_);
  nor _39426_ (_33494_, _33493_, _33492_);
  and _39427_ (_33495_, _33494_, _33463_);
  not _39428_ (_33496_, _33495_);
  nor _39429_ (_33497_, _33496_, _33489_);
  nor _39430_ (_33498_, _33497_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _39431_ (_33499_, _33498_, _33476_);
  not _39432_ (_33500_, _33499_);
  and _39433_ (_33501_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _39434_ (_33502_, _33501_);
  and _39435_ (_33503_, _33398_, _33383_);
  and _39436_ (_33504_, _33398_, _33376_);
  nand _39437_ (_33505_, _33398_, _33358_);
  not _39438_ (_33506_, _33505_);
  and _39439_ (_33507_, _33398_, _33388_);
  or _39440_ (_33508_, _33507_, _33506_);
  nor _39441_ (_33509_, _33508_, _33504_);
  not _39442_ (_33510_, _33466_);
  nand _39443_ (_33511_, _33398_, _33429_);
  and _39444_ (_33512_, _33511_, _33510_);
  nand _39445_ (_33513_, _33512_, _33509_);
  nor _39446_ (_33514_, _33513_, _33503_);
  and _39447_ (_33515_, _33398_, _33354_);
  nor _39448_ (_33516_, _33371_, _33381_);
  not _39449_ (_33517_, _33516_);
  nand _39450_ (_33518_, _33517_, _33515_);
  nand _39451_ (_33519_, _33418_, _33252_);
  nand _39452_ (_33520_, _33398_, _33417_);
  not _39453_ (_33521_, _33520_);
  and _39454_ (_33522_, _33398_, _33437_);
  nor _39455_ (_33523_, _33522_, _33521_);
  and _39456_ (_33524_, _33523_, _33519_);
  and _39457_ (_33525_, _33524_, _33518_);
  and _39458_ (_33526_, _33525_, _33487_);
  nand _39459_ (_33527_, _33526_, _33514_);
  nand _39460_ (_33528_, _33527_, _33131_);
  nor _39461_ (_33529_, _33469_, _33460_);
  nand _39462_ (_33530_, _33529_, _33528_);
  nand _39463_ (_33531_, _33530_, _33129_);
  and _39464_ (_33532_, _33531_, _33502_);
  nor _39465_ (_33533_, _33532_, _33500_);
  and _39466_ (_33534_, _33533_, _33475_);
  not _39467_ (_33535_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _39468_ (_33536_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _33129_);
  and _39469_ (_33537_, _33536_, _33535_);
  and _39470_ (_33538_, _33537_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _39471_ (_33539_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  not _39472_ (_33540_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _39473_ (_33541_, _33537_, _33540_);
  and _39474_ (_33542_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor _39475_ (_33543_, _33542_, _33539_);
  and _39476_ (_33544_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _33129_);
  nor _39477_ (_33545_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _39478_ (_33546_, _33545_, _33544_);
  and _39479_ (_33547_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not _39480_ (_33548_, _33547_);
  not _39481_ (_33549_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _39482_ (_33550_, _33544_, _33540_);
  and _39483_ (_33551_, _33550_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _39484_ (_33552_, _33551_, _33549_);
  and _39485_ (_33553_, _33545_, _33535_);
  or _39486_ (_33554_, _33553_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _39487_ (_33555_, _33554_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _39488_ (_33556_, _33555_, _33552_);
  and _39489_ (_33557_, _33556_, _33548_);
  and _39490_ (_33558_, _33557_, _33543_);
  not _39491_ (_33559_, _33558_);
  and _39492_ (_33560_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _39493_ (_33561_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _39494_ (_33562_, _33561_, _33560_);
  and _39495_ (_33563_, _33562_, _33551_);
  and _39496_ (_33564_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor _39497_ (_33565_, _33564_, _33563_);
  and _39498_ (_33566_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and _39499_ (_33567_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and _39500_ (_33568_, _33554_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or _39501_ (_33569_, _33568_, _33567_);
  nor _39502_ (_33570_, _33569_, _33566_);
  and _39503_ (_33571_, _33570_, _33565_);
  and _39504_ (_33572_, _33571_, _33559_);
  and _39505_ (_33573_, _33560_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _39506_ (_33574_, _33573_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _39507_ (_33575_, _33574_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _39508_ (_33576_, _33575_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _39509_ (_33577_, _33576_);
  not _39510_ (_33578_, _33551_);
  nor _39511_ (_33579_, _33575_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _39512_ (_33580_, _33579_, _33578_);
  and _39513_ (_33581_, _33580_, _33577_);
  not _39514_ (_33582_, _33581_);
  and _39515_ (_33583_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _39516_ (_33584_, _33583_, _33544_);
  and _39517_ (_33585_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor _39518_ (_33586_, _33585_, _33584_);
  and _39519_ (_33587_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _39520_ (_33588_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor _39521_ (_33589_, _33588_, _33587_);
  and _39522_ (_33590_, _33589_, _33586_);
  and _39523_ (_33591_, _33590_, _33582_);
  and _39524_ (_33592_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor _39525_ (_33593_, _33592_, _33584_);
  not _39526_ (_33594_, _33575_);
  nor _39527_ (_33595_, _33574_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _39528_ (_33596_, _33595_, _33578_);
  and _39529_ (_33597_, _33596_, _33594_);
  and _39530_ (_33598_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor _39531_ (_33599_, _33598_, _33597_);
  and _39532_ (_33600_, _33599_, _33593_);
  and _39533_ (_33601_, _33554_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and _39534_ (_33602_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _39535_ (_33603_, _33602_, _33601_);
  and _39536_ (_33604_, _33603_, _33600_);
  and _39537_ (_33605_, _33604_, _33591_);
  and _39538_ (_33606_, _33576_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  or _39539_ (_33607_, _33606_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand _39540_ (_33608_, _33606_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and _39541_ (_33609_, _33608_, _33551_);
  and _39542_ (_33610_, _33609_, _33607_);
  not _39543_ (_33611_, _33610_);
  and _39544_ (_33612_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor _39545_ (_33613_, _33612_, _33584_);
  and _39546_ (_33614_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  and _39547_ (_33615_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nor _39548_ (_33616_, _33615_, _33614_);
  and _39549_ (_33617_, _33616_, _33613_);
  and _39550_ (_33618_, _33617_, _33611_);
  not _39551_ (_33619_, _33606_);
  nor _39552_ (_33620_, _33576_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _39553_ (_33621_, _33620_, _33578_);
  and _39554_ (_33622_, _33621_, _33619_);
  not _39555_ (_33623_, _33622_);
  and _39556_ (_33624_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor _39557_ (_33625_, _33624_, _33584_);
  and _39558_ (_33626_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _39559_ (_33627_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor _39560_ (_33628_, _33627_, _33626_);
  and _39561_ (_33629_, _33628_, _33625_);
  and _39562_ (_33630_, _33629_, _33623_);
  not _39563_ (_33631_, _33630_);
  nor _39564_ (_33632_, _33631_, _33618_);
  and _39565_ (_33633_, _33632_, _33605_);
  nor _39566_ (_33634_, _33560_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _39567_ (_33635_, _33634_, _33573_);
  and _39568_ (_33636_, _33635_, _33551_);
  and _39569_ (_33637_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _39570_ (_33638_, _33637_, _33636_);
  and _39571_ (_33639_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and _39572_ (_33640_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and _39573_ (_33641_, _33554_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _39574_ (_33642_, _33641_, _33640_);
  nor _39575_ (_33643_, _33642_, _33639_);
  and _39576_ (_33644_, _33643_, _33638_);
  and _39577_ (_33645_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _39578_ (_33646_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor _39579_ (_33647_, _33646_, _33645_);
  not _39580_ (_33648_, _33574_);
  nor _39581_ (_33649_, _33573_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _39582_ (_33650_, _33649_, _33578_);
  and _39583_ (_33651_, _33650_, _33648_);
  not _39584_ (_33652_, _33651_);
  and _39585_ (_33653_, _33554_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and _39586_ (_33654_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _39587_ (_33655_, _33654_, _33653_);
  and _39588_ (_33656_, _33655_, _33652_);
  and _39589_ (_33657_, _33656_, _33647_);
  not _39590_ (_33658_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _39591_ (_33659_, \oc8051_top_1.oc8051_decoder1.wr , _33129_);
  not _39592_ (_33660_, _33659_);
  nor _39593_ (_33661_, _33660_, _33550_);
  and _39594_ (_33662_, _33661_, _33658_);
  and _39595_ (_33663_, _33662_, _33657_);
  and _39596_ (_33664_, _33663_, _33644_);
  and _39597_ (_33665_, _33664_, _33633_);
  and _39598_ (_33666_, _33665_, _33572_);
  not _39599_ (_33667_, _33666_);
  and _39600_ (_33668_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and _39601_ (_33669_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and _39602_ (_33670_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _33129_);
  and _39603_ (_33671_, _33670_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _39604_ (_33672_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _33129_);
  and _39605_ (_33673_, _33672_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _39606_ (_33674_, _33673_, _33671_);
  not _39607_ (_33675_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  nand _39608_ (_33676_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _33675_);
  nor _39609_ (_33677_, _33676_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not _39610_ (_33678_, _33677_);
  or _39611_ (_33679_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  not _39612_ (_33680_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or _39613_ (_33681_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _33680_);
  and _39614_ (_33682_, _33681_, _33679_);
  not _39615_ (_33683_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and _39616_ (_33684_, _33683_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _39617_ (_33685_, _33684_, _33682_);
  and _39618_ (_33686_, _33685_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  or _39619_ (_33687_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  or _39620_ (_33688_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _33680_);
  and _39621_ (_33689_, _33688_, _33687_);
  nor _39622_ (_33690_, _33683_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _39623_ (_33691_, _33690_, _33689_);
  or _39624_ (_33692_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or _39625_ (_33693_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _33680_);
  and _39626_ (_33694_, _33693_, _33692_);
  nor _39627_ (_33695_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _39628_ (_33696_, _33695_, _33694_);
  or _39629_ (_33697_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  or _39630_ (_33698_, _33680_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and _39631_ (_33699_, _33698_, _33697_);
  and _39632_ (_33700_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand _39633_ (_33701_, _33700_, _33699_);
  and _39634_ (_33702_, _33701_, _33696_);
  and _39635_ (_33703_, _33702_, _33691_);
  nand _39636_ (_33704_, _33703_, _33686_);
  not _39637_ (_33705_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  or _39638_ (_33706_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  or _39639_ (_33707_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _33680_);
  and _39640_ (_33708_, _33707_, _33706_);
  nand _39641_ (_33709_, _33708_, _33684_);
  and _39642_ (_33710_, _33709_, _33705_);
  or _39643_ (_33711_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or _39644_ (_33712_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _33680_);
  and _39645_ (_33713_, _33712_, _33711_);
  nand _39646_ (_33714_, _33713_, _33700_);
  or _39647_ (_33715_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or _39648_ (_33716_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _33680_);
  and _39649_ (_33717_, _33716_, _33715_);
  nand _39650_ (_33718_, _33717_, _33695_);
  or _39651_ (_33719_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or _39652_ (_33720_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _33680_);
  and _39653_ (_33721_, _33720_, _33719_);
  nand _39654_ (_33722_, _33721_, _33690_);
  and _39655_ (_33723_, _33722_, _33718_);
  and _39656_ (_33724_, _33723_, _33714_);
  nand _39657_ (_33725_, _33724_, _33710_);
  nand _39658_ (_33726_, _33725_, _33704_);
  nand _39659_ (_33727_, _33726_, _33676_);
  and _39660_ (_33728_, _33727_, _33678_);
  and _39661_ (_33729_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _39662_ (_33730_, _33729_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _39663_ (_33731_, _33730_);
  and _39664_ (_33732_, _33731_, _33728_);
  and _39665_ (_33733_, _33731_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _39666_ (_33734_, _33733_, _33732_);
  not _39667_ (_33735_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _39668_ (_33736_, _33735_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _39669_ (_33737_, _33736_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _39670_ (_33738_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _39671_ (_33739_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _39672_ (_33740_, _33739_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _39673_ (_33741_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _39674_ (_33742_, _33741_, _33738_);
  nor _39675_ (_33743_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _39676_ (_33744_, _33743_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _39677_ (_33745_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not _39678_ (_33746_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _39679_ (_33747_, _33736_, _33746_);
  and _39680_ (_33748_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor _39681_ (_33749_, _33748_, _33745_);
  and _39682_ (_33750_, _33749_, _33742_);
  and _39683_ (_33751_, _33739_, _33746_);
  not _39684_ (_33752_, _33751_);
  and _39685_ (_33753_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _33675_);
  or _39686_ (_33754_, _33682_, _33753_);
  or _39687_ (_33755_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _39688_ (_33756_, _33755_, _33754_);
  or _39689_ (_33757_, _33756_, _33752_);
  and _39690_ (_33758_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _39691_ (_33759_, _33758_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _39692_ (_33760_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and _39693_ (_33761_, _33758_, _33746_);
  and _39694_ (_33762_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _39695_ (_33763_, _33762_, _33760_);
  and _39696_ (_33764_, _33763_, _33757_);
  and _39697_ (_33765_, _33764_, _33750_);
  not _39698_ (_33766_, _33765_);
  and _39699_ (_33767_, _33766_, _33734_);
  nor _39700_ (_33768_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not _39701_ (_33769_, _33768_);
  or _39702_ (_33770_, _33769_, _33756_);
  and _39703_ (_33771_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _39704_ (_33772_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not _39705_ (_33773_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not _39706_ (_33774_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand _39707_ (_33775_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _33774_);
  nor _39708_ (_33776_, _33775_, _33773_);
  nor _39709_ (_33777_, _33776_, _33772_);
  and _39710_ (_33778_, _33777_, _33770_);
  nor _39711_ (_33779_, _33778_, _33734_);
  or _39712_ (_33780_, _33779_, _33767_);
  and _39713_ (_33781_, _33780_, _33674_);
  nand _39714_ (_33782_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nand _39715_ (_33783_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and _39716_ (_33784_, _33783_, _33782_);
  nand _39717_ (_33785_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _39718_ (_33786_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _39719_ (_33787_, _33786_, _33785_);
  and _39720_ (_33788_, _33787_, _33784_);
  or _39721_ (_33789_, _33689_, _33753_);
  or _39722_ (_33790_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _39723_ (_33791_, _33790_, _33789_);
  or _39724_ (_33792_, _33791_, _33752_);
  nand _39725_ (_33793_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  nand _39726_ (_33794_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _39727_ (_33795_, _33794_, _33793_);
  and _39728_ (_33796_, _33795_, _33792_);
  and _39729_ (_33797_, _33796_, _33788_);
  not _39730_ (_33798_, _33797_);
  and _39731_ (_33799_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and _39732_ (_33800_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  nor _39733_ (_33801_, _33800_, _33799_);
  and _39734_ (_33802_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _39735_ (_33803_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _39736_ (_33804_, _33803_, _33802_);
  and _39737_ (_33805_, _33804_, _33801_);
  or _39738_ (_33806_, _33713_, _33753_);
  or _39739_ (_33807_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _39740_ (_33808_, _33807_, _33806_);
  or _39741_ (_33809_, _33808_, _33752_);
  and _39742_ (_33810_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and _39743_ (_33811_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _39744_ (_33812_, _33811_, _33810_);
  and _39745_ (_33813_, _33812_, _33809_);
  and _39746_ (_33814_, _33813_, _33805_);
  not _39747_ (_33815_, _33814_);
  nand _39748_ (_33816_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand _39749_ (_33817_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _39750_ (_33818_, _33817_, _33816_);
  nand _39751_ (_33819_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nand _39752_ (_33820_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and _39753_ (_33821_, _33820_, _33819_);
  and _39754_ (_33822_, _33821_, _33818_);
  or _39755_ (_33823_, _33721_, _33753_);
  or _39756_ (_33824_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _39757_ (_33825_, _33824_, _33823_);
  or _39758_ (_33826_, _33825_, _33752_);
  nand _39759_ (_33827_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nand _39760_ (_33828_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and _39761_ (_33829_, _33828_, _33827_);
  and _39762_ (_33830_, _33829_, _33826_);
  and _39763_ (_33831_, _33830_, _33822_);
  and _39764_ (_33832_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _39765_ (_33833_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _39766_ (_33834_, _33833_, _33832_);
  and _39767_ (_33835_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and _39768_ (_33836_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor _39769_ (_33837_, _33836_, _33835_);
  and _39770_ (_33838_, _33837_, _33834_);
  or _39771_ (_33839_, _33717_, _33753_);
  or _39772_ (_33840_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and _39773_ (_33841_, _33840_, _33839_);
  and _39774_ (_33842_, _33841_, _33751_);
  and _39775_ (_33843_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and _39776_ (_33844_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _39777_ (_33845_, _33844_, _33843_);
  not _39778_ (_33846_, _33845_);
  nor _39779_ (_33847_, _33846_, _33842_);
  and _39780_ (_33848_, _33847_, _33838_);
  nor _39781_ (_33849_, _33848_, _33831_);
  nand _39782_ (_33850_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nand _39783_ (_33851_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _39784_ (_33852_, _33851_, _33850_);
  nand _39785_ (_33853_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand _39786_ (_33854_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _39787_ (_33855_, _33854_, _33853_);
  and _39788_ (_33856_, _33855_, _33852_);
  or _39789_ (_33857_, _33708_, _33753_);
  or _39790_ (_33858_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _39791_ (_33859_, _33858_, _33857_);
  or _39792_ (_33860_, _33859_, _33752_);
  nand _39793_ (_33861_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nand _39794_ (_33862_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and _39795_ (_33863_, _33862_, _33861_);
  and _39796_ (_33864_, _33863_, _33860_);
  nand _39797_ (_33865_, _33864_, _33856_);
  and _39798_ (_33866_, _33865_, _33849_);
  and _39799_ (_33867_, _33866_, _33815_);
  and _39800_ (_33868_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _39801_ (_33869_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _39802_ (_33870_, _33869_, _33868_);
  and _39803_ (_33871_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _39804_ (_33872_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor _39805_ (_33873_, _33872_, _33871_);
  and _39806_ (_33874_, _33873_, _33870_);
  or _39807_ (_33875_, _33694_, _33753_);
  or _39808_ (_33876_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _39809_ (_33877_, _33876_, _33875_);
  or _39810_ (_33878_, _33877_, _33752_);
  and _39811_ (_33879_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and _39812_ (_33880_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor _39813_ (_33881_, _33880_, _33879_);
  and _39814_ (_33882_, _33881_, _33878_);
  and _39815_ (_33883_, _33882_, _33874_);
  not _39816_ (_33884_, _33883_);
  and _39817_ (_33885_, _33884_, _33867_);
  and _39818_ (_33886_, _33885_, _33798_);
  and _39819_ (_33887_, _33886_, _33734_);
  not _39820_ (_33888_, _33734_);
  nand _39821_ (_33889_, _33848_, _33831_);
  nor _39822_ (_33890_, _33889_, _33865_);
  and _39823_ (_33891_, _33890_, _33814_);
  and _39824_ (_33892_, _33891_, _33883_);
  and _39825_ (_33893_, _33892_, _33797_);
  and _39826_ (_33894_, _33893_, _33888_);
  or _39827_ (_33895_, _33894_, _33887_);
  and _39828_ (_33896_, _33895_, _33766_);
  not _39829_ (_33897_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _39830_ (_33898_, _33672_, _33897_);
  and _39831_ (_33899_, _33671_, _33898_);
  or _39832_ (_33900_, _33895_, _33766_);
  nand _39833_ (_33901_, _33900_, _33899_);
  nor _39834_ (_33902_, _33901_, _33896_);
  nor _39835_ (_33903_, _33902_, _33781_);
  not _39836_ (_33904_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _39837_ (_33905_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _33129_);
  and _39838_ (_33906_, _33905_, _33904_);
  not _39839_ (_33907_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _39840_ (_33908_, _33670_, _33907_);
  and _39841_ (_33909_, _33908_, _33906_);
  not _39842_ (_33910_, _33909_);
  and _39843_ (_33911_, _33778_, _33765_);
  nor _39844_ (_33912_, _33911_, _33910_);
  nor _39845_ (_33913_, _33905_, _33672_);
  and _39846_ (_33914_, _33913_, _33908_);
  nor _39847_ (_33915_, _33778_, _33765_);
  nor _39848_ (_33916_, _33915_, _33911_);
  and _39849_ (_33917_, _33916_, _33914_);
  nor _39850_ (_33918_, _33917_, _33912_);
  not _39851_ (_33919_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _39852_ (_33920_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _33129_);
  and _39853_ (_33921_, _33920_, _33919_);
  and _39854_ (_33922_, _33921_, _33673_);
  and _39855_ (_33923_, _33915_, _33922_);
  and _39856_ (_33924_, _33921_, _33898_);
  and _39857_ (_33925_, _33924_, _33765_);
  nor _39858_ (_33926_, _33925_, _33923_);
  and _39859_ (_33927_, _33908_, _33672_);
  not _39860_ (_33928_, _33927_);
  nor _39861_ (_33929_, _33928_, _33765_);
  nor _39862_ (_33930_, _33670_, _33920_);
  and _39863_ (_33931_, _33930_, _33905_);
  and _39864_ (_33932_, _33921_, _33904_);
  nor _39865_ (_33933_, _33932_, _33931_);
  and _39866_ (_33934_, _33671_, _33904_);
  and _39867_ (_33935_, _33930_, _33913_);
  nor _39868_ (_33936_, _33935_, _33934_);
  and _39869_ (_33937_, _33936_, _33933_);
  nor _39870_ (_33938_, _33937_, _33765_);
  nor _39871_ (_33939_, _33938_, _33929_);
  and _39872_ (_33940_, _33939_, _33926_);
  and _39873_ (_33941_, _33940_, _33918_);
  nand _39874_ (_33942_, _33941_, _33903_);
  and _39875_ (_33943_, _33942_, _33666_);
  nor _39876_ (_33944_, _33943_, _33669_);
  and _39877_ (_33945_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  or _39878_ (_33946_, _33769_, _33791_);
  nand _39879_ (_33947_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  not _39880_ (_33948_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _39881_ (_33949_, _33775_, _33948_);
  and _39882_ (_33950_, _33949_, _33947_);
  and _39883_ (_33951_, _33950_, _33946_);
  nor _39884_ (_33952_, _33951_, _33734_);
  and _39885_ (_33953_, _33798_, _33734_);
  or _39886_ (_33954_, _33953_, _33952_);
  and _39887_ (_33955_, _33954_, _33674_);
  nor _39888_ (_33956_, _33885_, _33888_);
  nor _39889_ (_33957_, _33892_, _33734_);
  nor _39890_ (_33958_, _33957_, _33956_);
  and _39891_ (_33959_, _33958_, _33798_);
  or _39892_ (_33960_, _33958_, _33798_);
  nand _39893_ (_33961_, _33960_, _33899_);
  nor _39894_ (_33962_, _33961_, _33959_);
  nor _39895_ (_33963_, _33962_, _33955_);
  and _39896_ (_33964_, _33951_, _33797_);
  nor _39897_ (_33965_, _33964_, _33910_);
  nor _39898_ (_33966_, _33951_, _33797_);
  nor _39899_ (_33967_, _33966_, _33964_);
  and _39900_ (_33968_, _33967_, _33914_);
  nor _39901_ (_33969_, _33968_, _33965_);
  and _39902_ (_33970_, _33966_, _33922_);
  and _39903_ (_33971_, _33924_, _33797_);
  nor _39904_ (_33972_, _33971_, _33970_);
  nor _39905_ (_33973_, _33928_, _33797_);
  nor _39906_ (_33974_, _33937_, _33797_);
  nor _39907_ (_33975_, _33974_, _33973_);
  and _39908_ (_33976_, _33975_, _33972_);
  and _39909_ (_33977_, _33976_, _33969_);
  nand _39910_ (_33978_, _33977_, _33963_);
  and _39911_ (_33979_, _33978_, _33666_);
  nor _39912_ (_33980_, _33979_, _33945_);
  and _39913_ (_33981_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or _39914_ (_33982_, _33769_, _33877_);
  nand _39915_ (_33983_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not _39916_ (_33984_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _39917_ (_33985_, _33775_, _33984_);
  and _39918_ (_33986_, _33985_, _33983_);
  and _39919_ (_33987_, _33986_, _33982_);
  and _39920_ (_33988_, _33987_, _33883_);
  nor _39921_ (_33989_, _33988_, _33910_);
  nor _39922_ (_33990_, _33987_, _33883_);
  nor _39923_ (_33991_, _33990_, _33988_);
  and _39924_ (_33992_, _33991_, _33914_);
  nor _39925_ (_33993_, _33992_, _33989_);
  nor _39926_ (_33994_, _33928_, _33883_);
  nor _39927_ (_33995_, _33937_, _33883_);
  nor _39928_ (_33996_, _33995_, _33994_);
  and _39929_ (_33997_, _33996_, _33993_);
  nand _39930_ (_33998_, _33867_, _33734_);
  nand _39931_ (_33999_, _33891_, _33888_);
  and _39932_ (_34000_, _33999_, _33998_);
  and _39933_ (_34001_, _34000_, _33883_);
  or _39934_ (_34002_, _34000_, _33883_);
  nand _39935_ (_34003_, _34002_, _33899_);
  or _39936_ (_34004_, _34003_, _34001_);
  and _39937_ (_34005_, _33883_, _33734_);
  not _39938_ (_34006_, _33674_);
  nand _39939_ (_34007_, _33986_, _33982_);
  nor _39940_ (_34008_, _34007_, _33734_);
  or _39941_ (_34009_, _34008_, _34006_);
  nor _39942_ (_34010_, _34009_, _34005_);
  and _39943_ (_34011_, _33990_, _33922_);
  and _39944_ (_34012_, _33924_, _33883_);
  nor _39945_ (_34013_, _34012_, _34011_);
  not _39946_ (_34014_, _34013_);
  nor _39947_ (_34015_, _34014_, _34010_);
  and _39948_ (_34016_, _34015_, _34004_);
  and _39949_ (_34017_, _34016_, _33997_);
  nor _39950_ (_34018_, _34017_, _33667_);
  nor _39951_ (_34019_, _34018_, _33981_);
  nor _39952_ (_34020_, _33928_, _33814_);
  nor _39953_ (_34021_, _33937_, _33814_);
  nor _39954_ (_34022_, _34021_, _34020_);
  or _39955_ (_34023_, _33890_, _33734_);
  or _39956_ (_34024_, _33866_, _33888_);
  and _39957_ (_34025_, _34024_, _34023_);
  or _39958_ (_34026_, _34025_, _33814_);
  nand _39959_ (_34027_, _34025_, _33814_);
  nand _39960_ (_34028_, _34027_, _34026_);
  nand _39961_ (_34029_, _34028_, _33899_);
  or _39962_ (_34030_, _33769_, _33808_);
  nand _39963_ (_34031_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  not _39964_ (_34032_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _39965_ (_34033_, _33775_, _34032_);
  and _39966_ (_34034_, _34033_, _34031_);
  and _39967_ (_34035_, _34034_, _34030_);
  and _39968_ (_34036_, _34035_, _33814_);
  nor _39969_ (_34037_, _34036_, _33910_);
  nor _39970_ (_34038_, _34035_, _33814_);
  or _39971_ (_34039_, _34038_, _34036_);
  not _39972_ (_34040_, _34039_);
  and _39973_ (_34041_, _34040_, _33914_);
  or _39974_ (_34042_, _34041_, _34037_);
  and _39975_ (_34043_, _34038_, _33922_);
  not _39976_ (_34044_, _34043_);
  nor _39977_ (_34045_, _34035_, _34006_);
  and _39978_ (_34046_, _33924_, _33814_);
  nor _39979_ (_34047_, _34046_, _34045_);
  and _39980_ (_34048_, _34047_, _34044_);
  not _39981_ (_34049_, _34048_);
  nor _39982_ (_34050_, _34049_, _34042_);
  and _39983_ (_34051_, _34050_, _34029_);
  and _39984_ (_34052_, _34051_, _34022_);
  nor _39985_ (_34053_, _34052_, _33667_);
  and _39986_ (_34054_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _39987_ (_34055_, _34054_, _34053_);
  and _39988_ (_34056_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  or _39989_ (_34057_, _33769_, _33859_);
  nand _39990_ (_34058_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not _39991_ (_34059_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _39992_ (_34060_, _33775_, _34059_);
  and _39993_ (_34061_, _34060_, _34058_);
  nand _39994_ (_34062_, _34061_, _34057_);
  and _39995_ (_34063_, _34062_, _33674_);
  not _39996_ (_34064_, _33865_);
  not _39997_ (_34065_, _33849_);
  and _39998_ (_34066_, _34065_, _33734_);
  and _39999_ (_34067_, _33889_, _33888_);
  nor _40000_ (_34068_, _34067_, _34066_);
  nand _40001_ (_34069_, _34068_, _34064_);
  or _40002_ (_34070_, _34068_, _34064_);
  nand _40003_ (_34071_, _34070_, _34069_);
  and _40004_ (_34072_, _34071_, _33899_);
  nor _40005_ (_34073_, _34072_, _34063_);
  nor _40006_ (_34074_, _34062_, _33865_);
  nor _40007_ (_34075_, _34074_, _33910_);
  and _40008_ (_34076_, _34062_, _33865_);
  nor _40009_ (_34077_, _34076_, _34074_);
  and _40010_ (_34078_, _34077_, _33914_);
  nor _40011_ (_34079_, _34078_, _34075_);
  and _40012_ (_34080_, _34076_, _33922_);
  and _40013_ (_34081_, _33924_, _34064_);
  nor _40014_ (_34082_, _34081_, _34080_);
  and _40015_ (_34083_, _33927_, _33865_);
  not _40016_ (_34084_, _33937_);
  and _40017_ (_34085_, _34084_, _33865_);
  nor _40018_ (_34086_, _34085_, _34083_);
  and _40019_ (_34087_, _34086_, _34082_);
  and _40020_ (_34088_, _34087_, _34079_);
  nand _40021_ (_34089_, _34088_, _34073_);
  and _40022_ (_34090_, _34089_, _33666_);
  nor _40023_ (_34091_, _34090_, _34056_);
  and _40024_ (_34092_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  or _40025_ (_34093_, _33769_, _33825_);
  nand _40026_ (_34094_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  not _40027_ (_34095_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _40028_ (_34096_, _33775_, _34095_);
  and _40029_ (_34097_, _34096_, _34094_);
  nand _40030_ (_34098_, _34097_, _34093_);
  and _40031_ (_34099_, _34098_, _33674_);
  not _40032_ (_34100_, _33899_);
  and _40033_ (_34101_, _33889_, _34065_);
  nand _40034_ (_34102_, _34101_, _33734_);
  or _40035_ (_34103_, _34101_, _33734_);
  and _40036_ (_34104_, _34103_, _34102_);
  nor _40037_ (_34105_, _34104_, _34100_);
  nor _40038_ (_34106_, _34105_, _34099_);
  not _40039_ (_34107_, _34098_);
  and _40040_ (_34108_, _34107_, _33831_);
  nor _40041_ (_34109_, _34108_, _33910_);
  nor _40042_ (_34110_, _34107_, _33831_);
  nor _40043_ (_34111_, _34110_, _34108_);
  and _40044_ (_34112_, _34111_, _33914_);
  nor _40045_ (_34113_, _34112_, _34109_);
  and _40046_ (_34114_, _34110_, _33922_);
  and _40047_ (_34115_, _33924_, _33831_);
  nor _40048_ (_34116_, _34115_, _34114_);
  nor _40049_ (_34117_, _33928_, _33831_);
  nor _40050_ (_34118_, _33937_, _33831_);
  nor _40051_ (_34119_, _34118_, _34117_);
  and _40052_ (_34120_, _34119_, _34116_);
  and _40053_ (_34121_, _34120_, _34113_);
  nand _40054_ (_34122_, _34121_, _34106_);
  and _40055_ (_34123_, _34122_, _33666_);
  nor _40056_ (_34124_, _34123_, _34092_);
  or _40057_ (_34125_, _33666_, _33549_);
  nand _40058_ (_34126_, _33768_, _33841_);
  nand _40059_ (_34127_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  not _40060_ (_34128_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _40061_ (_34129_, _33775_, _34128_);
  and _40062_ (_34130_, _34129_, _34127_);
  nand _40063_ (_34131_, _34130_, _34126_);
  not _40064_ (_34132_, _34131_);
  and _40065_ (_34133_, _34132_, _33848_);
  nor _40066_ (_34134_, _34132_, _33848_);
  nor _40067_ (_34135_, _34134_, _34133_);
  nand _40068_ (_34136_, _34135_, _33914_);
  nand _40069_ (_34137_, _34134_, _33922_);
  nor _40070_ (_34138_, _34133_, _33910_);
  and _40071_ (_34139_, _34131_, _33674_);
  and _40072_ (_34140_, _33920_, _33898_);
  and _40073_ (_34141_, _34140_, _33848_);
  or _40074_ (_34142_, _34141_, _34139_);
  nor _40075_ (_34143_, _34142_, _34138_);
  and _40076_ (_34144_, _34143_, _34137_);
  and _40077_ (_34145_, _34144_, _34136_);
  and _40078_ (_34146_, _33937_, _33928_);
  or _40079_ (_34147_, _34146_, _33848_);
  and _40080_ (_34148_, _34147_, _34145_);
  not _40081_ (_34149_, _34148_);
  nand _40082_ (_34150_, _34149_, _33666_);
  and _40083_ (_34151_, _34150_, _34125_);
  and _40084_ (_34152_, _34151_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _40085_ (_34153_, _34152_, _34124_);
  and _40086_ (_34154_, _34153_, _34091_);
  and _40087_ (_34155_, _34154_, _34055_);
  and _40088_ (_34156_, _34155_, _34019_);
  and _40089_ (_34157_, _34156_, _33980_);
  and _40090_ (_34158_, _34157_, _33944_);
  nand _40091_ (_34159_, _34158_, _33668_);
  or _40092_ (_34160_, _34158_, _33668_);
  and _40093_ (_34161_, _34160_, _33578_);
  nand _40094_ (_34162_, _34161_, _34159_);
  nor _40095_ (_34163_, _33666_, _33610_);
  and _40096_ (_34164_, _34163_, _34162_);
  and _40097_ (_34165_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _40098_ (_34166_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _40099_ (_34167_, _34166_, _34165_);
  and _40100_ (_34168_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and _40101_ (_34169_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor _40102_ (_34170_, _34169_, _34168_);
  and _40103_ (_34171_, _34170_, _34167_);
  or _40104_ (_34172_, _33699_, _33753_);
  or _40105_ (_34173_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand _40106_ (_34174_, _34173_, _34172_);
  or _40107_ (_34175_, _34174_, _33752_);
  and _40108_ (_34176_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _40109_ (_34177_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor _40110_ (_34178_, _34177_, _34176_);
  and _40111_ (_34179_, _34178_, _34175_);
  and _40112_ (_34180_, _34179_, _34171_);
  and _40113_ (_34181_, _33886_, _33766_);
  nor _40114_ (_34182_, _34181_, _33888_);
  and _40115_ (_34183_, _33797_, _33765_);
  and _40116_ (_34184_, _34183_, _33892_);
  nor _40117_ (_34185_, _34184_, _33734_);
  or _40118_ (_34186_, _34185_, _34182_);
  and _40119_ (_34187_, _34186_, _34180_);
  nor _40120_ (_34188_, _34186_, _34180_);
  nor _40121_ (_34189_, _34188_, _34187_);
  and _40122_ (_34190_, _34189_, _33899_);
  or _40123_ (_34191_, _33769_, _34174_);
  and _40124_ (_34192_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not _40125_ (_34193_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _40126_ (_34194_, _33775_, _34193_);
  nor _40127_ (_34195_, _34194_, _34192_);
  and _40128_ (_34196_, _34195_, _34191_);
  not _40129_ (_34197_, _34196_);
  nor _40130_ (_34198_, _34197_, _33734_);
  not _40131_ (_34199_, _34198_);
  and _40132_ (_34200_, _33734_, _34180_);
  nor _40133_ (_34201_, _34200_, _34006_);
  and _40134_ (_34202_, _34201_, _34199_);
  nor _40135_ (_34203_, _34202_, _34190_);
  and _40136_ (_34204_, _34196_, _34180_);
  nor _40137_ (_34205_, _34204_, _33910_);
  nor _40138_ (_34206_, _34196_, _34180_);
  nor _40139_ (_34207_, _34206_, _34204_);
  and _40140_ (_34208_, _34207_, _33914_);
  nor _40141_ (_34209_, _34208_, _34205_);
  and _40142_ (_34210_, _33922_, _34206_);
  and _40143_ (_34211_, _33924_, _34180_);
  nor _40144_ (_34212_, _34211_, _34210_);
  not _40145_ (_34213_, _33934_);
  nor _40146_ (_34214_, _34213_, _34180_);
  nor _40147_ (_34215_, _33927_, _33935_);
  and _40148_ (_34216_, _34215_, _33933_);
  nor _40149_ (_34217_, _34216_, _34180_);
  nor _40150_ (_34218_, _34217_, _34214_);
  and _40151_ (_34219_, _34218_, _34212_);
  and _40152_ (_34220_, _34219_, _34209_);
  and _40153_ (_34221_, _34220_, _34203_);
  and _40154_ (_34222_, _34221_, _33666_);
  nor _40155_ (_34223_, _34222_, _34164_);
  nand _40156_ (_34224_, _34223_, _33534_);
  not _40157_ (_34225_, _33532_);
  and _40158_ (_34226_, _34225_, _33474_);
  not _40159_ (_34227_, _33604_);
  and _40160_ (_34228_, _33571_, _33558_);
  and _40161_ (_34229_, _34228_, _33644_);
  and _40162_ (_34230_, _34229_, _33663_);
  nor _40163_ (_34231_, _33630_, _33618_);
  not _40164_ (_34232_, _33591_);
  nor _40165_ (_34233_, _33604_, _34232_);
  and _40166_ (_34234_, _34233_, _34231_);
  and _40167_ (_34235_, _34234_, _34230_);
  not _40168_ (_34236_, _34235_);
  and _40169_ (_34237_, _34236_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor _40170_ (_34238_, _34236_, _34017_);
  nor _40171_ (_34239_, _34238_, _34237_);
  nor _40172_ (_34240_, _34239_, _34227_);
  and _40173_ (_34241_, _34239_, _34227_);
  nor _40174_ (_34242_, _34241_, _34240_);
  nand _40175_ (_34243_, _33559_, _33226_);
  or _40176_ (_34244_, _33559_, _33226_);
  and _40177_ (_34245_, _34244_, _34243_);
  not _40178_ (_34246_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _40179_ (_34247_, _33659_, _34246_);
  not _40180_ (_34248_, _34247_);
  and _40181_ (_34249_, _33630_, _33618_);
  and _40182_ (_34250_, _34249_, _33605_);
  not _40183_ (_34251_, _33657_);
  and _40184_ (_34252_, _33644_, _33571_);
  and _40185_ (_34253_, _34252_, _33559_);
  and _40186_ (_34254_, _34253_, _34251_);
  and _40187_ (_34255_, _34254_, _34250_);
  not _40188_ (_34256_, _34255_);
  and _40189_ (_34257_, _34229_, _33657_);
  and _40190_ (_34258_, _34250_, _34257_);
  and _40191_ (_34259_, _34253_, _33657_);
  and _40192_ (_34260_, _34250_, _34259_);
  nor _40193_ (_34261_, _34260_, _34258_);
  and _40194_ (_34262_, _34229_, _34251_);
  and _40195_ (_34263_, _34262_, _34250_);
  not _40196_ (_34264_, _34263_);
  and _40197_ (_34265_, _34264_, _34261_);
  and _40198_ (_34266_, _34265_, _34256_);
  and _40199_ (_34267_, _34249_, _34233_);
  and _40200_ (_34268_, _34267_, _34257_);
  and _40201_ (_34269_, _34267_, _34259_);
  nor _40202_ (_34270_, _34269_, _34268_);
  and _40203_ (_34271_, _34267_, _34262_);
  not _40204_ (_34272_, _34271_);
  and _40205_ (_34273_, _34272_, _34270_);
  and _40206_ (_34274_, _34273_, _34266_);
  or _40207_ (_34275_, _34274_, _34248_);
  and _40208_ (_34276_, _34254_, _34247_);
  and _40209_ (_34277_, _34276_, _34267_);
  not _40210_ (_34278_, _34277_);
  and _40211_ (_34279_, _34278_, _34275_);
  nor _40212_ (_34280_, _34279_, _34245_);
  and _40213_ (_34281_, _34236_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _40214_ (_34282_, _34236_, _34052_);
  nor _40215_ (_34283_, _34282_, _34281_);
  and _40216_ (_34284_, _34283_, _34251_);
  nor _40217_ (_34285_, _34283_, _34251_);
  nor _40218_ (_34286_, _34285_, _34284_);
  and _40219_ (_34287_, _34286_, _34280_);
  and _40220_ (_34288_, _34287_, _34242_);
  and _40221_ (_34289_, _34283_, _33226_);
  and _40222_ (_34290_, _34289_, _34239_);
  nand _40223_ (_34291_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _40224_ (_34292_, _34283_, _33464_);
  and _40225_ (_34293_, _34292_, _34239_);
  nand _40226_ (_34294_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _40227_ (_34295_, _34294_, _34291_);
  nor _40228_ (_34296_, _34283_, _33464_);
  and _40229_ (_34297_, _34296_, _34239_);
  nand _40230_ (_34298_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor _40231_ (_34299_, _34283_, _33226_);
  and _40232_ (_34300_, _34299_, _34239_);
  nand _40233_ (_34301_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _40234_ (_34302_, _34301_, _34298_);
  and _40235_ (_34303_, _34302_, _34295_);
  not _40236_ (_34304_, _34239_);
  and _40237_ (_34305_, _34299_, _34304_);
  nand _40238_ (_34306_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and _40239_ (_34307_, _34296_, _34304_);
  nand _40240_ (_34308_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and _40241_ (_34309_, _34308_, _34306_);
  and _40242_ (_34310_, _34289_, _34304_);
  nand _40243_ (_34311_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _40244_ (_34312_, _34292_, _34304_);
  nand _40245_ (_34313_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _40246_ (_34314_, _34313_, _34311_);
  and _40247_ (_34315_, _34314_, _34309_);
  and _40248_ (_34316_, _34315_, _34303_);
  nor _40249_ (_34317_, _34316_, _34288_);
  not _40250_ (_34318_, _34221_);
  and _40251_ (_34319_, _34288_, _34318_);
  or _40252_ (_34320_, _34319_, _34317_);
  nand _40253_ (_34321_, _34320_, _34226_);
  and _40254_ (_34322_, _33532_, _33499_);
  not _40255_ (_34323_, _34322_);
  or _40256_ (_34324_, _34323_, _33474_);
  not _40257_ (_34325_, _33135_);
  and _40258_ (_34326_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and _40259_ (_34327_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _40260_ (_34328_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _40261_ (_34329_, _34328_, _34327_);
  and _40262_ (_34330_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _40263_ (_34331_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _40264_ (_34332_, _34331_, _34330_);
  and _40265_ (_34333_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not _40266_ (_34334_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _40267_ (_34335_, _33146_, _34334_);
  nor _40268_ (_34336_, _34335_, _34333_);
  and _40269_ (_34337_, _34336_, _34332_);
  and _40270_ (_34338_, _34337_, _34329_);
  and _40271_ (_34339_, _33141_, _33135_);
  not _40272_ (_34340_, _34339_);
  nor _40273_ (_34341_, _34340_, _34338_);
  nor _40274_ (_34342_, _34341_, _34326_);
  or _40275_ (_34343_, _34342_, _34324_);
  and _40276_ (_34344_, _34343_, _33499_);
  and _40277_ (_34345_, _34344_, _34321_);
  nand _40278_ (_34346_, _34345_, _34224_);
  and _40279_ (_34347_, _33376_, _33385_);
  and _40280_ (_34348_, _34347_, _33464_);
  and _40281_ (_34349_, _33423_, _33465_);
  or _40282_ (_34350_, _34349_, _34348_);
  and _40283_ (_34351_, _33437_, _33465_);
  nor _40284_ (_34352_, _34351_, _34350_);
  and _40285_ (_34353_, _34352_, _33362_);
  and _40286_ (_34354_, _33418_, _33385_);
  and _40287_ (_34355_, _34354_, _33464_);
  and _40288_ (_34356_, _33397_, _33465_);
  or _40289_ (_34357_, _34356_, _34355_);
  and _40290_ (_34358_, _33388_, _33465_);
  and _40291_ (_34359_, _33465_, _33408_);
  or _40292_ (_34360_, _33416_, _33405_);
  or _40293_ (_34361_, _34360_, _34359_);
  or _40294_ (_34362_, _34361_, _34358_);
  nor _40295_ (_34363_, _34362_, _34357_);
  and _40296_ (_34364_, _34363_, _34353_);
  nor _40297_ (_34365_, _34364_, _33477_);
  and _40298_ (_34366_, _33360_, _33353_);
  not _40299_ (_34367_, _33458_);
  nor _40300_ (_34368_, _34367_, _34366_);
  nor _40301_ (_34369_, _34368_, _34365_);
  or _40302_ (_34370_, _34369_, _34346_);
  and _40303_ (_34371_, _34226_, _33499_);
  not _40304_ (_34372_, _34371_);
  and _40305_ (_34373_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _40306_ (_34374_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor _40307_ (_34375_, _34374_, _34373_);
  and _40308_ (_34376_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _40309_ (_34377_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor _40310_ (_34378_, _34377_, _34376_);
  and _40311_ (_34379_, _34378_, _34375_);
  and _40312_ (_34380_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _40313_ (_34381_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor _40314_ (_34382_, _34381_, _34380_);
  and _40315_ (_34383_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _40316_ (_34384_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _40317_ (_34385_, _34384_, _34383_);
  and _40318_ (_34386_, _34385_, _34382_);
  and _40319_ (_34387_, _34386_, _34379_);
  nor _40320_ (_34388_, _34387_, _34288_);
  not _40321_ (_34389_, _34052_);
  and _40322_ (_34390_, _34288_, _34389_);
  nor _40323_ (_34391_, _34390_, _34388_);
  or _40324_ (_34392_, _34391_, _34372_);
  not _40325_ (_34393_, _34283_);
  and _40326_ (_34394_, _34322_, _33474_);
  and _40327_ (_34395_, _34394_, _34393_);
  nor _40328_ (_34396_, _34154_, _34055_);
  or _40329_ (_34397_, _34396_, _34155_);
  nand _40330_ (_34398_, _34397_, _33578_);
  nand _40331_ (_34399_, _34398_, _33652_);
  and _40332_ (_34400_, _34399_, _33667_);
  or _40333_ (_34401_, _34400_, _34053_);
  nand _40334_ (_34402_, _34401_, _33534_);
  and _40335_ (_34403_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and _40336_ (_34404_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  not _40337_ (_34405_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _40338_ (_34406_, _33146_, _34405_);
  nor _40339_ (_34407_, _34406_, _34404_);
  and _40340_ (_34408_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _40341_ (_34409_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _40342_ (_34410_, _34409_, _34408_);
  and _40343_ (_34411_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _40344_ (_34412_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _40345_ (_34413_, _34412_, _34411_);
  and _40346_ (_34414_, _34413_, _34410_);
  and _40347_ (_34415_, _34414_, _34407_);
  nor _40348_ (_34416_, _34415_, _34340_);
  nor _40349_ (_34417_, _34416_, _34403_);
  or _40350_ (_34418_, _34417_, _34324_);
  nand _40351_ (_34419_, _34418_, _34402_);
  nor _40352_ (_34420_, _34419_, _34395_);
  and _40353_ (_34421_, _34420_, _34392_);
  or _40354_ (_34422_, _34421_, _34370_);
  not _40355_ (_34423_, _34369_);
  and _40356_ (_34424_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _40357_ (_34425_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor _40358_ (_34426_, _34425_, _34424_);
  and _40359_ (_34427_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _40360_ (_34428_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor _40361_ (_34429_, _34428_, _34427_);
  and _40362_ (_34430_, _34429_, _34426_);
  and _40363_ (_34431_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _40364_ (_34432_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor _40365_ (_34433_, _34432_, _34431_);
  and _40366_ (_34434_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _40367_ (_34435_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor _40368_ (_34436_, _34435_, _34434_);
  and _40369_ (_34437_, _34436_, _34433_);
  and _40370_ (_34438_, _34437_, _34430_);
  nor _40371_ (_34439_, _34438_, _34288_);
  and _40372_ (_34440_, _34288_, _34149_);
  nor _40373_ (_34441_, _34440_, _34439_);
  or _40374_ (_34442_, _34441_, _34372_);
  and _40375_ (_34443_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and _40376_ (_34444_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  not _40377_ (_34445_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _40378_ (_34446_, _33146_, _34445_);
  nor _40379_ (_34447_, _34446_, _34444_);
  and _40380_ (_34448_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _40381_ (_34449_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _40382_ (_34450_, _34449_, _34448_);
  and _40383_ (_34451_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _40384_ (_34452_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _40385_ (_34453_, _34452_, _34451_);
  and _40386_ (_34454_, _34453_, _34450_);
  and _40387_ (_34455_, _34454_, _34447_);
  nor _40388_ (_34456_, _34455_, _34340_);
  nor _40389_ (_34457_, _34456_, _34443_);
  nor _40390_ (_34458_, _34457_, _34324_);
  not _40391_ (_34459_, _33534_);
  nor _40392_ (_34460_, _34151_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor _40393_ (_34461_, _34460_, _34152_);
  nor _40394_ (_34462_, _34461_, _33551_);
  nor _40395_ (_34463_, _34462_, _33552_);
  nor _40396_ (_34464_, _34463_, _33666_);
  not _40397_ (_34465_, _34464_);
  and _40398_ (_34466_, _34465_, _34150_);
  or _40399_ (_34467_, _34466_, _34459_);
  nand _40400_ (_34468_, _34394_, _33226_);
  nand _40401_ (_34469_, _34468_, _34467_);
  nor _40402_ (_34470_, _34469_, _34458_);
  and _40403_ (_34471_, _34470_, _34442_);
  or _40404_ (_34472_, _34471_, _34423_);
  nand _40405_ (_34473_, _34472_, _34422_);
  and _40406_ (_34474_, _33618_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _40407_ (_34475_, _34474_, _34251_);
  nor _40408_ (_34476_, _33558_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _40409_ (_34477_, _34476_, _34475_);
  nor _40410_ (_34478_, _34477_, _34473_);
  and _40411_ (_34479_, _34477_, _34473_);
  nor _40412_ (_34480_, _34479_, _34478_);
  and _40413_ (_34481_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and _40414_ (_34482_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  not _40415_ (_34483_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _40416_ (_34484_, _33146_, _34483_);
  nor _40417_ (_34485_, _34484_, _34482_);
  and _40418_ (_34486_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _40419_ (_34487_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _40420_ (_34488_, _34487_, _34486_);
  and _40421_ (_34489_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _40422_ (_34490_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _40423_ (_34491_, _34490_, _34489_);
  and _40424_ (_34492_, _34491_, _34488_);
  and _40425_ (_34493_, _34492_, _34485_);
  nor _40426_ (_34494_, _34493_, _34340_);
  nor _40427_ (_34495_, _34494_, _34481_);
  nor _40428_ (_34496_, _34495_, _34324_);
  and _40429_ (_34497_, _34394_, _34304_);
  nor _40430_ (_34498_, _34497_, _34496_);
  and _40431_ (_34499_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _40432_ (_34500_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _40433_ (_34501_, _34500_, _34499_);
  and _40434_ (_34502_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _40435_ (_34503_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor _40436_ (_34504_, _34503_, _34502_);
  and _40437_ (_34505_, _34504_, _34501_);
  and _40438_ (_34506_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and _40439_ (_34507_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor _40440_ (_34508_, _34507_, _34506_);
  and _40441_ (_34509_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _40442_ (_34510_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor _40443_ (_34511_, _34510_, _34509_);
  and _40444_ (_34512_, _34511_, _34508_);
  and _40445_ (_34513_, _34512_, _34505_);
  nor _40446_ (_34514_, _34513_, _34288_);
  not _40447_ (_34515_, _34017_);
  and _40448_ (_34516_, _34288_, _34515_);
  nor _40449_ (_34517_, _34516_, _34514_);
  or _40450_ (_34518_, _34517_, _34372_);
  and _40451_ (_34519_, _33532_, _33500_);
  nor _40452_ (_34520_, _34155_, _34019_);
  or _40453_ (_34521_, _34520_, _34156_);
  and _40454_ (_34522_, _34521_, _33578_);
  or _40455_ (_34523_, _34522_, _33597_);
  and _40456_ (_34524_, _34523_, _33667_);
  or _40457_ (_34525_, _34524_, _34018_);
  and _40458_ (_34526_, _34525_, _33534_);
  nor _40459_ (_34527_, _34526_, _34519_);
  and _40460_ (_34528_, _34527_, _34518_);
  and _40461_ (_34529_, _34528_, _34498_);
  or _40462_ (_34530_, _34529_, _34370_);
  and _40463_ (_34531_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _40464_ (_34532_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor _40465_ (_34533_, _34532_, _34531_);
  and _40466_ (_34534_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _40467_ (_34535_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor _40468_ (_34536_, _34535_, _34534_);
  and _40469_ (_34537_, _34536_, _34533_);
  and _40470_ (_34538_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _40471_ (_34539_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor _40472_ (_34540_, _34539_, _34538_);
  and _40473_ (_34541_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _40474_ (_34542_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _40475_ (_34543_, _34542_, _34541_);
  and _40476_ (_34544_, _34543_, _34540_);
  and _40477_ (_34545_, _34544_, _34537_);
  nor _40478_ (_34546_, _34545_, _34288_);
  and _40479_ (_34547_, _34288_, _34122_);
  nor _40480_ (_34548_, _34547_, _34546_);
  nor _40481_ (_34549_, _34548_, _34372_);
  not _40482_ (_34550_, _34549_);
  and _40483_ (_34551_, _34226_, _33500_);
  nor _40484_ (_34552_, _34152_, _34124_);
  nor _40485_ (_34553_, _34552_, _34153_);
  nor _40486_ (_34554_, _34553_, _33551_);
  nor _40487_ (_34555_, _34554_, _33563_);
  nor _40488_ (_34556_, _34555_, _33666_);
  nor _40489_ (_34557_, _34556_, _34123_);
  not _40490_ (_34558_, _34557_);
  and _40491_ (_34559_, _34558_, _33534_);
  nor _40492_ (_34560_, _34559_, _34551_);
  and _40493_ (_34561_, _34394_, _33250_);
  and _40494_ (_34562_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and _40495_ (_34563_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _40496_ (_34564_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _40497_ (_34565_, _34564_, _34563_);
  and _40498_ (_34566_, _33236_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and _40499_ (_34567_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _40500_ (_34568_, _34567_, _34566_);
  and _40501_ (_34569_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _40502_ (_34570_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _40503_ (_34571_, _34570_, _34569_);
  and _40504_ (_34572_, _34571_, _34568_);
  and _40505_ (_34573_, _34572_, _34565_);
  nor _40506_ (_34574_, _34573_, _34340_);
  nor _40507_ (_34575_, _34574_, _34562_);
  nor _40508_ (_34576_, _34575_, _34324_);
  nor _40509_ (_34577_, _34576_, _34561_);
  and _40510_ (_34578_, _34577_, _34560_);
  and _40511_ (_34579_, _34578_, _34550_);
  or _40512_ (_34580_, _34579_, _34423_);
  and _40513_ (_34581_, _34580_, _34530_);
  and _40514_ (_34582_, _34474_, _34227_);
  nor _40515_ (_34583_, _33571_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _40516_ (_34584_, _34583_, _34582_);
  and _40517_ (_34585_, _34584_, _34581_);
  nor _40518_ (_34586_, _34584_, _34581_);
  or _40519_ (_34587_, _34586_, _34585_);
  and _40520_ (_34588_, _34587_, _34480_);
  and _40521_ (_34589_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and _40522_ (_34590_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  not _40523_ (_34591_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _40524_ (_34592_, _33146_, _34591_);
  nor _40525_ (_34593_, _34592_, _34590_);
  and _40526_ (_34594_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _40527_ (_34595_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _40528_ (_34596_, _34595_, _34594_);
  and _40529_ (_34597_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _40530_ (_34598_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _40531_ (_34599_, _34598_, _34597_);
  and _40532_ (_34600_, _34599_, _34596_);
  and _40533_ (_34601_, _34600_, _34593_);
  nor _40534_ (_34602_, _34601_, _34340_);
  nor _40535_ (_34603_, _34602_, _34589_);
  nor _40536_ (_34604_, _34603_, _34324_);
  nor _40537_ (_34605_, _34225_, _33474_);
  not _40538_ (_34606_, _34605_);
  nor _40539_ (_34607_, _34226_, _33499_);
  and _40540_ (_34608_, _34607_, _34606_);
  or _40541_ (_34609_, _34608_, _34604_);
  nor _40542_ (_34610_, _34156_, _33980_);
  nor _40543_ (_34611_, _34610_, _34157_);
  nor _40544_ (_34612_, _34611_, _33551_);
  nor _40545_ (_34613_, _34612_, _33581_);
  nor _40546_ (_34614_, _34613_, _33666_);
  nor _40547_ (_34615_, _34614_, _33979_);
  nor _40548_ (_34616_, _34615_, _34459_);
  and _40549_ (_34617_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _40550_ (_34618_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor _40551_ (_34619_, _34618_, _34617_);
  and _40552_ (_34620_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and _40553_ (_34621_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor _40554_ (_34622_, _34621_, _34620_);
  and _40555_ (_34623_, _34622_, _34619_);
  and _40556_ (_34624_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _40557_ (_34625_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _40558_ (_34626_, _34625_, _34624_);
  and _40559_ (_34627_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _40560_ (_34628_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor _40561_ (_34629_, _34628_, _34627_);
  and _40562_ (_34630_, _34629_, _34626_);
  and _40563_ (_34631_, _34630_, _34623_);
  nor _40564_ (_34632_, _34631_, _34288_);
  and _40565_ (_34633_, _34288_, _33978_);
  nor _40566_ (_34634_, _34633_, _34632_);
  nor _40567_ (_34635_, _34634_, _34372_);
  or _40568_ (_34636_, _34635_, _34616_);
  nor _40569_ (_34637_, _34636_, _34609_);
  and _40570_ (_34638_, _34637_, _34370_);
  nor _40571_ (_34639_, _34474_, _34232_);
  not _40572_ (_34640_, _34639_);
  nor _40573_ (_34641_, _34640_, _34638_);
  not _40574_ (_34642_, _34641_);
  not _40575_ (_34643_, _34370_);
  nor _40576_ (_34644_, _34157_, _33944_);
  nor _40577_ (_34645_, _34644_, _34158_);
  nor _40578_ (_34646_, _34645_, _33551_);
  nor _40579_ (_34647_, _34646_, _33622_);
  nor _40580_ (_34648_, _34647_, _33666_);
  nor _40581_ (_34649_, _34648_, _33943_);
  nor _40582_ (_34650_, _34649_, _34459_);
  not _40583_ (_34651_, _34650_);
  and _40584_ (_34652_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _40585_ (_34653_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor _40586_ (_34654_, _34653_, _34652_);
  and _40587_ (_34655_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and _40588_ (_34656_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor _40589_ (_34657_, _34656_, _34655_);
  and _40590_ (_34658_, _34657_, _34654_);
  and _40591_ (_34659_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _40592_ (_34660_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor _40593_ (_34661_, _34660_, _34659_);
  and _40594_ (_34662_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and _40595_ (_34663_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor _40596_ (_34664_, _34663_, _34662_);
  and _40597_ (_34665_, _34664_, _34661_);
  and _40598_ (_34666_, _34665_, _34658_);
  nor _40599_ (_34667_, _34666_, _34288_);
  and _40600_ (_34668_, _34288_, _33942_);
  nor _40601_ (_34669_, _34668_, _34667_);
  nor _40602_ (_34670_, _34669_, _34372_);
  and _40603_ (_34671_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and _40604_ (_34672_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  not _40605_ (_34673_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _40606_ (_34674_, _33146_, _34673_);
  nor _40607_ (_34675_, _34674_, _34672_);
  and _40608_ (_34676_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _40609_ (_34677_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _40610_ (_34678_, _34677_, _34676_);
  and _40611_ (_34679_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _40612_ (_34680_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _40613_ (_34681_, _34680_, _34679_);
  and _40614_ (_34682_, _34681_, _34678_);
  and _40615_ (_34683_, _34682_, _34675_);
  nor _40616_ (_34684_, _34683_, _34340_);
  nor _40617_ (_34685_, _34684_, _34671_);
  not _40618_ (_34686_, _34685_);
  and _40619_ (_34687_, _34686_, _34605_);
  nor _40620_ (_34688_, _34607_, _34687_);
  not _40621_ (_34689_, _34688_);
  nor _40622_ (_34690_, _34689_, _34670_);
  and _40623_ (_34691_, _34690_, _34651_);
  nor _40624_ (_34692_, _34691_, _34643_);
  nor _40625_ (_34693_, _34474_, _33630_);
  not _40626_ (_34694_, _34693_);
  and _40627_ (_34695_, _34694_, _34692_);
  nor _40628_ (_34696_, _34694_, _34692_);
  nor _40629_ (_34697_, _34696_, _34695_);
  and _40630_ (_34698_, _34697_, _34642_);
  not _40631_ (_34699_, _34529_);
  and _40632_ (_34700_, _34699_, _34370_);
  nor _40633_ (_34701_, _34474_, _33604_);
  not _40634_ (_34702_, _34701_);
  and _40635_ (_34703_, _34702_, _34700_);
  and _40636_ (_34704_, _34640_, _34638_);
  nor _40637_ (_34705_, _34704_, _34703_);
  not _40638_ (_34706_, _33618_);
  and _40639_ (_34707_, _34346_, _34706_);
  nor _40640_ (_34708_, _34346_, _34706_);
  nor _40641_ (_34709_, _34708_, _34707_);
  not _40642_ (_34710_, _34709_);
  and _40643_ (_34711_, _34710_, _34705_);
  and _40644_ (_34712_, _34711_, _34698_);
  and _40645_ (_34713_, _34712_, _34588_);
  and _40646_ (_34714_, _34474_, _33631_);
  nor _40647_ (_34715_, _34474_, _33657_);
  nor _40648_ (_34716_, _34715_, _34714_);
  and _40649_ (_34717_, _34691_, _34643_);
  and _40650_ (_34718_, _34421_, _34370_);
  nor _40651_ (_34719_, _34718_, _34717_);
  and _40652_ (_34720_, _34719_, _34716_);
  nor _40653_ (_34721_, _34719_, _34716_);
  or _40654_ (_34722_, _34721_, _34720_);
  nor _40655_ (_34723_, _34637_, _34370_);
  and _40656_ (_34724_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _40657_ (_34725_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor _40658_ (_34726_, _34725_, _34724_);
  and _40659_ (_34727_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _40660_ (_34728_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor _40661_ (_34729_, _34728_, _34727_);
  and _40662_ (_34730_, _34729_, _34726_);
  and _40663_ (_34731_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and _40664_ (_34732_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor _40665_ (_34733_, _34732_, _34731_);
  and _40666_ (_34734_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and _40667_ (_34735_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _40668_ (_34736_, _34735_, _34734_);
  and _40669_ (_34737_, _34736_, _34733_);
  and _40670_ (_34738_, _34737_, _34730_);
  nor _40671_ (_34739_, _34738_, _34288_);
  and _40672_ (_34740_, _34288_, _34089_);
  nor _40673_ (_34741_, _34740_, _34739_);
  nor _40674_ (_34742_, _34741_, _34372_);
  and _40675_ (_34743_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and _40676_ (_34744_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _40677_ (_34745_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _40678_ (_34746_, _34745_, _34744_);
  not _40679_ (_34747_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _40680_ (_34748_, _33146_, _34747_);
  and _40681_ (_34749_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _40682_ (_34750_, _34749_, _34748_);
  and _40683_ (_34751_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _40684_ (_34752_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _40685_ (_34753_, _34752_, _34751_);
  and _40686_ (_34754_, _34753_, _34750_);
  and _40687_ (_34755_, _34754_, _34746_);
  nor _40688_ (_34756_, _34755_, _34340_);
  nor _40689_ (_34757_, _34756_, _34743_);
  nor _40690_ (_34758_, _34757_, _34324_);
  nor _40691_ (_34759_, _34758_, _34742_);
  and _40692_ (_34760_, _34394_, _33177_);
  nor _40693_ (_34761_, _34153_, _34091_);
  nor _40694_ (_34762_, _34761_, _34154_);
  nor _40695_ (_34763_, _34762_, _33551_);
  nor _40696_ (_34764_, _34763_, _33636_);
  nor _40697_ (_34765_, _34764_, _33666_);
  nor _40698_ (_34766_, _34765_, _34090_);
  not _40699_ (_34767_, _34766_);
  and _40700_ (_34768_, _34767_, _33534_);
  nor _40701_ (_34769_, _34768_, _34760_);
  and _40702_ (_34770_, _34769_, _34759_);
  nor _40703_ (_34771_, _34770_, _34423_);
  nor _40704_ (_34772_, _34771_, _34723_);
  and _40705_ (_34773_, _34474_, _34232_);
  nor _40706_ (_34774_, _33644_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _40707_ (_34775_, _34774_, _34773_);
  not _40708_ (_34776_, _34775_);
  and _40709_ (_34777_, _34776_, _34772_);
  nor _40710_ (_34778_, _34776_, _34772_);
  nor _40711_ (_34779_, _34778_, _34777_);
  not _40712_ (_34780_, _34779_);
  nor _40713_ (_34781_, _34780_, _34722_);
  nor _40714_ (_34782_, _34702_, _34700_);
  nor _40715_ (_34783_, _33618_, _33550_);
  nor _40716_ (_34784_, _34783_, _33660_);
  not _40717_ (_34785_, _34784_);
  nor _40718_ (_34786_, _34785_, _34782_);
  and _40719_ (_34787_, _34786_, _34781_);
  and _40720_ (_34788_, _34787_, _34713_);
  not _40721_ (_34789_, _34700_);
  not _40722_ (_34790_, _34772_);
  and _40723_ (_34791_, _34472_, _34422_);
  and _40724_ (_34792_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and _40725_ (_34793_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or _40726_ (_34794_, _34793_, _34792_);
  and _40727_ (_34795_, _34794_, _34581_);
  not _40728_ (_34796_, _34581_);
  and _40729_ (_34797_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and _40730_ (_34798_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or _40731_ (_34799_, _34798_, _34797_);
  and _40732_ (_34800_, _34799_, _34796_);
  or _40733_ (_34801_, _34800_, _34795_);
  or _40734_ (_34802_, _34801_, _34790_);
  not _40735_ (_34803_, _34719_);
  and _40736_ (_34804_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  and _40737_ (_34805_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or _40738_ (_34806_, _34805_, _34804_);
  and _40739_ (_34807_, _34806_, _34581_);
  and _40740_ (_34808_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and _40741_ (_34809_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or _40742_ (_34810_, _34809_, _34808_);
  and _40743_ (_34811_, _34810_, _34796_);
  or _40744_ (_34812_, _34811_, _34807_);
  or _40745_ (_34813_, _34812_, _34772_);
  and _40746_ (_34814_, _34813_, _34803_);
  and _40747_ (_34815_, _34814_, _34802_);
  or _40748_ (_34816_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or _40749_ (_34817_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and _40750_ (_34818_, _34817_, _34816_);
  and _40751_ (_34819_, _34818_, _34581_);
  or _40752_ (_34820_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or _40753_ (_34821_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and _40754_ (_34822_, _34821_, _34820_);
  and _40755_ (_34823_, _34822_, _34796_);
  or _40756_ (_34824_, _34823_, _34819_);
  or _40757_ (_34825_, _34824_, _34790_);
  or _40758_ (_34826_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or _40759_ (_34827_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and _40760_ (_34828_, _34827_, _34826_);
  and _40761_ (_34829_, _34828_, _34581_);
  or _40762_ (_34830_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or _40763_ (_34831_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  and _40764_ (_34832_, _34831_, _34830_);
  and _40765_ (_34833_, _34832_, _34796_);
  or _40766_ (_34834_, _34833_, _34829_);
  or _40767_ (_34835_, _34834_, _34772_);
  and _40768_ (_34836_, _34835_, _34719_);
  and _40769_ (_34837_, _34836_, _34825_);
  or _40770_ (_34838_, _34837_, _34815_);
  or _40771_ (_34839_, _34838_, _34789_);
  not _40772_ (_34840_, _34638_);
  and _40773_ (_34841_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and _40774_ (_34842_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or _40775_ (_34843_, _34842_, _34841_);
  and _40776_ (_34844_, _34843_, _34581_);
  and _40777_ (_34845_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and _40778_ (_34846_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or _40779_ (_34847_, _34846_, _34845_);
  and _40780_ (_34848_, _34847_, _34796_);
  or _40781_ (_34849_, _34848_, _34844_);
  or _40782_ (_34850_, _34849_, _34790_);
  and _40783_ (_34851_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and _40784_ (_34852_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or _40785_ (_34853_, _34852_, _34851_);
  and _40786_ (_34854_, _34853_, _34581_);
  and _40787_ (_34855_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and _40788_ (_34856_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or _40789_ (_34857_, _34856_, _34855_);
  and _40790_ (_34858_, _34857_, _34796_);
  or _40791_ (_34859_, _34858_, _34854_);
  or _40792_ (_34860_, _34859_, _34772_);
  and _40793_ (_34861_, _34860_, _34803_);
  and _40794_ (_34862_, _34861_, _34850_);
  or _40795_ (_34863_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or _40796_ (_34864_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and _40797_ (_34865_, _34864_, _34796_);
  and _40798_ (_34866_, _34865_, _34863_);
  or _40799_ (_34867_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or _40800_ (_34868_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and _40801_ (_34869_, _34868_, _34581_);
  and _40802_ (_34870_, _34869_, _34867_);
  or _40803_ (_34871_, _34870_, _34866_);
  or _40804_ (_34872_, _34871_, _34790_);
  or _40805_ (_34873_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or _40806_ (_34874_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  and _40807_ (_34875_, _34874_, _34796_);
  and _40808_ (_34876_, _34875_, _34873_);
  or _40809_ (_34877_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or _40810_ (_34878_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  and _40811_ (_34879_, _34878_, _34581_);
  and _40812_ (_34880_, _34879_, _34877_);
  or _40813_ (_34881_, _34880_, _34876_);
  or _40814_ (_34882_, _34881_, _34772_);
  and _40815_ (_34883_, _34882_, _34719_);
  and _40816_ (_34884_, _34883_, _34872_);
  or _40817_ (_34885_, _34884_, _34862_);
  or _40818_ (_34886_, _34885_, _34700_);
  and _40819_ (_34887_, _34886_, _34840_);
  and _40820_ (_34888_, _34887_, _34839_);
  and _40821_ (_34889_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and _40822_ (_34890_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or _40823_ (_34891_, _34890_, _34889_);
  and _40824_ (_34892_, _34891_, _34581_);
  and _40825_ (_34893_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and _40826_ (_34894_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or _40827_ (_34895_, _34894_, _34893_);
  and _40828_ (_34896_, _34895_, _34796_);
  or _40829_ (_34897_, _34896_, _34892_);
  and _40830_ (_34898_, _34897_, _34772_);
  and _40831_ (_34899_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and _40832_ (_34900_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or _40833_ (_34901_, _34900_, _34899_);
  and _40834_ (_34902_, _34901_, _34581_);
  and _40835_ (_34903_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and _40836_ (_34904_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or _40837_ (_34905_, _34904_, _34903_);
  and _40838_ (_34906_, _34905_, _34796_);
  or _40839_ (_34907_, _34906_, _34902_);
  and _40840_ (_34908_, _34907_, _34790_);
  or _40841_ (_34909_, _34908_, _34719_);
  or _40842_ (_34910_, _34909_, _34898_);
  or _40843_ (_34911_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or _40844_ (_34912_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and _40845_ (_34913_, _34912_, _34796_);
  and _40846_ (_34914_, _34913_, _34911_);
  or _40847_ (_34915_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or _40848_ (_34916_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and _40849_ (_34917_, _34916_, _34581_);
  and _40850_ (_34918_, _34917_, _34915_);
  or _40851_ (_34919_, _34918_, _34914_);
  and _40852_ (_34920_, _34919_, _34772_);
  or _40853_ (_34921_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or _40854_ (_34922_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and _40855_ (_34923_, _34922_, _34796_);
  and _40856_ (_34924_, _34923_, _34921_);
  or _40857_ (_34925_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or _40858_ (_34926_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and _40859_ (_34927_, _34926_, _34581_);
  and _40860_ (_34928_, _34927_, _34925_);
  or _40861_ (_34929_, _34928_, _34924_);
  and _40862_ (_34930_, _34929_, _34790_);
  or _40863_ (_34931_, _34930_, _34803_);
  or _40864_ (_34932_, _34931_, _34920_);
  and _40865_ (_34933_, _34932_, _34910_);
  or _40866_ (_34934_, _34933_, _34700_);
  and _40867_ (_34935_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and _40868_ (_34936_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or _40869_ (_34937_, _34936_, _34935_);
  and _40870_ (_34938_, _34937_, _34581_);
  and _40871_ (_34939_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and _40872_ (_34940_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or _40873_ (_34941_, _34940_, _34939_);
  and _40874_ (_34942_, _34941_, _34796_);
  or _40875_ (_34943_, _34942_, _34938_);
  and _40876_ (_34944_, _34943_, _34772_);
  and _40877_ (_34945_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  and _40878_ (_34946_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or _40879_ (_34947_, _34946_, _34945_);
  and _40880_ (_34948_, _34947_, _34581_);
  and _40881_ (_34949_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and _40882_ (_34950_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or _40883_ (_34951_, _34950_, _34949_);
  and _40884_ (_34952_, _34951_, _34796_);
  or _40885_ (_34953_, _34952_, _34948_);
  and _40886_ (_34954_, _34953_, _34790_);
  or _40887_ (_34955_, _34954_, _34719_);
  or _40888_ (_34956_, _34955_, _34944_);
  or _40889_ (_34957_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or _40890_ (_34958_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and _40891_ (_34959_, _34958_, _34957_);
  and _40892_ (_34960_, _34959_, _34581_);
  or _40893_ (_34961_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or _40894_ (_34962_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and _40895_ (_34963_, _34962_, _34961_);
  and _40896_ (_34964_, _34963_, _34796_);
  or _40897_ (_34965_, _34964_, _34960_);
  and _40898_ (_34966_, _34965_, _34772_);
  or _40899_ (_34967_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or _40900_ (_34968_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and _40901_ (_34969_, _34968_, _34967_);
  and _40902_ (_34970_, _34969_, _34581_);
  or _40903_ (_34971_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or _40904_ (_34972_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and _40905_ (_34973_, _34972_, _34971_);
  and _40906_ (_34974_, _34973_, _34796_);
  or _40907_ (_34975_, _34974_, _34970_);
  and _40908_ (_34976_, _34975_, _34790_);
  or _40909_ (_34977_, _34976_, _34803_);
  or _40910_ (_34978_, _34977_, _34966_);
  and _40911_ (_34979_, _34978_, _34956_);
  or _40912_ (_34980_, _34979_, _34789_);
  and _40913_ (_34981_, _34980_, _34638_);
  and _40914_ (_34982_, _34981_, _34934_);
  or _40915_ (_34983_, _34982_, _34888_);
  or _40916_ (_34984_, _34983_, _34692_);
  not _40917_ (_34985_, _34692_);
  and _40918_ (_34986_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  and _40919_ (_34987_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  or _40920_ (_34988_, _34987_, _34986_);
  and _40921_ (_34989_, _34988_, _34581_);
  and _40922_ (_34990_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  and _40923_ (_34991_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  or _40924_ (_34992_, _34991_, _34990_);
  and _40925_ (_34993_, _34992_, _34796_);
  or _40926_ (_34994_, _34993_, _34989_);
  and _40927_ (_34995_, _34994_, _34772_);
  and _40928_ (_34996_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  and _40929_ (_34997_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or _40930_ (_34998_, _34997_, _34996_);
  and _40931_ (_34999_, _34998_, _34581_);
  and _40932_ (_35000_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  and _40933_ (_35001_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  or _40934_ (_35002_, _35001_, _35000_);
  and _40935_ (_35003_, _35002_, _34796_);
  or _40936_ (_35004_, _35003_, _34999_);
  and _40937_ (_35005_, _35004_, _34790_);
  or _40938_ (_35006_, _35005_, _34719_);
  or _40939_ (_35007_, _35006_, _34995_);
  or _40940_ (_35008_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  or _40941_ (_35009_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  and _40942_ (_35010_, _35009_, _35008_);
  and _40943_ (_35011_, _35010_, _34581_);
  or _40944_ (_35012_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or _40945_ (_35013_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  and _40946_ (_35014_, _35013_, _35012_);
  and _40947_ (_35015_, _35014_, _34796_);
  or _40948_ (_35016_, _35015_, _35011_);
  and _40949_ (_35017_, _35016_, _34772_);
  or _40950_ (_35018_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  or _40951_ (_35019_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  and _40952_ (_35020_, _35019_, _35018_);
  and _40953_ (_35021_, _35020_, _34581_);
  or _40954_ (_35022_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  or _40955_ (_35023_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  and _40956_ (_35024_, _35023_, _35022_);
  and _40957_ (_35025_, _35024_, _34796_);
  or _40958_ (_35026_, _35025_, _35021_);
  and _40959_ (_35027_, _35026_, _34790_);
  or _40960_ (_35028_, _35027_, _34803_);
  or _40961_ (_35029_, _35028_, _35017_);
  and _40962_ (_35030_, _35029_, _35007_);
  or _40963_ (_35031_, _35030_, _34700_);
  and _40964_ (_35032_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  and _40965_ (_35033_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or _40966_ (_35034_, _35033_, _35032_);
  and _40967_ (_35035_, _35034_, _34581_);
  and _40968_ (_35036_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  and _40969_ (_35037_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or _40970_ (_35038_, _35037_, _35036_);
  and _40971_ (_35039_, _35038_, _34796_);
  or _40972_ (_35040_, _35039_, _35035_);
  and _40973_ (_35041_, _35040_, _34772_);
  and _40974_ (_35042_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and _40975_ (_35043_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or _40976_ (_35044_, _35043_, _35042_);
  and _40977_ (_35045_, _35044_, _34581_);
  and _40978_ (_35046_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and _40979_ (_35047_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or _40980_ (_35048_, _35047_, _35046_);
  and _40981_ (_35049_, _35048_, _34796_);
  or _40982_ (_35050_, _35049_, _35045_);
  and _40983_ (_35051_, _35050_, _34790_);
  or _40984_ (_35052_, _35051_, _34719_);
  or _40985_ (_35053_, _35052_, _35041_);
  or _40986_ (_35054_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or _40987_ (_35055_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and _40988_ (_35056_, _35055_, _35054_);
  and _40989_ (_35057_, _35056_, _34581_);
  or _40990_ (_35058_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or _40991_ (_35059_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and _40992_ (_35060_, _35059_, _35058_);
  and _40993_ (_35061_, _35060_, _34796_);
  or _40994_ (_35062_, _35061_, _35057_);
  and _40995_ (_35063_, _35062_, _34772_);
  or _40996_ (_35064_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or _40997_ (_35065_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and _40998_ (_35066_, _35065_, _35064_);
  and _40999_ (_35067_, _35066_, _34581_);
  or _41000_ (_35068_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or _41001_ (_35069_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  and _41002_ (_35070_, _35069_, _35068_);
  and _41003_ (_35071_, _35070_, _34796_);
  or _41004_ (_35072_, _35071_, _35067_);
  and _41005_ (_35073_, _35072_, _34790_);
  or _41006_ (_35074_, _35073_, _34803_);
  or _41007_ (_35075_, _35074_, _35063_);
  and _41008_ (_35076_, _35075_, _35053_);
  or _41009_ (_35077_, _35076_, _34789_);
  and _41010_ (_35078_, _35077_, _34638_);
  and _41011_ (_35079_, _35078_, _35031_);
  and _41012_ (_35080_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and _41013_ (_35081_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or _41014_ (_35082_, _35081_, _35080_);
  and _41015_ (_35083_, _35082_, _34796_);
  and _41016_ (_35084_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  and _41017_ (_35085_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or _41018_ (_35086_, _35085_, _35084_);
  and _41019_ (_35087_, _35086_, _34581_);
  or _41020_ (_35088_, _35087_, _35083_);
  or _41021_ (_35089_, _35088_, _34790_);
  and _41022_ (_35090_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and _41023_ (_35091_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or _41024_ (_35092_, _35091_, _35090_);
  and _41025_ (_35093_, _35092_, _34796_);
  and _41026_ (_35094_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  and _41027_ (_35095_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or _41028_ (_35096_, _35095_, _35094_);
  and _41029_ (_35097_, _35096_, _34581_);
  or _41030_ (_35098_, _35097_, _35093_);
  or _41031_ (_35099_, _35098_, _34772_);
  and _41032_ (_35100_, _35099_, _34803_);
  and _41033_ (_35101_, _35100_, _35089_);
  or _41034_ (_35102_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or _41035_ (_35103_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  and _41036_ (_35104_, _35103_, _34581_);
  and _41037_ (_35105_, _35104_, _35102_);
  or _41038_ (_35106_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or _41039_ (_35107_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and _41040_ (_35108_, _35107_, _34796_);
  and _41041_ (_35109_, _35108_, _35106_);
  or _41042_ (_35110_, _35109_, _35105_);
  or _41043_ (_35111_, _35110_, _34790_);
  or _41044_ (_35112_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or _41045_ (_35113_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  and _41046_ (_35114_, _35113_, _34581_);
  and _41047_ (_35115_, _35114_, _35112_);
  or _41048_ (_35116_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or _41049_ (_35117_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and _41050_ (_35118_, _35117_, _34796_);
  and _41051_ (_35119_, _35118_, _35116_);
  or _41052_ (_35120_, _35119_, _35115_);
  or _41053_ (_35121_, _35120_, _34772_);
  and _41054_ (_35122_, _35121_, _34719_);
  and _41055_ (_35123_, _35122_, _35111_);
  or _41056_ (_35124_, _35123_, _35101_);
  and _41057_ (_35125_, _35124_, _34789_);
  and _41058_ (_35126_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and _41059_ (_35127_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or _41060_ (_35128_, _35127_, _34581_);
  or _41061_ (_35129_, _35128_, _35126_);
  and _41062_ (_35130_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and _41063_ (_35131_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or _41064_ (_35132_, _35131_, _34796_);
  or _41065_ (_35133_, _35132_, _35130_);
  and _41066_ (_35134_, _35133_, _35129_);
  or _41067_ (_35135_, _35134_, _34790_);
  and _41068_ (_35136_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and _41069_ (_35137_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or _41070_ (_35138_, _35137_, _34581_);
  or _41071_ (_35139_, _35138_, _35136_);
  and _41072_ (_35140_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and _41073_ (_35141_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or _41074_ (_35142_, _35141_, _34796_);
  or _41075_ (_35143_, _35142_, _35140_);
  and _41076_ (_35144_, _35143_, _35139_);
  or _41077_ (_35145_, _35144_, _34772_);
  and _41078_ (_35146_, _35145_, _34803_);
  and _41079_ (_35147_, _35146_, _35135_);
  or _41080_ (_35148_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or _41081_ (_35149_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and _41082_ (_35150_, _35149_, _35148_);
  or _41083_ (_35151_, _35150_, _34796_);
  or _41084_ (_35152_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or _41085_ (_35153_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and _41086_ (_35154_, _35153_, _35152_);
  or _41087_ (_35155_, _35154_, _34581_);
  and _41088_ (_35156_, _35155_, _35151_);
  or _41089_ (_35157_, _35156_, _34790_);
  or _41090_ (_35158_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or _41091_ (_35159_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and _41092_ (_35160_, _35159_, _35158_);
  or _41093_ (_35161_, _35160_, _34796_);
  or _41094_ (_35162_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or _41095_ (_35163_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and _41096_ (_35164_, _35163_, _35162_);
  or _41097_ (_35165_, _35164_, _34581_);
  and _41098_ (_35166_, _35165_, _35161_);
  or _41099_ (_35167_, _35166_, _34772_);
  and _41100_ (_35168_, _35167_, _34719_);
  and _41101_ (_35169_, _35168_, _35157_);
  or _41102_ (_35170_, _35169_, _35147_);
  and _41103_ (_35171_, _35170_, _34700_);
  or _41104_ (_35172_, _35171_, _35125_);
  and _41105_ (_35173_, _35172_, _34840_);
  or _41106_ (_35174_, _35173_, _35079_);
  or _41107_ (_35175_, _35174_, _34985_);
  and _41108_ (_35176_, _35175_, _34984_);
  or _41109_ (_35177_, _35176_, _34346_);
  not _41110_ (_35178_, _34346_);
  and _41111_ (_35179_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and _41112_ (_35180_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or _41113_ (_35181_, _35180_, _35179_);
  and _41114_ (_35182_, _35181_, _34796_);
  and _41115_ (_35183_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and _41116_ (_35184_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or _41117_ (_35185_, _35184_, _35183_);
  and _41118_ (_35186_, _35185_, _34581_);
  or _41119_ (_35187_, _35186_, _35182_);
  or _41120_ (_35188_, _35187_, _34790_);
  and _41121_ (_35189_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and _41122_ (_35190_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or _41123_ (_35191_, _35190_, _35189_);
  and _41124_ (_35192_, _35191_, _34796_);
  and _41125_ (_35193_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and _41126_ (_35194_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or _41127_ (_35195_, _35194_, _35193_);
  and _41128_ (_35196_, _35195_, _34581_);
  or _41129_ (_35197_, _35196_, _35192_);
  or _41130_ (_35198_, _35197_, _34772_);
  and _41131_ (_35199_, _35198_, _34803_);
  and _41132_ (_35200_, _35199_, _35188_);
  or _41133_ (_35201_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or _41134_ (_35202_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and _41135_ (_35203_, _35202_, _34581_);
  and _41136_ (_35204_, _35203_, _35201_);
  or _41137_ (_35205_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or _41138_ (_35206_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and _41139_ (_35207_, _35206_, _34796_);
  and _41140_ (_35208_, _35207_, _35205_);
  or _41141_ (_35209_, _35208_, _35204_);
  or _41142_ (_35210_, _35209_, _34790_);
  or _41143_ (_35211_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or _41144_ (_35212_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and _41145_ (_35213_, _35212_, _34581_);
  and _41146_ (_35214_, _35213_, _35211_);
  or _41147_ (_35215_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or _41148_ (_35216_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and _41149_ (_35217_, _35216_, _34796_);
  and _41150_ (_35218_, _35217_, _35215_);
  or _41151_ (_35219_, _35218_, _35214_);
  or _41152_ (_35220_, _35219_, _34772_);
  and _41153_ (_35221_, _35220_, _34719_);
  and _41154_ (_35222_, _35221_, _35210_);
  or _41155_ (_35223_, _35222_, _35200_);
  and _41156_ (_35224_, _35223_, _34789_);
  and _41157_ (_35225_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and _41158_ (_35226_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or _41159_ (_35227_, _35226_, _34581_);
  or _41160_ (_35228_, _35227_, _35225_);
  and _41161_ (_35229_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and _41162_ (_35230_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or _41163_ (_35231_, _35230_, _34796_);
  or _41164_ (_35232_, _35231_, _35229_);
  and _41165_ (_35233_, _35232_, _35228_);
  or _41166_ (_35234_, _35233_, _34790_);
  and _41167_ (_35235_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and _41168_ (_35236_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or _41169_ (_35237_, _35236_, _34581_);
  or _41170_ (_35238_, _35237_, _35235_);
  and _41171_ (_35239_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and _41172_ (_35240_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or _41173_ (_35241_, _35240_, _34796_);
  or _41174_ (_35242_, _35241_, _35239_);
  and _41175_ (_35243_, _35242_, _35238_);
  or _41176_ (_35244_, _35243_, _34772_);
  and _41177_ (_35245_, _35244_, _34803_);
  and _41178_ (_35246_, _35245_, _35234_);
  or _41179_ (_35247_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or _41180_ (_35248_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and _41181_ (_35249_, _35248_, _35247_);
  or _41182_ (_35250_, _35249_, _34796_);
  or _41183_ (_35251_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or _41184_ (_35252_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and _41185_ (_35253_, _35252_, _35251_);
  or _41186_ (_35254_, _35253_, _34581_);
  and _41187_ (_35255_, _35254_, _35250_);
  or _41188_ (_35256_, _35255_, _34790_);
  or _41189_ (_35257_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or _41190_ (_35258_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and _41191_ (_35259_, _35258_, _35257_);
  or _41192_ (_35260_, _35259_, _34796_);
  or _41193_ (_35261_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or _41194_ (_35262_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and _41195_ (_35263_, _35262_, _35261_);
  or _41196_ (_35264_, _35263_, _34581_);
  and _41197_ (_35265_, _35264_, _35260_);
  or _41198_ (_35266_, _35265_, _34772_);
  and _41199_ (_35267_, _35266_, _34719_);
  and _41200_ (_35268_, _35267_, _35256_);
  or _41201_ (_35269_, _35268_, _35246_);
  and _41202_ (_35270_, _35269_, _34700_);
  or _41203_ (_35271_, _35270_, _35224_);
  and _41204_ (_35272_, _35271_, _34840_);
  and _41205_ (_35273_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  and _41206_ (_35274_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  or _41207_ (_35275_, _35274_, _35273_);
  and _41208_ (_35276_, _35275_, _34581_);
  and _41209_ (_35277_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  and _41210_ (_35278_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  or _41211_ (_35279_, _35278_, _35277_);
  and _41212_ (_35280_, _35279_, _34796_);
  or _41213_ (_35281_, _35280_, _35276_);
  and _41214_ (_35282_, _35281_, _34772_);
  and _41215_ (_35283_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  and _41216_ (_35284_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  or _41217_ (_35285_, _35284_, _35283_);
  and _41218_ (_35286_, _35285_, _34581_);
  and _41219_ (_35287_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  and _41220_ (_35288_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  or _41221_ (_35289_, _35288_, _35287_);
  and _41222_ (_35290_, _35289_, _34796_);
  or _41223_ (_35291_, _35290_, _35286_);
  and _41224_ (_35292_, _35291_, _34790_);
  or _41225_ (_35293_, _35292_, _35282_);
  and _41226_ (_35294_, _35293_, _34803_);
  or _41227_ (_35295_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  or _41228_ (_35296_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  and _41229_ (_35297_, _35296_, _35295_);
  and _41230_ (_35298_, _35297_, _34581_);
  or _41231_ (_35299_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  or _41232_ (_35300_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  and _41233_ (_35301_, _35300_, _35299_);
  and _41234_ (_35302_, _35301_, _34796_);
  or _41235_ (_35303_, _35302_, _35298_);
  and _41236_ (_35304_, _35303_, _34772_);
  or _41237_ (_35305_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  or _41238_ (_35306_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  and _41239_ (_35307_, _35306_, _35305_);
  and _41240_ (_35308_, _35307_, _34581_);
  or _41241_ (_35309_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  or _41242_ (_35310_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  and _41243_ (_35311_, _35310_, _35309_);
  and _41244_ (_35312_, _35311_, _34796_);
  or _41245_ (_35313_, _35312_, _35308_);
  and _41246_ (_35314_, _35313_, _34790_);
  or _41247_ (_35315_, _35314_, _35304_);
  and _41248_ (_35316_, _35315_, _34719_);
  or _41249_ (_35317_, _35316_, _35294_);
  and _41250_ (_35318_, _35317_, _34789_);
  and _41251_ (_35319_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and _41252_ (_35320_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or _41253_ (_35321_, _35320_, _35319_);
  and _41254_ (_35322_, _35321_, _34581_);
  and _41255_ (_35323_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and _41256_ (_35324_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or _41257_ (_35325_, _35324_, _35323_);
  and _41258_ (_35326_, _35325_, _34796_);
  or _41259_ (_35327_, _35326_, _35322_);
  and _41260_ (_35328_, _35327_, _34772_);
  and _41261_ (_35329_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and _41262_ (_35330_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or _41263_ (_35331_, _35330_, _35329_);
  and _41264_ (_35332_, _35331_, _34581_);
  and _41265_ (_35333_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and _41266_ (_35334_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or _41267_ (_35335_, _35334_, _35333_);
  and _41268_ (_35336_, _35335_, _34796_);
  or _41269_ (_35337_, _35336_, _35332_);
  and _41270_ (_35338_, _35337_, _34790_);
  or _41271_ (_35339_, _35338_, _35328_);
  and _41272_ (_35340_, _35339_, _34803_);
  or _41273_ (_35341_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or _41274_ (_35342_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and _41275_ (_35343_, _35342_, _35341_);
  and _41276_ (_35344_, _35343_, _34581_);
  or _41277_ (_35345_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or _41278_ (_35346_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and _41279_ (_35347_, _35346_, _35345_);
  and _41280_ (_35348_, _35347_, _34796_);
  or _41281_ (_35349_, _35348_, _35344_);
  and _41282_ (_35350_, _35349_, _34772_);
  or _41283_ (_35351_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or _41284_ (_35352_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and _41285_ (_35353_, _35352_, _35351_);
  and _41286_ (_35354_, _35353_, _34581_);
  or _41287_ (_35355_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or _41288_ (_35356_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and _41289_ (_35357_, _35356_, _35355_);
  and _41290_ (_35358_, _35357_, _34796_);
  or _41291_ (_35359_, _35358_, _35354_);
  and _41292_ (_35360_, _35359_, _34790_);
  or _41293_ (_35361_, _35360_, _35350_);
  and _41294_ (_35362_, _35361_, _34719_);
  or _41295_ (_35363_, _35362_, _35340_);
  and _41296_ (_35364_, _35363_, _34700_);
  or _41297_ (_35365_, _35364_, _35318_);
  and _41298_ (_35366_, _35365_, _34638_);
  or _41299_ (_35367_, _35366_, _35272_);
  or _41300_ (_35368_, _35367_, _34692_);
  and _41301_ (_35369_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and _41302_ (_35370_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or _41303_ (_35371_, _35370_, _35369_);
  and _41304_ (_35372_, _35371_, _34581_);
  and _41305_ (_35373_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and _41306_ (_35374_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or _41307_ (_35375_, _35374_, _35373_);
  and _41308_ (_35376_, _35375_, _34796_);
  or _41309_ (_35377_, _35376_, _35372_);
  or _41310_ (_35378_, _35377_, _34790_);
  and _41311_ (_35379_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and _41312_ (_35380_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or _41313_ (_35381_, _35380_, _35379_);
  and _41314_ (_35382_, _35381_, _34581_);
  and _41315_ (_35383_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and _41316_ (_35384_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or _41317_ (_35385_, _35384_, _35383_);
  and _41318_ (_35386_, _35385_, _34796_);
  or _41319_ (_35387_, _35386_, _35382_);
  or _41320_ (_35388_, _35387_, _34772_);
  and _41321_ (_35389_, _35388_, _34803_);
  and _41322_ (_35390_, _35389_, _35378_);
  or _41323_ (_35391_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or _41324_ (_35392_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and _41325_ (_35393_, _35392_, _34796_);
  and _41326_ (_35394_, _35393_, _35391_);
  or _41327_ (_35395_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or _41328_ (_35396_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and _41329_ (_35397_, _35396_, _34581_);
  and _41330_ (_35398_, _35397_, _35395_);
  or _41331_ (_35399_, _35398_, _35394_);
  or _41332_ (_35400_, _35399_, _34790_);
  or _41333_ (_35401_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or _41334_ (_35402_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and _41335_ (_35403_, _35402_, _34796_);
  and _41336_ (_35404_, _35403_, _35401_);
  or _41337_ (_35405_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or _41338_ (_35406_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and _41339_ (_35407_, _35406_, _34581_);
  and _41340_ (_35408_, _35407_, _35405_);
  or _41341_ (_35409_, _35408_, _35404_);
  or _41342_ (_35410_, _35409_, _34772_);
  and _41343_ (_35411_, _35410_, _34719_);
  and _41344_ (_35412_, _35411_, _35400_);
  or _41345_ (_35413_, _35412_, _35390_);
  and _41346_ (_35414_, _35413_, _34789_);
  and _41347_ (_35415_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and _41348_ (_35416_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or _41349_ (_35417_, _35416_, _35415_);
  and _41350_ (_35418_, _35417_, _34581_);
  and _41351_ (_35419_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and _41352_ (_35420_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or _41353_ (_35421_, _35420_, _35419_);
  and _41354_ (_35422_, _35421_, _34796_);
  or _41355_ (_35423_, _35422_, _35418_);
  or _41356_ (_35424_, _35423_, _34790_);
  and _41357_ (_35425_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and _41358_ (_35426_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or _41359_ (_35427_, _35426_, _35425_);
  and _41360_ (_35428_, _35427_, _34581_);
  and _41361_ (_35429_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and _41362_ (_35430_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or _41363_ (_35431_, _35430_, _35429_);
  and _41364_ (_35432_, _35431_, _34796_);
  or _41365_ (_35433_, _35432_, _35428_);
  or _41366_ (_35434_, _35433_, _34772_);
  and _41367_ (_35435_, _35434_, _34803_);
  and _41368_ (_35436_, _35435_, _35424_);
  or _41369_ (_35437_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or _41370_ (_35438_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and _41371_ (_35439_, _35438_, _35437_);
  and _41372_ (_35440_, _35439_, _34581_);
  or _41373_ (_35441_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or _41374_ (_35442_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and _41375_ (_35443_, _35442_, _35441_);
  and _41376_ (_35444_, _35443_, _34796_);
  or _41377_ (_35445_, _35444_, _35440_);
  or _41378_ (_35446_, _35445_, _34790_);
  or _41379_ (_35447_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or _41380_ (_35448_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and _41381_ (_35449_, _35448_, _35447_);
  and _41382_ (_35450_, _35449_, _34581_);
  or _41383_ (_35451_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or _41384_ (_35452_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and _41385_ (_35453_, _35452_, _35451_);
  and _41386_ (_35454_, _35453_, _34796_);
  or _41387_ (_35455_, _35454_, _35450_);
  or _41388_ (_35456_, _35455_, _34772_);
  and _41389_ (_35457_, _35456_, _34719_);
  and _41390_ (_35458_, _35457_, _35446_);
  or _41391_ (_35459_, _35458_, _35436_);
  and _41392_ (_35460_, _35459_, _34700_);
  or _41393_ (_35461_, _35460_, _35414_);
  and _41394_ (_35462_, _35461_, _34840_);
  or _41395_ (_35463_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or _41396_ (_35464_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and _41397_ (_35465_, _35464_, _35463_);
  and _41398_ (_35466_, _35465_, _34581_);
  or _41399_ (_35467_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or _41400_ (_35468_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and _41401_ (_35469_, _35468_, _35467_);
  and _41402_ (_35470_, _35469_, _34796_);
  or _41403_ (_35471_, _35470_, _35466_);
  and _41404_ (_35472_, _35471_, _34790_);
  or _41405_ (_35473_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or _41406_ (_35474_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and _41407_ (_35475_, _35474_, _35473_);
  and _41408_ (_35476_, _35475_, _34581_);
  or _41409_ (_35477_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or _41410_ (_35478_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and _41411_ (_35479_, _35478_, _35477_);
  and _41412_ (_35480_, _35479_, _34796_);
  or _41413_ (_35481_, _35480_, _35476_);
  and _41414_ (_35482_, _35481_, _34772_);
  or _41415_ (_35483_, _35482_, _35472_);
  and _41416_ (_35484_, _35483_, _34719_);
  and _41417_ (_35485_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and _41418_ (_35486_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or _41419_ (_35487_, _35486_, _35485_);
  and _41420_ (_35488_, _35487_, _34581_);
  and _41421_ (_35489_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and _41422_ (_35490_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or _41423_ (_35491_, _35490_, _35489_);
  and _41424_ (_35492_, _35491_, _34796_);
  or _41425_ (_35493_, _35492_, _35488_);
  and _41426_ (_35494_, _35493_, _34790_);
  and _41427_ (_35495_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and _41428_ (_35496_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or _41429_ (_35497_, _35496_, _35495_);
  and _41430_ (_35498_, _35497_, _34581_);
  and _41431_ (_35499_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and _41432_ (_35500_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or _41433_ (_35501_, _35500_, _35499_);
  and _41434_ (_35502_, _35501_, _34796_);
  or _41435_ (_35503_, _35502_, _35498_);
  and _41436_ (_35504_, _35503_, _34772_);
  or _41437_ (_35505_, _35504_, _35494_);
  and _41438_ (_35506_, _35505_, _34803_);
  or _41439_ (_35507_, _35506_, _35484_);
  and _41440_ (_35508_, _35507_, _34700_);
  or _41441_ (_35509_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or _41442_ (_35510_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  and _41443_ (_35511_, _35510_, _34796_);
  and _41444_ (_35512_, _35511_, _35509_);
  or _41445_ (_35513_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or _41446_ (_35514_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and _41447_ (_35515_, _35514_, _34581_);
  and _41448_ (_35516_, _35515_, _35513_);
  or _41449_ (_35517_, _35516_, _35512_);
  and _41450_ (_35518_, _35517_, _34790_);
  or _41451_ (_35519_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or _41452_ (_35520_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and _41453_ (_35521_, _35520_, _34796_);
  and _41454_ (_35522_, _35521_, _35519_);
  or _41455_ (_35523_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or _41456_ (_35524_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  and _41457_ (_35525_, _35524_, _34581_);
  and _41458_ (_35526_, _35525_, _35523_);
  or _41459_ (_35527_, _35526_, _35522_);
  and _41460_ (_35528_, _35527_, _34772_);
  or _41461_ (_35529_, _35528_, _35518_);
  and _41462_ (_35530_, _35529_, _34719_);
  and _41463_ (_35531_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and _41464_ (_35532_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or _41465_ (_35533_, _35532_, _35531_);
  and _41466_ (_35534_, _35533_, _34581_);
  and _41467_ (_35535_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and _41468_ (_35536_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or _41469_ (_35537_, _35536_, _35535_);
  and _41470_ (_35538_, _35537_, _34796_);
  or _41471_ (_35539_, _35538_, _35534_);
  and _41472_ (_35540_, _35539_, _34790_);
  and _41473_ (_35541_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and _41474_ (_35542_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or _41475_ (_35543_, _35542_, _35541_);
  and _41476_ (_35544_, _35543_, _34581_);
  and _41477_ (_35545_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and _41478_ (_35546_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or _41479_ (_35547_, _35546_, _35545_);
  and _41480_ (_35548_, _35547_, _34796_);
  or _41481_ (_35549_, _35548_, _35544_);
  and _41482_ (_35550_, _35549_, _34772_);
  or _41483_ (_35551_, _35550_, _35540_);
  and _41484_ (_35552_, _35551_, _34803_);
  or _41485_ (_35553_, _35552_, _35530_);
  and _41486_ (_35554_, _35553_, _34789_);
  or _41487_ (_35555_, _35554_, _35508_);
  and _41488_ (_35556_, _35555_, _34638_);
  or _41489_ (_35557_, _35556_, _35462_);
  or _41490_ (_35558_, _35557_, _34985_);
  and _41491_ (_35559_, _35558_, _35368_);
  or _41492_ (_35560_, _35559_, _35178_);
  and _41493_ (_35561_, _35560_, _35177_);
  or _41494_ (_35562_, _35561_, _34788_);
  not _41495_ (_38997_, rst);
  not _41496_ (_35563_, _34788_);
  or _41497_ (_35564_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and _41498_ (_35565_, _35564_, _38997_);
  and _41499_ (_38984_[7], _35565_, _35562_);
  nor _41500_ (_35566_, _34785_, _34477_);
  nor _41501_ (_35567_, _34785_, _34584_);
  nor _41502_ (_35568_, _35567_, _35566_);
  nor _41503_ (_35569_, _34785_, _34775_);
  nor _41504_ (_35570_, _34785_, _34716_);
  nor _41505_ (_35571_, _35570_, _35569_);
  and _41506_ (_35572_, _35571_, _35568_);
  and _41507_ (_35573_, _34784_, _34701_);
  and _41508_ (_35574_, _34784_, _34640_);
  nor _41509_ (_35575_, _35574_, _35573_);
  nor _41510_ (_35576_, _34474_, _34249_);
  and _41511_ (_35577_, _35576_, _34784_);
  not _41512_ (_35578_, _35577_);
  and _41513_ (_35579_, _35578_, _35575_);
  and _41514_ (_35580_, _35579_, _34784_);
  and _41515_ (_35581_, _35580_, _35572_);
  and _41516_ (_35582_, _33930_, _33898_);
  not _41517_ (_35583_, _35582_);
  and _41518_ (_35584_, _34197_, _34180_);
  not _41519_ (_35585_, _33778_);
  nor _41520_ (_35586_, _35585_, _33765_);
  not _41521_ (_35587_, _33951_);
  nor _41522_ (_35588_, _35587_, _33797_);
  and _41523_ (_35589_, _34007_, _33883_);
  nor _41524_ (_35590_, _35589_, _33967_);
  nor _41525_ (_35591_, _35590_, _35588_);
  nor _41526_ (_35592_, _35591_, _33916_);
  nor _41527_ (_35593_, _35592_, _35586_);
  and _41528_ (_35594_, _35591_, _33916_);
  nor _41529_ (_35595_, _35594_, _35592_);
  not _41530_ (_35596_, _35595_);
  and _41531_ (_35597_, _35589_, _33967_);
  nor _41532_ (_35598_, _35597_, _35590_);
  not _41533_ (_35599_, _35598_);
  not _41534_ (_35600_, _33991_);
  and _41535_ (_35601_, _34061_, _34057_);
  and _41536_ (_35602_, _35601_, _33865_);
  nor _41537_ (_35603_, _34098_, _33831_);
  and _41538_ (_35604_, _34131_, _33848_);
  nor _41539_ (_35605_, _35604_, _34111_);
  nor _41540_ (_35606_, _35605_, _35603_);
  nor _41541_ (_35607_, _35606_, _34077_);
  nor _41542_ (_35608_, _35607_, _35602_);
  nor _41543_ (_35609_, _35608_, _34040_);
  and _41544_ (_35610_, _35608_, _34040_);
  nor _41545_ (_35611_, _35610_, _35609_);
  not _41546_ (_35612_, _35611_);
  and _41547_ (_35613_, _35606_, _34077_);
  nor _41548_ (_35614_, _35613_, _35607_);
  not _41549_ (_35615_, _35614_);
  and _41550_ (_35616_, _35604_, _34111_);
  nor _41551_ (_35617_, _35616_, _35605_);
  not _41552_ (_35618_, _35617_);
  nor _41553_ (_35619_, _34135_, _33734_);
  and _41554_ (_35620_, _35619_, _35618_);
  and _41555_ (_35621_, _35620_, _35615_);
  and _41556_ (_35622_, _35621_, _35612_);
  not _41557_ (_35623_, _34035_);
  or _41558_ (_35624_, _35623_, _33814_);
  and _41559_ (_35625_, _35623_, _33814_);
  or _41560_ (_35626_, _35608_, _35625_);
  and _41561_ (_35627_, _35626_, _35624_);
  or _41562_ (_35628_, _35627_, _35622_);
  and _41563_ (_35629_, _35628_, _35600_);
  and _41564_ (_35630_, _35629_, _35599_);
  and _41565_ (_35631_, _35630_, _35596_);
  nor _41566_ (_35632_, _35631_, _35593_);
  nor _41567_ (_35633_, _35632_, _34207_);
  nor _41568_ (_35634_, _35633_, _35584_);
  nor _41569_ (_35635_, _35634_, _35583_);
  not _41570_ (_35636_, _35635_);
  and _41571_ (_35637_, _33930_, _33906_);
  not _41572_ (_35638_, _35637_);
  not _41573_ (_35639_, _34207_);
  not _41574_ (_35640_, _34077_);
  and _41575_ (_35641_, _34134_, _34111_);
  nor _41576_ (_35642_, _35641_, _34110_);
  nor _41577_ (_35643_, _35642_, _35640_);
  nor _41578_ (_35644_, _35643_, _34076_);
  nor _41579_ (_35645_, _35644_, _34040_);
  and _41580_ (_35646_, _35644_, _34040_);
  nor _41581_ (_35647_, _35646_, _35645_);
  not _41582_ (_35648_, _34135_);
  nor _41583_ (_35649_, _35648_, _33734_);
  and _41584_ (_35650_, _35649_, _34111_);
  and _41585_ (_35651_, _35642_, _35640_);
  nor _41586_ (_35652_, _35651_, _35643_);
  and _41587_ (_35653_, _35652_, _35650_);
  not _41588_ (_35654_, _35653_);
  nor _41589_ (_35655_, _35654_, _35647_);
  nor _41590_ (_35656_, _35644_, _34036_);
  or _41591_ (_35657_, _35656_, _34038_);
  or _41592_ (_35658_, _35657_, _35655_);
  and _41593_ (_35659_, _35658_, _33991_);
  and _41594_ (_35660_, _35659_, _33967_);
  not _41595_ (_35661_, _33916_);
  and _41596_ (_35662_, _33990_, _33967_);
  nor _41597_ (_35663_, _35662_, _33966_);
  nor _41598_ (_35664_, _35663_, _35661_);
  and _41599_ (_35665_, _35663_, _35661_);
  nor _41600_ (_35666_, _35665_, _35664_);
  and _41601_ (_35667_, _35666_, _35660_);
  not _41602_ (_35668_, _35667_);
  nor _41603_ (_35669_, _35664_, _33915_);
  and _41604_ (_35670_, _35669_, _35668_);
  nor _41605_ (_35671_, _35670_, _35639_);
  nor _41606_ (_35672_, _35671_, _34206_);
  nor _41607_ (_35673_, _35672_, _35638_);
  and _41608_ (_35674_, _33730_, _33728_);
  and _41609_ (_35675_, _33908_, _33898_);
  and _41610_ (_35676_, _33922_, _33728_);
  nor _41611_ (_35677_, _35676_, _35675_);
  nor _41612_ (_35678_, _35677_, _35674_);
  nor _41613_ (_35679_, _33924_, _33888_);
  not _41614_ (_35680_, _33733_);
  and _41615_ (_35681_, _33913_, _33671_);
  nor _41616_ (_35682_, _35681_, _35680_);
  nor _41617_ (_35683_, _35682_, _33732_);
  not _41618_ (_35684_, _35683_);
  nor _41619_ (_35685_, _35684_, _35679_);
  nor _41620_ (_35686_, _35685_, _35678_);
  not _41621_ (_35687_, _34183_);
  and _41622_ (_35688_, _33921_, _33906_);
  and _41623_ (_35689_, _34064_, _33831_);
  nor _41624_ (_35690_, _35689_, _33814_);
  and _41625_ (_35691_, _35690_, _35688_);
  and _41626_ (_35692_, _35691_, _33884_);
  nor _41627_ (_35693_, _35692_, _35687_);
  and _41628_ (_35694_, _35693_, _33734_);
  nor _41629_ (_35695_, _35694_, _34200_);
  not _41630_ (_35696_, _35688_);
  nor _41631_ (_35697_, _33734_, _34180_);
  not _41632_ (_35698_, _35697_);
  nor _41633_ (_35699_, _35698_, _35693_);
  nor _41634_ (_35700_, _35699_, _35696_);
  and _41635_ (_35701_, _35700_, _35695_);
  nor _41636_ (_35702_, _33733_, _33728_);
  not _41637_ (_35703_, _33914_);
  nor _41638_ (_35704_, _35703_, _33732_);
  nor _41639_ (_35705_, _35704_, _33909_);
  nor _41640_ (_35706_, _35705_, _35702_);
  not _41641_ (_35707_, _34180_);
  and _41642_ (_35708_, _33908_, _33673_);
  and _41643_ (_35709_, _35708_, _35707_);
  and _41644_ (_35710_, _33935_, _33888_);
  not _41645_ (_35711_, _33848_);
  and _41646_ (_35712_, _33906_, _33671_);
  and _41647_ (_35713_, _35712_, _35711_);
  or _41648_ (_35714_, _35691_, _35713_);
  or _41649_ (_35715_, _35714_, _35710_);
  or _41650_ (_35716_, _35715_, _35709_);
  or _41651_ (_35717_, _35716_, _35706_);
  nor _41652_ (_35718_, _35717_, _35701_);
  and _41653_ (_35719_, _35718_, _35686_);
  not _41654_ (_35720_, _35719_);
  nor _41655_ (_35721_, _35720_, _35673_);
  and _41656_ (_35722_, _35721_, _35636_);
  not _41657_ (_35723_, _35722_);
  and _41658_ (_35724_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _33705_);
  and _41659_ (_35725_, _35724_, _33695_);
  and _41660_ (_35726_, _35725_, _35723_);
  nor _41661_ (_35727_, _34148_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  not _41662_ (_35728_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _41663_ (_35729_, _35725_, _35728_);
  and _41664_ (_35730_, _35729_, _33717_);
  or _41665_ (_35731_, _35730_, _35727_);
  or _41666_ (_35732_, _35731_, _35726_);
  and _41667_ (_35733_, _35732_, _35581_);
  not _41668_ (_35734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor _41669_ (_35735_, _35581_, _35734_);
  or _41670_ (_36928_, _35735_, _35733_);
  not _41671_ (_35736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _41672_ (_35737_, _35581_, _35736_);
  nand _41673_ (_35738_, _35724_, _33690_);
  nor _41674_ (_35739_, _35738_, _35722_);
  and _41675_ (_35740_, _34122_, _35728_);
  and _41676_ (_35741_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _41677_ (_35742_, _35724_, _33700_);
  or _41678_ (_35743_, _35742_, _35741_);
  and _41679_ (_35744_, _35724_, _33683_);
  or _41680_ (_35745_, _35744_, _35743_);
  and _41681_ (_35746_, _35745_, _33721_);
  or _41682_ (_35747_, _35746_, _35740_);
  or _41683_ (_35748_, _35747_, _35739_);
  and _41684_ (_35749_, _35748_, _35581_);
  or _41685_ (_36929_, _35749_, _35737_);
  nand _41686_ (_35750_, _35724_, _33684_);
  nor _41687_ (_35751_, _35750_, _35722_);
  and _41688_ (_35752_, _34089_, _35728_);
  nand _41689_ (_35753_, _33684_, _33705_);
  and _41690_ (_35754_, _33708_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _41691_ (_35755_, _35754_, _35753_);
  or _41692_ (_35756_, _35755_, _35752_);
  or _41693_ (_35757_, _35756_, _35751_);
  and _41694_ (_35758_, _35757_, _35581_);
  not _41695_ (_35759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor _41696_ (_35760_, _35581_, _35759_);
  or _41697_ (_36930_, _35760_, _35758_);
  and _41698_ (_35761_, _35742_, _35723_);
  nor _41699_ (_35762_, _34052_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _41700_ (_35763_, _33700_, _33705_);
  and _41701_ (_35764_, _33713_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _41702_ (_35765_, _35764_, _35763_);
  or _41703_ (_35766_, _35765_, _35762_);
  or _41704_ (_35767_, _35766_, _35761_);
  and _41705_ (_35768_, _35767_, _35581_);
  not _41706_ (_35769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor _41707_ (_35770_, _35581_, _35769_);
  or _41708_ (_36931_, _35770_, _35768_);
  nand _41709_ (_35771_, _35741_, _33695_);
  nor _41710_ (_35772_, _35771_, _35722_);
  nor _41711_ (_35773_, _34017_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _41712_ (_35774_, _33695_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _41713_ (_35775_, _33694_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _41714_ (_35776_, _35775_, _35774_);
  or _41715_ (_35777_, _35776_, _35773_);
  or _41716_ (_35778_, _35777_, _35772_);
  and _41717_ (_35779_, _35778_, _35581_);
  not _41718_ (_35780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _41719_ (_35781_, _35581_, _35780_);
  or _41720_ (_36932_, _35781_, _35779_);
  not _41721_ (_35782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _41722_ (_35783_, _35581_, _35782_);
  nand _41723_ (_35784_, _35741_, _33690_);
  nor _41724_ (_35785_, _35784_, _35722_);
  and _41725_ (_35786_, _33978_, _35728_);
  nand _41726_ (_35787_, _33690_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _41727_ (_35788_, _33689_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _41728_ (_35789_, _35788_, _35787_);
  or _41729_ (_35790_, _35789_, _35786_);
  or _41730_ (_35791_, _35790_, _35785_);
  and _41731_ (_35792_, _35791_, _35581_);
  or _41732_ (_36933_, _35792_, _35783_);
  not _41733_ (_35793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _41734_ (_35794_, _35581_, _35793_);
  nand _41735_ (_35795_, _35741_, _33684_);
  nor _41736_ (_35796_, _35795_, _35722_);
  and _41737_ (_35797_, _33942_, _35728_);
  nand _41738_ (_35798_, _33684_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _41739_ (_35799_, _33682_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _41740_ (_35800_, _35799_, _35798_);
  or _41741_ (_35801_, _35800_, _35797_);
  or _41742_ (_35802_, _35801_, _35796_);
  and _41743_ (_35803_, _35802_, _35581_);
  or _41744_ (_36934_, _35803_, _35794_);
  not _41745_ (_35804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor _41746_ (_35805_, _35581_, _35804_);
  and _41747_ (_35806_, _35741_, _33700_);
  not _41748_ (_35807_, _35806_);
  nor _41749_ (_35808_, _35807_, _35722_);
  nand _41750_ (_35809_, _34221_, _35728_);
  or _41751_ (_35810_, _33699_, _35728_);
  and _41752_ (_35811_, _35810_, _35807_);
  and _41753_ (_35812_, _35811_, _35809_);
  or _41754_ (_35813_, _35812_, _35808_);
  and _41755_ (_35814_, _35813_, _35581_);
  or _41756_ (_36935_, _35814_, _35805_);
  and _41757_ (_35815_, _35732_, _34784_);
  and _41758_ (_35816_, _35566_, _34584_);
  and _41759_ (_35817_, _35816_, _35571_);
  and _41760_ (_35818_, _35817_, _35579_);
  and _41761_ (_35819_, _35818_, _35815_);
  not _41762_ (_35820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor _41763_ (_35821_, _35818_, _35820_);
  or _41764_ (_37816_, _35821_, _35819_);
  and _41765_ (_35822_, _35748_, _34784_);
  and _41766_ (_35823_, _35818_, _35822_);
  not _41767_ (_35824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor _41768_ (_35825_, _35818_, _35824_);
  or _41769_ (_37817_, _35825_, _35823_);
  and _41770_ (_35826_, _35757_, _34784_);
  and _41771_ (_35827_, _35818_, _35826_);
  not _41772_ (_35828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor _41773_ (_35829_, _35818_, _35828_);
  or _41774_ (_37818_, _35829_, _35827_);
  and _41775_ (_35830_, _35767_, _34784_);
  and _41776_ (_35831_, _35818_, _35830_);
  not _41777_ (_35832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor _41778_ (_35833_, _35818_, _35832_);
  or _41779_ (_37819_, _35833_, _35831_);
  and _41780_ (_35834_, _35778_, _34784_);
  and _41781_ (_35835_, _35818_, _35834_);
  not _41782_ (_35836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor _41783_ (_35837_, _35818_, _35836_);
  or _41784_ (_37820_, _35837_, _35835_);
  and _41785_ (_35838_, _35791_, _34784_);
  and _41786_ (_35839_, _35818_, _35838_);
  not _41787_ (_35840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor _41788_ (_35841_, _35818_, _35840_);
  or _41789_ (_37821_, _35841_, _35839_);
  and _41790_ (_35842_, _35802_, _34784_);
  and _41791_ (_35843_, _35818_, _35842_);
  not _41792_ (_35844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor _41793_ (_35845_, _35818_, _35844_);
  or _41794_ (_37822_, _35845_, _35843_);
  and _41795_ (_35846_, _35813_, _34784_);
  and _41796_ (_35847_, _35818_, _35846_);
  not _41797_ (_35848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor _41798_ (_35849_, _35818_, _35848_);
  or _41799_ (_37823_, _35849_, _35847_);
  and _41800_ (_35850_, _35567_, _34477_);
  and _41801_ (_35851_, _35850_, _35571_);
  and _41802_ (_35852_, _35851_, _35579_);
  and _41803_ (_35853_, _35852_, _35815_);
  not _41804_ (_35854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor _41805_ (_35855_, _35852_, _35854_);
  or _41806_ (_38360_, _35855_, _35853_);
  and _41807_ (_35856_, _35852_, _35822_);
  not _41808_ (_35857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor _41809_ (_35858_, _35852_, _35857_);
  or _41810_ (_38361_, _35858_, _35856_);
  and _41811_ (_35859_, _35852_, _35826_);
  not _41812_ (_35860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor _41813_ (_35861_, _35852_, _35860_);
  or _41814_ (_38362_, _35861_, _35859_);
  and _41815_ (_35862_, _35852_, _35830_);
  not _41816_ (_35863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor _41817_ (_35864_, _35852_, _35863_);
  or _41818_ (_38363_, _35864_, _35862_);
  and _41819_ (_35865_, _35852_, _35834_);
  not _41820_ (_35866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor _41821_ (_35867_, _35852_, _35866_);
  or _41822_ (_38364_, _35867_, _35865_);
  and _41823_ (_35868_, _35852_, _35838_);
  not _41824_ (_35869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor _41825_ (_35870_, _35852_, _35869_);
  or _41826_ (_38365_, _35870_, _35868_);
  and _41827_ (_35871_, _35852_, _35842_);
  not _41828_ (_35872_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor _41829_ (_35873_, _35852_, _35872_);
  or _41830_ (_38366_, _35873_, _35871_);
  and _41831_ (_35874_, _35852_, _35846_);
  not _41832_ (_35875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor _41833_ (_35876_, _35852_, _35875_);
  or _41834_ (_38367_, _35876_, _35874_);
  and _41835_ (_35877_, _35567_, _35566_);
  and _41836_ (_35878_, _35877_, _35571_);
  and _41837_ (_35879_, _35878_, _35579_);
  and _41838_ (_35880_, _35879_, _35815_);
  not _41839_ (_35881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor _41840_ (_35882_, _35879_, _35881_);
  or _41841_ (_38448_, _35882_, _35880_);
  and _41842_ (_35883_, _35879_, _35822_);
  not _41843_ (_35884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor _41844_ (_35885_, _35879_, _35884_);
  or _41845_ (_38449_, _35885_, _35883_);
  and _41846_ (_35886_, _35879_, _35826_);
  not _41847_ (_35887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor _41848_ (_35888_, _35879_, _35887_);
  or _41849_ (_38450_, _35888_, _35886_);
  and _41850_ (_35889_, _35879_, _35830_);
  not _41851_ (_35890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor _41852_ (_35891_, _35879_, _35890_);
  or _41853_ (_38451_, _35891_, _35889_);
  and _41854_ (_35892_, _35879_, _35834_);
  not _41855_ (_35893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor _41856_ (_35894_, _35879_, _35893_);
  or _41857_ (_38452_, _35894_, _35892_);
  and _41858_ (_35895_, _35879_, _35838_);
  not _41859_ (_35896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor _41860_ (_35897_, _35879_, _35896_);
  or _41861_ (_38453_, _35897_, _35895_);
  and _41862_ (_35898_, _35879_, _35842_);
  not _41863_ (_35899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor _41864_ (_35900_, _35879_, _35899_);
  or _41865_ (_38454_, _35900_, _35898_);
  and _41866_ (_35901_, _35879_, _35846_);
  not _41867_ (_35902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor _41868_ (_35903_, _35879_, _35902_);
  or _41869_ (_38455_, _35903_, _35901_);
  and _41870_ (_35904_, _35569_, _34716_);
  and _41871_ (_35905_, _35904_, _35568_);
  and _41872_ (_35906_, _35905_, _35579_);
  and _41873_ (_35907_, _35906_, _35815_);
  not _41874_ (_35908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor _41875_ (_35909_, _35906_, _35908_);
  or _41876_ (_38536_, _35909_, _35907_);
  and _41877_ (_35910_, _35906_, _35822_);
  not _41878_ (_35911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor _41879_ (_35912_, _35906_, _35911_);
  or _41880_ (_38537_, _35912_, _35910_);
  and _41881_ (_35913_, _35906_, _35826_);
  not _41882_ (_35914_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor _41883_ (_35915_, _35906_, _35914_);
  or _41884_ (_38538_, _35915_, _35913_);
  and _41885_ (_35916_, _35906_, _35830_);
  not _41886_ (_35917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor _41887_ (_35918_, _35906_, _35917_);
  or _41888_ (_38539_, _35918_, _35916_);
  and _41889_ (_35919_, _35906_, _35834_);
  not _41890_ (_35920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor _41891_ (_35921_, _35906_, _35920_);
  or _41892_ (_38540_, _35921_, _35919_);
  and _41893_ (_35922_, _35906_, _35838_);
  not _41894_ (_35923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor _41895_ (_35924_, _35906_, _35923_);
  or _41896_ (_38541_, _35924_, _35922_);
  and _41897_ (_35925_, _35906_, _35842_);
  not _41898_ (_35926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor _41899_ (_35927_, _35906_, _35926_);
  or _41900_ (_38542_, _35927_, _35925_);
  and _41901_ (_35928_, _35906_, _35846_);
  not _41902_ (_35929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor _41903_ (_35930_, _35906_, _35929_);
  or _41904_ (_38543_, _35930_, _35928_);
  and _41905_ (_35931_, _35904_, _35816_);
  and _41906_ (_35932_, _35931_, _35579_);
  and _41907_ (_35933_, _35932_, _35815_);
  not _41908_ (_35934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor _41909_ (_35935_, _35932_, _35934_);
  or _41910_ (_38624_, _35935_, _35933_);
  and _41911_ (_35936_, _35932_, _35822_);
  not _41912_ (_35937_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor _41913_ (_35938_, _35932_, _35937_);
  or _41914_ (_38625_, _35938_, _35936_);
  and _41915_ (_35939_, _35932_, _35826_);
  not _41916_ (_35940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor _41917_ (_35941_, _35932_, _35940_);
  or _41918_ (_38626_, _35941_, _35939_);
  and _41919_ (_35942_, _35932_, _35830_);
  not _41920_ (_35943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor _41921_ (_35944_, _35932_, _35943_);
  or _41922_ (_38627_, _35944_, _35942_);
  and _41923_ (_35945_, _35932_, _35834_);
  not _41924_ (_35946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor _41925_ (_35947_, _35932_, _35946_);
  or _41926_ (_38628_, _35947_, _35945_);
  and _41927_ (_35948_, _35932_, _35838_);
  not _41928_ (_35949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor _41929_ (_35950_, _35932_, _35949_);
  or _41930_ (_38629_, _35950_, _35948_);
  and _41931_ (_35951_, _35932_, _35842_);
  not _41932_ (_35952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor _41933_ (_35953_, _35932_, _35952_);
  or _41934_ (_38630_, _35953_, _35951_);
  and _41935_ (_35954_, _35932_, _35846_);
  not _41936_ (_35955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor _41937_ (_35956_, _35932_, _35955_);
  or _41938_ (_38631_, _35956_, _35954_);
  and _41939_ (_35957_, _35904_, _35850_);
  and _41940_ (_35958_, _35957_, _35579_);
  and _41941_ (_35959_, _35958_, _35815_);
  not _41942_ (_35960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor _41943_ (_35961_, _35958_, _35960_);
  or _41944_ (_38712_, _35961_, _35959_);
  and _41945_ (_35962_, _35958_, _35822_);
  not _41946_ (_35963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor _41947_ (_35964_, _35958_, _35963_);
  or _41948_ (_38713_, _35964_, _35962_);
  and _41949_ (_35965_, _35958_, _35826_);
  not _41950_ (_35966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor _41951_ (_35967_, _35958_, _35966_);
  or _41952_ (_38714_, _35967_, _35965_);
  and _41953_ (_35968_, _35958_, _35830_);
  not _41954_ (_35969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor _41955_ (_35970_, _35958_, _35969_);
  or _41956_ (_38715_, _35970_, _35968_);
  and _41957_ (_35971_, _35958_, _35834_);
  not _41958_ (_35972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor _41959_ (_35973_, _35958_, _35972_);
  or _41960_ (_38716_, _35973_, _35971_);
  and _41961_ (_35974_, _35958_, _35838_);
  not _41962_ (_35975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor _41963_ (_35976_, _35958_, _35975_);
  or _41964_ (_38717_, _35976_, _35974_);
  and _41965_ (_35977_, _35958_, _35842_);
  not _41966_ (_35978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor _41967_ (_35979_, _35958_, _35978_);
  or _41968_ (_38718_, _35979_, _35977_);
  and _41969_ (_35980_, _35958_, _35846_);
  not _41970_ (_35981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor _41971_ (_35982_, _35958_, _35981_);
  or _41972_ (_38719_, _35982_, _35980_);
  and _41973_ (_35983_, _35904_, _35877_);
  and _41974_ (_35984_, _35983_, _35579_);
  and _41975_ (_35985_, _35984_, _35815_);
  not _41976_ (_35986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor _41977_ (_35987_, _35984_, _35986_);
  or _41978_ (_38800_, _35987_, _35985_);
  and _41979_ (_35988_, _35984_, _35822_);
  not _41980_ (_35989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor _41981_ (_35990_, _35984_, _35989_);
  or _41982_ (_38801_, _35990_, _35988_);
  and _41983_ (_35991_, _35984_, _35826_);
  not _41984_ (_35992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor _41985_ (_35993_, _35984_, _35992_);
  or _41986_ (_38802_, _35993_, _35991_);
  and _41987_ (_35994_, _35984_, _35830_);
  not _41988_ (_35995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor _41989_ (_35996_, _35984_, _35995_);
  or _41990_ (_38803_, _35996_, _35994_);
  and _41991_ (_35997_, _35984_, _35834_);
  not _41992_ (_35998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor _41993_ (_35999_, _35984_, _35998_);
  or _41994_ (_38804_, _35999_, _35997_);
  and _41995_ (_36000_, _35984_, _35838_);
  not _41996_ (_36001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor _41997_ (_36002_, _35984_, _36001_);
  or _41998_ (_38805_, _36002_, _36000_);
  and _41999_ (_36003_, _35984_, _35842_);
  not _42000_ (_36004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor _42001_ (_36005_, _35984_, _36004_);
  or _42002_ (_38806_, _36005_, _36003_);
  and _42003_ (_36006_, _35984_, _35846_);
  not _42004_ (_36007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor _42005_ (_36008_, _35984_, _36007_);
  or _42006_ (_38807_, _36008_, _36006_);
  and _42007_ (_36009_, _35570_, _34775_);
  and _42008_ (_36010_, _36009_, _35568_);
  and _42009_ (_36011_, _36010_, _35579_);
  and _42010_ (_36012_, _36011_, _35815_);
  not _42011_ (_36013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor _42012_ (_36014_, _36011_, _36013_);
  or _42013_ (_38888_, _36014_, _36012_);
  and _42014_ (_36015_, _36011_, _35822_);
  not _42015_ (_36016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor _42016_ (_36017_, _36011_, _36016_);
  or _42017_ (_38889_, _36017_, _36015_);
  and _42018_ (_36018_, _36011_, _35826_);
  not _42019_ (_36019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor _42020_ (_36020_, _36011_, _36019_);
  or _42021_ (_38890_, _36020_, _36018_);
  and _42022_ (_36021_, _36011_, _35830_);
  not _42023_ (_36022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor _42024_ (_36023_, _36011_, _36022_);
  or _42025_ (_38891_, _36023_, _36021_);
  and _42026_ (_36024_, _36011_, _35834_);
  not _42027_ (_36025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor _42028_ (_36026_, _36011_, _36025_);
  or _42029_ (_38892_, _36026_, _36024_);
  and _42030_ (_36027_, _36011_, _35838_);
  not _42031_ (_36028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor _42032_ (_36029_, _36011_, _36028_);
  or _42033_ (_38893_, _36029_, _36027_);
  and _42034_ (_36030_, _36011_, _35842_);
  not _42035_ (_36031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor _42036_ (_36032_, _36011_, _36031_);
  or _42037_ (_38894_, _36032_, _36030_);
  and _42038_ (_36033_, _36011_, _35846_);
  not _42039_ (_36034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor _42040_ (_36035_, _36011_, _36034_);
  or _42041_ (_38895_, _36035_, _36033_);
  and _42042_ (_36036_, _36009_, _35816_);
  and _42043_ (_36037_, _36036_, _35579_);
  and _42044_ (_36038_, _36037_, _35815_);
  not _42045_ (_36039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor _42046_ (_36040_, _36037_, _36039_);
  or _42047_ (_38976_, _36040_, _36038_);
  and _42048_ (_36041_, _36037_, _35822_);
  not _42049_ (_36042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor _42050_ (_36043_, _36037_, _36042_);
  or _42051_ (_38977_, _36043_, _36041_);
  and _42052_ (_36044_, _36037_, _35826_);
  not _42053_ (_36045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor _42054_ (_36046_, _36037_, _36045_);
  or _42055_ (_38978_, _36046_, _36044_);
  and _42056_ (_36047_, _36037_, _35830_);
  not _42057_ (_36048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor _42058_ (_36049_, _36037_, _36048_);
  or _42059_ (_38979_, _36049_, _36047_);
  and _42060_ (_36050_, _36037_, _35834_);
  not _42061_ (_36051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor _42062_ (_36052_, _36037_, _36051_);
  or _42063_ (_38980_, _36052_, _36050_);
  and _42064_ (_36053_, _36037_, _35838_);
  not _42065_ (_36054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor _42066_ (_36055_, _36037_, _36054_);
  or _42067_ (_38981_, _36055_, _36053_);
  and _42068_ (_36056_, _36037_, _35842_);
  not _42069_ (_36057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor _42070_ (_36058_, _36037_, _36057_);
  or _42071_ (_38982_, _36058_, _36056_);
  and _42072_ (_36059_, _36037_, _35846_);
  not _42073_ (_36060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor _42074_ (_36061_, _36037_, _36060_);
  or _42075_ (_38983_, _36061_, _36059_);
  and _42076_ (_36062_, _36009_, _35850_);
  and _42077_ (_36063_, _36062_, _35579_);
  and _42078_ (_36064_, _36063_, _35815_);
  not _42079_ (_36065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor _42080_ (_36066_, _36063_, _36065_);
  or _42081_ (_37016_, _36066_, _36064_);
  and _42082_ (_36067_, _36063_, _35822_);
  not _42083_ (_36068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor _42084_ (_36069_, _36063_, _36068_);
  or _42085_ (_37017_, _36069_, _36067_);
  and _42086_ (_36070_, _36063_, _35826_);
  not _42087_ (_36071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor _42088_ (_36072_, _36063_, _36071_);
  or _42089_ (_37018_, _36072_, _36070_);
  and _42090_ (_36073_, _36063_, _35830_);
  not _42091_ (_36074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor _42092_ (_36075_, _36063_, _36074_);
  or _42093_ (_37019_, _36075_, _36073_);
  and _42094_ (_36076_, _36063_, _35834_);
  not _42095_ (_36077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor _42096_ (_36078_, _36063_, _36077_);
  or _42097_ (_37020_, _36078_, _36076_);
  and _42098_ (_36079_, _36063_, _35838_);
  not _42099_ (_36080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor _42100_ (_36081_, _36063_, _36080_);
  or _42101_ (_37021_, _36081_, _36079_);
  and _42102_ (_36082_, _36063_, _35842_);
  not _42103_ (_36083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor _42104_ (_36084_, _36063_, _36083_);
  or _42105_ (_37022_, _36084_, _36082_);
  and _42106_ (_36085_, _36063_, _35846_);
  not _42107_ (_36086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nor _42108_ (_36087_, _36063_, _36086_);
  or _42109_ (_37023_, _36087_, _36085_);
  and _42110_ (_36088_, _36009_, _35877_);
  and _42111_ (_36089_, _36088_, _35579_);
  and _42112_ (_36090_, _36089_, _35815_);
  not _42113_ (_36091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor _42114_ (_36092_, _36089_, _36091_);
  or _42115_ (_37104_, _36092_, _36090_);
  and _42116_ (_36093_, _36089_, _35822_);
  not _42117_ (_36094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor _42118_ (_36095_, _36089_, _36094_);
  or _42119_ (_37105_, _36095_, _36093_);
  and _42120_ (_36096_, _36089_, _35826_);
  not _42121_ (_36097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor _42122_ (_36098_, _36089_, _36097_);
  or _42123_ (_37106_, _36098_, _36096_);
  and _42124_ (_36099_, _36089_, _35830_);
  not _42125_ (_36100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor _42126_ (_36101_, _36089_, _36100_);
  or _42127_ (_37107_, _36101_, _36099_);
  and _42128_ (_36102_, _36089_, _35834_);
  not _42129_ (_36103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor _42130_ (_36104_, _36089_, _36103_);
  or _42131_ (_37108_, _36104_, _36102_);
  and _42132_ (_36105_, _36089_, _35838_);
  not _42133_ (_36106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor _42134_ (_36107_, _36089_, _36106_);
  or _42135_ (_37109_, _36107_, _36105_);
  and _42136_ (_36108_, _36089_, _35842_);
  not _42137_ (_36109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor _42138_ (_36110_, _36089_, _36109_);
  or _42139_ (_37110_, _36110_, _36108_);
  and _42140_ (_36111_, _36089_, _35846_);
  not _42141_ (_36112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor _42142_ (_36113_, _36089_, _36112_);
  or _42143_ (_37111_, _36113_, _36111_);
  and _42144_ (_36114_, _35570_, _35569_);
  and _42145_ (_36115_, _36114_, _35568_);
  and _42146_ (_36116_, _36115_, _35579_);
  and _42147_ (_36117_, _36116_, _35815_);
  not _42148_ (_36118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor _42149_ (_36119_, _36116_, _36118_);
  or _42150_ (_37192_, _36119_, _36117_);
  and _42151_ (_36120_, _36116_, _35822_);
  not _42152_ (_36121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor _42153_ (_36122_, _36116_, _36121_);
  or _42154_ (_37193_, _36122_, _36120_);
  and _42155_ (_36123_, _36116_, _35826_);
  not _42156_ (_36124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor _42157_ (_36125_, _36116_, _36124_);
  or _42158_ (_37194_, _36125_, _36123_);
  and _42159_ (_36126_, _36116_, _35830_);
  not _42160_ (_36127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor _42161_ (_36128_, _36116_, _36127_);
  or _42162_ (_37195_, _36128_, _36126_);
  and _42163_ (_36129_, _36116_, _35834_);
  not _42164_ (_36130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor _42165_ (_36131_, _36116_, _36130_);
  or _42166_ (_37196_, _36131_, _36129_);
  and _42167_ (_36132_, _36116_, _35838_);
  not _42168_ (_36133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor _42169_ (_36134_, _36116_, _36133_);
  or _42170_ (_37197_, _36134_, _36132_);
  and _42171_ (_36135_, _36116_, _35842_);
  not _42172_ (_36136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor _42173_ (_36137_, _36116_, _36136_);
  or _42174_ (_37198_, _36137_, _36135_);
  and _42175_ (_36138_, _36116_, _35846_);
  not _42176_ (_36139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nor _42177_ (_36140_, _36116_, _36139_);
  or _42178_ (_37199_, _36140_, _36138_);
  and _42179_ (_36141_, _36114_, _35816_);
  and _42180_ (_36142_, _36141_, _35579_);
  and _42181_ (_36143_, _36142_, _35815_);
  not _42182_ (_36144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor _42183_ (_36145_, _36142_, _36144_);
  or _42184_ (_37280_, _36145_, _36143_);
  and _42185_ (_36146_, _36142_, _35822_);
  not _42186_ (_36147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor _42187_ (_36148_, _36142_, _36147_);
  or _42188_ (_37281_, _36148_, _36146_);
  and _42189_ (_36149_, _36142_, _35826_);
  not _42190_ (_36150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor _42191_ (_36151_, _36142_, _36150_);
  or _42192_ (_37282_, _36151_, _36149_);
  and _42193_ (_36152_, _36142_, _35830_);
  not _42194_ (_36153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor _42195_ (_36154_, _36142_, _36153_);
  or _42196_ (_37283_, _36154_, _36152_);
  and _42197_ (_36155_, _36142_, _35834_);
  not _42198_ (_36156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor _42199_ (_36157_, _36142_, _36156_);
  or _42200_ (_37284_, _36157_, _36155_);
  and _42201_ (_36158_, _36142_, _35838_);
  not _42202_ (_36159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor _42203_ (_36160_, _36142_, _36159_);
  or _42204_ (_37285_, _36160_, _36158_);
  and _42205_ (_36161_, _36142_, _35842_);
  not _42206_ (_36162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor _42207_ (_36163_, _36142_, _36162_);
  or _42208_ (_37286_, _36163_, _36161_);
  and _42209_ (_36164_, _36142_, _35846_);
  not _42210_ (_36165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor _42211_ (_36166_, _36142_, _36165_);
  or _42212_ (_37287_, _36166_, _36164_);
  and _42213_ (_36167_, _36114_, _35850_);
  and _42214_ (_36168_, _36167_, _35579_);
  and _42215_ (_36169_, _36168_, _35815_);
  not _42216_ (_36170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor _42217_ (_36171_, _36168_, _36170_);
  or _42218_ (_37368_, _36171_, _36169_);
  and _42219_ (_36172_, _36168_, _35822_);
  not _42220_ (_36173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor _42221_ (_36174_, _36168_, _36173_);
  or _42222_ (_37369_, _36174_, _36172_);
  and _42223_ (_36175_, _36168_, _35826_);
  not _42224_ (_36176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor _42225_ (_36177_, _36168_, _36176_);
  or _42226_ (_37370_, _36177_, _36175_);
  and _42227_ (_36178_, _36168_, _35830_);
  not _42228_ (_36179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor _42229_ (_36180_, _36168_, _36179_);
  or _42230_ (_37371_, _36180_, _36178_);
  and _42231_ (_36181_, _36168_, _35834_);
  not _42232_ (_36182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor _42233_ (_36183_, _36168_, _36182_);
  or _42234_ (_37372_, _36183_, _36181_);
  and _42235_ (_36184_, _36168_, _35838_);
  not _42236_ (_36185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor _42237_ (_36186_, _36168_, _36185_);
  or _42238_ (_37373_, _36186_, _36184_);
  and _42239_ (_36187_, _36168_, _35842_);
  not _42240_ (_36188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor _42241_ (_36189_, _36168_, _36188_);
  or _42242_ (_37374_, _36189_, _36187_);
  and _42243_ (_36190_, _36168_, _35846_);
  not _42244_ (_36191_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nor _42245_ (_36192_, _36168_, _36191_);
  or _42246_ (_37375_, _36192_, _36190_);
  and _42247_ (_36193_, _36114_, _35877_);
  and _42248_ (_36194_, _36193_, _35579_);
  and _42249_ (_36195_, _36194_, _35815_);
  not _42250_ (_36196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor _42251_ (_36197_, _36194_, _36196_);
  or _42252_ (_37456_, _36197_, _36195_);
  and _42253_ (_36198_, _36194_, _35822_);
  not _42254_ (_36199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor _42255_ (_36200_, _36194_, _36199_);
  or _42256_ (_37457_, _36200_, _36198_);
  and _42257_ (_36201_, _36194_, _35826_);
  not _42258_ (_36202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor _42259_ (_36203_, _36194_, _36202_);
  or _42260_ (_37458_, _36203_, _36201_);
  and _42261_ (_36204_, _36194_, _35830_);
  not _42262_ (_36205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor _42263_ (_36206_, _36194_, _36205_);
  or _42264_ (_37459_, _36206_, _36204_);
  and _42265_ (_36207_, _36194_, _35834_);
  not _42266_ (_36208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor _42267_ (_36209_, _36194_, _36208_);
  or _42268_ (_37460_, _36209_, _36207_);
  and _42269_ (_36210_, _36194_, _35838_);
  not _42270_ (_36211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor _42271_ (_36212_, _36194_, _36211_);
  or _42272_ (_37461_, _36212_, _36210_);
  and _42273_ (_36213_, _36194_, _35842_);
  not _42274_ (_36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor _42275_ (_36215_, _36194_, _36214_);
  or _42276_ (_37462_, _36215_, _36213_);
  and _42277_ (_36216_, _36194_, _35846_);
  not _42278_ (_36217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor _42279_ (_36218_, _36194_, _36217_);
  or _42280_ (_37463_, _36218_, _36216_);
  not _42281_ (_36219_, _35576_);
  and _42282_ (_36220_, _35573_, _33591_);
  and _42283_ (_36221_, _36220_, _36219_);
  and _42284_ (_36222_, _36221_, _35572_);
  and _42285_ (_36223_, _36222_, _35815_);
  not _42286_ (_36224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  nor _42287_ (_36225_, _36222_, _36224_);
  or _42288_ (_37544_, _36225_, _36223_);
  and _42289_ (_36226_, _36222_, _35822_);
  not _42290_ (_36227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  nor _42291_ (_36228_, _36222_, _36227_);
  or _42292_ (_37545_, _36228_, _36226_);
  and _42293_ (_36229_, _36222_, _35826_);
  not _42294_ (_36230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  nor _42295_ (_36231_, _36222_, _36230_);
  or _42296_ (_37546_, _36231_, _36229_);
  and _42297_ (_36232_, _36222_, _35830_);
  not _42298_ (_36233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  nor _42299_ (_36234_, _36222_, _36233_);
  or _42300_ (_37547_, _36234_, _36232_);
  and _42301_ (_36235_, _36222_, _35834_);
  not _42302_ (_36236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  nor _42303_ (_36237_, _36222_, _36236_);
  or _42304_ (_37548_, _36237_, _36235_);
  and _42305_ (_36238_, _36222_, _35838_);
  not _42306_ (_36239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  nor _42307_ (_36240_, _36222_, _36239_);
  or _42308_ (_37549_, _36240_, _36238_);
  and _42309_ (_36241_, _36222_, _35842_);
  not _42310_ (_36242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  nor _42311_ (_36243_, _36222_, _36242_);
  or _42312_ (_37550_, _36243_, _36241_);
  and _42313_ (_36244_, _36222_, _35846_);
  not _42314_ (_36245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  nor _42315_ (_36246_, _36222_, _36245_);
  or _42316_ (_37551_, _36246_, _36244_);
  and _42317_ (_36247_, _36221_, _35817_);
  and _42318_ (_36248_, _36247_, _35815_);
  not _42319_ (_36249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  nor _42320_ (_36250_, _36247_, _36249_);
  or _42321_ (_37632_, _36250_, _36248_);
  and _42322_ (_36251_, _36247_, _35822_);
  not _42323_ (_36252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  nor _42324_ (_36253_, _36247_, _36252_);
  or _42325_ (_37633_, _36253_, _36251_);
  and _42326_ (_36254_, _36247_, _35826_);
  not _42327_ (_36255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  nor _42328_ (_36256_, _36247_, _36255_);
  or _42329_ (_37634_, _36256_, _36254_);
  and _42330_ (_36257_, _36247_, _35830_);
  not _42331_ (_36258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  nor _42332_ (_36259_, _36247_, _36258_);
  or _42333_ (_37635_, _36259_, _36257_);
  and _42334_ (_36260_, _36247_, _35834_);
  not _42335_ (_36261_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  nor _42336_ (_36262_, _36247_, _36261_);
  or _42337_ (_37636_, _36262_, _36260_);
  and _42338_ (_36263_, _36247_, _35838_);
  not _42339_ (_36264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  nor _42340_ (_36265_, _36247_, _36264_);
  or _42341_ (_37637_, _36265_, _36263_);
  and _42342_ (_36266_, _36247_, _35842_);
  not _42343_ (_36267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  nor _42344_ (_36268_, _36247_, _36267_);
  or _42345_ (_37638_, _36268_, _36266_);
  and _42346_ (_36269_, _36247_, _35846_);
  not _42347_ (_36270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  nor _42348_ (_36271_, _36247_, _36270_);
  or _42349_ (_37639_, _36271_, _36269_);
  and _42350_ (_36272_, _36221_, _35851_);
  and _42351_ (_36273_, _36272_, _35815_);
  not _42352_ (_36274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  nor _42353_ (_36275_, _36272_, _36274_);
  or _42354_ (_37720_, _36275_, _36273_);
  and _42355_ (_36276_, _36272_, _35822_);
  not _42356_ (_36277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  nor _42357_ (_36278_, _36272_, _36277_);
  or _42358_ (_37721_, _36278_, _36276_);
  and _42359_ (_36279_, _36272_, _35826_);
  not _42360_ (_36280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  nor _42361_ (_36281_, _36272_, _36280_);
  or _42362_ (_37722_, _36281_, _36279_);
  and _42363_ (_36282_, _36272_, _35830_);
  not _42364_ (_36283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  nor _42365_ (_36284_, _36272_, _36283_);
  or _42366_ (_37723_, _36284_, _36282_);
  and _42367_ (_36285_, _36272_, _35834_);
  not _42368_ (_36286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  nor _42369_ (_36287_, _36272_, _36286_);
  or _42370_ (_37724_, _36287_, _36285_);
  and _42371_ (_36288_, _36272_, _35838_);
  not _42372_ (_36289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  nor _42373_ (_36290_, _36272_, _36289_);
  or _42374_ (_37725_, _36290_, _36288_);
  and _42375_ (_36291_, _36272_, _35842_);
  not _42376_ (_36292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  nor _42377_ (_36293_, _36272_, _36292_);
  or _42378_ (_37726_, _36293_, _36291_);
  and _42379_ (_36294_, _36272_, _35846_);
  not _42380_ (_36295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  nor _42381_ (_36296_, _36272_, _36295_);
  or _42382_ (_37727_, _36296_, _36294_);
  and _42383_ (_36297_, _36221_, _35878_);
  and _42384_ (_36298_, _36297_, _35815_);
  not _42385_ (_36299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  nor _42386_ (_36300_, _36297_, _36299_);
  or _42387_ (_37808_, _36300_, _36298_);
  and _42388_ (_36301_, _36297_, _35822_);
  not _42389_ (_36302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  nor _42390_ (_36303_, _36297_, _36302_);
  or _42391_ (_37809_, _36303_, _36301_);
  and _42392_ (_36304_, _36297_, _35826_);
  not _42393_ (_36305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  nor _42394_ (_36306_, _36297_, _36305_);
  or _42395_ (_37810_, _36306_, _36304_);
  and _42396_ (_36307_, _36297_, _35830_);
  not _42397_ (_36308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  nor _42398_ (_36309_, _36297_, _36308_);
  or _42399_ (_37811_, _36309_, _36307_);
  and _42400_ (_36310_, _36297_, _35834_);
  not _42401_ (_36311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  nor _42402_ (_36312_, _36297_, _36311_);
  or _42403_ (_37812_, _36312_, _36310_);
  and _42404_ (_36313_, _36297_, _35838_);
  not _42405_ (_36314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  nor _42406_ (_36315_, _36297_, _36314_);
  or _42407_ (_37813_, _36315_, _36313_);
  and _42408_ (_36316_, _36297_, _35842_);
  not _42409_ (_36317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  nor _42410_ (_36318_, _36297_, _36317_);
  or _42411_ (_37814_, _36318_, _36316_);
  and _42412_ (_36319_, _36297_, _35846_);
  not _42413_ (_36320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  nor _42414_ (_36321_, _36297_, _36320_);
  or _42415_ (_37815_, _36321_, _36319_);
  and _42416_ (_36322_, _36221_, _35905_);
  and _42417_ (_36323_, _36322_, _35815_);
  not _42418_ (_36324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  nor _42419_ (_36325_, _36322_, _36324_);
  or _42420_ (_37904_, _36325_, _36323_);
  and _42421_ (_36326_, _36322_, _35822_);
  not _42422_ (_36327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  nor _42423_ (_36328_, _36322_, _36327_);
  or _42424_ (_37905_, _36328_, _36326_);
  and _42425_ (_36329_, _36322_, _35826_);
  not _42426_ (_36330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  nor _42427_ (_36331_, _36322_, _36330_);
  or _42428_ (_37906_, _36331_, _36329_);
  and _42429_ (_36332_, _36322_, _35830_);
  not _42430_ (_36333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  nor _42431_ (_36334_, _36322_, _36333_);
  or _42432_ (_37907_, _36334_, _36332_);
  and _42433_ (_36335_, _36322_, _35834_);
  not _42434_ (_36336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  nor _42435_ (_36337_, _36322_, _36336_);
  or _42436_ (_37908_, _36337_, _36335_);
  and _42437_ (_36338_, _36322_, _35838_);
  not _42438_ (_36339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  nor _42439_ (_36340_, _36322_, _36339_);
  or _42440_ (_37909_, _36340_, _36338_);
  and _42441_ (_36341_, _36322_, _35842_);
  not _42442_ (_36342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  nor _42443_ (_36343_, _36322_, _36342_);
  or _42444_ (_37910_, _36343_, _36341_);
  and _42445_ (_36344_, _36322_, _35846_);
  not _42446_ (_36345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  nor _42447_ (_36346_, _36322_, _36345_);
  or _42448_ (_37911_, _36346_, _36344_);
  and _42449_ (_36347_, _36221_, _35931_);
  and _42450_ (_36348_, _36347_, _35815_);
  not _42451_ (_36349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  nor _42452_ (_36350_, _36347_, _36349_);
  or _42453_ (_37992_, _36350_, _36348_);
  and _42454_ (_36351_, _36347_, _35822_);
  not _42455_ (_36352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  nor _42456_ (_36353_, _36347_, _36352_);
  or _42457_ (_37993_, _36353_, _36351_);
  and _42458_ (_36354_, _36347_, _35826_);
  not _42459_ (_36355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  nor _42460_ (_36356_, _36347_, _36355_);
  or _42461_ (_37994_, _36356_, _36354_);
  and _42462_ (_36357_, _36347_, _35830_);
  not _42463_ (_36358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  nor _42464_ (_36359_, _36347_, _36358_);
  or _42465_ (_37995_, _36359_, _36357_);
  and _42466_ (_36360_, _36347_, _35834_);
  not _42467_ (_36361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  nor _42468_ (_36362_, _36347_, _36361_);
  or _42469_ (_37996_, _36362_, _36360_);
  and _42470_ (_36363_, _36347_, _35838_);
  not _42471_ (_36364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  nor _42472_ (_36365_, _36347_, _36364_);
  or _42473_ (_37997_, _36365_, _36363_);
  and _42474_ (_36366_, _36347_, _35842_);
  not _42475_ (_36367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  nor _42476_ (_36368_, _36347_, _36367_);
  or _42477_ (_37998_, _36368_, _36366_);
  and _42478_ (_36369_, _36347_, _35846_);
  not _42479_ (_36370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  nor _42480_ (_36371_, _36347_, _36370_);
  or _42481_ (_37999_, _36371_, _36369_);
  and _42482_ (_36372_, _36221_, _35957_);
  and _42483_ (_36373_, _36372_, _35815_);
  not _42484_ (_36374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  nor _42485_ (_36375_, _36372_, _36374_);
  or _42486_ (_38080_, _36375_, _36373_);
  and _42487_ (_36376_, _36372_, _35822_);
  not _42488_ (_36377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  nor _42489_ (_36378_, _36372_, _36377_);
  or _42490_ (_38081_, _36378_, _36376_);
  and _42491_ (_36379_, _36372_, _35826_);
  not _42492_ (_36380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  nor _42493_ (_36381_, _36372_, _36380_);
  or _42494_ (_38082_, _36381_, _36379_);
  and _42495_ (_36382_, _36372_, _35830_);
  not _42496_ (_36383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  nor _42497_ (_36384_, _36372_, _36383_);
  or _42498_ (_38083_, _36384_, _36382_);
  and _42499_ (_36385_, _36372_, _35834_);
  not _42500_ (_36386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  nor _42501_ (_36387_, _36372_, _36386_);
  or _42502_ (_38084_, _36387_, _36385_);
  and _42503_ (_36388_, _36372_, _35838_);
  not _42504_ (_36389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  nor _42505_ (_36390_, _36372_, _36389_);
  or _42506_ (_38085_, _36390_, _36388_);
  and _42507_ (_36391_, _36372_, _35842_);
  not _42508_ (_36392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  nor _42509_ (_36393_, _36372_, _36392_);
  or _42510_ (_38086_, _36393_, _36391_);
  and _42511_ (_36394_, _36372_, _35846_);
  not _42512_ (_36395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  nor _42513_ (_36396_, _36372_, _36395_);
  or _42514_ (_38087_, _36396_, _36394_);
  and _42515_ (_36397_, _36221_, _35983_);
  and _42516_ (_36398_, _36397_, _35815_);
  not _42517_ (_36399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  nor _42518_ (_36400_, _36397_, _36399_);
  or _42519_ (_38168_, _36400_, _36398_);
  and _42520_ (_36401_, _36397_, _35822_);
  not _42521_ (_36402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  nor _42522_ (_36403_, _36397_, _36402_);
  or _42523_ (_38169_, _36403_, _36401_);
  and _42524_ (_36404_, _36397_, _35826_);
  not _42525_ (_36405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  nor _42526_ (_36406_, _36397_, _36405_);
  or _42527_ (_38170_, _36406_, _36404_);
  and _42528_ (_36407_, _36397_, _35830_);
  not _42529_ (_36408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  nor _42530_ (_36409_, _36397_, _36408_);
  or _42531_ (_38171_, _36409_, _36407_);
  and _42532_ (_36410_, _36397_, _35834_);
  not _42533_ (_36411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  nor _42534_ (_36412_, _36397_, _36411_);
  or _42535_ (_38172_, _36412_, _36410_);
  and _42536_ (_36413_, _36397_, _35838_);
  not _42537_ (_36414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  nor _42538_ (_36415_, _36397_, _36414_);
  or _42539_ (_38173_, _36415_, _36413_);
  and _42540_ (_36416_, _36397_, _35842_);
  not _42541_ (_36417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  nor _42542_ (_36418_, _36397_, _36417_);
  or _42543_ (_38174_, _36418_, _36416_);
  and _42544_ (_36419_, _36397_, _35846_);
  not _42545_ (_36420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  nor _42546_ (_36421_, _36397_, _36420_);
  or _42547_ (_38175_, _36421_, _36419_);
  and _42548_ (_36422_, _36221_, _36010_);
  and _42549_ (_36423_, _36422_, _35815_);
  not _42550_ (_36424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  nor _42551_ (_36425_, _36422_, _36424_);
  or _42552_ (_38256_, _36425_, _36423_);
  and _42553_ (_36426_, _36422_, _35822_);
  not _42554_ (_36427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  nor _42555_ (_36428_, _36422_, _36427_);
  or _42556_ (_38257_, _36428_, _36426_);
  and _42557_ (_36429_, _36422_, _35826_);
  not _42558_ (_36430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  nor _42559_ (_36431_, _36422_, _36430_);
  or _42560_ (_38258_, _36431_, _36429_);
  and _42561_ (_36432_, _36422_, _35830_);
  not _42562_ (_36433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  nor _42563_ (_36434_, _36422_, _36433_);
  or _42564_ (_38259_, _36434_, _36432_);
  and _42565_ (_36435_, _36422_, _35834_);
  not _42566_ (_36436_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  nor _42567_ (_36437_, _36422_, _36436_);
  or _42568_ (_38260_, _36437_, _36435_);
  and _42569_ (_36438_, _36422_, _35838_);
  not _42570_ (_36439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  nor _42571_ (_36440_, _36422_, _36439_);
  or _42572_ (_38261_, _36440_, _36438_);
  and _42573_ (_36441_, _36422_, _35842_);
  not _42574_ (_36442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  nor _42575_ (_36443_, _36422_, _36442_);
  or _42576_ (_38262_, _36443_, _36441_);
  and _42577_ (_36444_, _36422_, _35846_);
  not _42578_ (_36445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  nor _42579_ (_36446_, _36422_, _36445_);
  or _42580_ (_38263_, _36446_, _36444_);
  and _42581_ (_36447_, _36221_, _36036_);
  and _42582_ (_36448_, _36447_, _35815_);
  not _42583_ (_36449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  nor _42584_ (_36450_, _36447_, _36449_);
  or _42585_ (_38320_, _36450_, _36448_);
  and _42586_ (_36451_, _36447_, _35822_);
  not _42587_ (_36452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  nor _42588_ (_36453_, _36447_, _36452_);
  or _42589_ (_38321_, _36453_, _36451_);
  and _42590_ (_36454_, _36447_, _35826_);
  not _42591_ (_36455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  nor _42592_ (_36456_, _36447_, _36455_);
  or _42593_ (_38322_, _36456_, _36454_);
  and _42594_ (_36457_, _36447_, _35830_);
  not _42595_ (_36458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  nor _42596_ (_36459_, _36447_, _36458_);
  or _42597_ (_38323_, _36459_, _36457_);
  and _42598_ (_36460_, _36447_, _35834_);
  not _42599_ (_36461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  nor _42600_ (_36462_, _36447_, _36461_);
  or _42601_ (_38324_, _36462_, _36460_);
  and _42602_ (_36463_, _36447_, _35838_);
  not _42603_ (_36464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  nor _42604_ (_36465_, _36447_, _36464_);
  or _42605_ (_38325_, _36465_, _36463_);
  and _42606_ (_36466_, _36447_, _35842_);
  not _42607_ (_36467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  nor _42608_ (_36468_, _36447_, _36467_);
  or _42609_ (_38326_, _36468_, _36466_);
  and _42610_ (_36469_, _36447_, _35846_);
  not _42611_ (_36470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  nor _42612_ (_36471_, _36447_, _36470_);
  or _42613_ (_38327_, _36471_, _36469_);
  and _42614_ (_36472_, _36221_, _36062_);
  and _42615_ (_36473_, _36472_, _35815_);
  not _42616_ (_36474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  nor _42617_ (_36475_, _36472_, _36474_);
  or _42618_ (_38328_, _36475_, _36473_);
  and _42619_ (_36476_, _36472_, _35822_);
  not _42620_ (_36477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  nor _42621_ (_36478_, _36472_, _36477_);
  or _42622_ (_38329_, _36478_, _36476_);
  and _42623_ (_36479_, _36472_, _35826_);
  not _42624_ (_36480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  nor _42625_ (_36481_, _36472_, _36480_);
  or _42626_ (_38330_, _36481_, _36479_);
  and _42627_ (_36482_, _36472_, _35830_);
  not _42628_ (_36483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  nor _42629_ (_36484_, _36472_, _36483_);
  or _42630_ (_38331_, _36484_, _36482_);
  and _42631_ (_36485_, _36472_, _35834_);
  not _42632_ (_36486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  nor _42633_ (_36487_, _36472_, _36486_);
  or _42634_ (_38332_, _36487_, _36485_);
  and _42635_ (_36488_, _36472_, _35838_);
  not _42636_ (_36489_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  nor _42637_ (_36490_, _36472_, _36489_);
  or _42638_ (_38333_, _36490_, _36488_);
  and _42639_ (_36491_, _36472_, _35842_);
  not _42640_ (_36492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  nor _42641_ (_36493_, _36472_, _36492_);
  or _42642_ (_38334_, _36493_, _36491_);
  and _42643_ (_36494_, _36472_, _35846_);
  not _42644_ (_36495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  nor _42645_ (_36496_, _36472_, _36495_);
  or _42646_ (_38335_, _36496_, _36494_);
  and _42647_ (_36497_, _36221_, _36088_);
  and _42648_ (_36498_, _36497_, _35815_);
  not _42649_ (_36499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  nor _42650_ (_36500_, _36497_, _36499_);
  or _42651_ (_38336_, _36500_, _36498_);
  and _42652_ (_36501_, _36497_, _35822_);
  not _42653_ (_36502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  nor _42654_ (_36503_, _36497_, _36502_);
  or _42655_ (_38337_, _36503_, _36501_);
  and _42656_ (_36504_, _36497_, _35826_);
  not _42657_ (_36505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  nor _42658_ (_36506_, _36497_, _36505_);
  or _42659_ (_38338_, _36506_, _36504_);
  and _42660_ (_36507_, _36497_, _35830_);
  not _42661_ (_36508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  nor _42662_ (_36509_, _36497_, _36508_);
  or _42663_ (_38339_, _36509_, _36507_);
  and _42664_ (_36510_, _36497_, _35834_);
  not _42665_ (_36511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  nor _42666_ (_36512_, _36497_, _36511_);
  or _42667_ (_38340_, _36512_, _36510_);
  and _42668_ (_36513_, _36497_, _35838_);
  not _42669_ (_36514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  nor _42670_ (_36515_, _36497_, _36514_);
  or _42671_ (_38341_, _36515_, _36513_);
  and _42672_ (_36516_, _36497_, _35842_);
  not _42673_ (_36517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  nor _42674_ (_36518_, _36497_, _36517_);
  or _42675_ (_38342_, _36518_, _36516_);
  and _42676_ (_36519_, _36497_, _35846_);
  not _42677_ (_36520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  nor _42678_ (_36521_, _36497_, _36520_);
  or _42679_ (_38343_, _36521_, _36519_);
  and _42680_ (_36522_, _36221_, _36115_);
  and _42681_ (_36523_, _36522_, _35815_);
  not _42682_ (_36524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  nor _42683_ (_36525_, _36522_, _36524_);
  or _42684_ (_38344_, _36525_, _36523_);
  and _42685_ (_36526_, _36522_, _35822_);
  not _42686_ (_36527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  nor _42687_ (_36528_, _36522_, _36527_);
  or _42688_ (_38345_, _36528_, _36526_);
  and _42689_ (_36529_, _36522_, _35826_);
  not _42690_ (_36530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  nor _42691_ (_36531_, _36522_, _36530_);
  or _42692_ (_38346_, _36531_, _36529_);
  and _42693_ (_36532_, _36522_, _35830_);
  not _42694_ (_36533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  nor _42695_ (_36534_, _36522_, _36533_);
  or _42696_ (_38347_, _36534_, _36532_);
  and _42697_ (_36535_, _36522_, _35834_);
  not _42698_ (_36536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  nor _42699_ (_36537_, _36522_, _36536_);
  or _42700_ (_38348_, _36537_, _36535_);
  and _42701_ (_36538_, _36522_, _35838_);
  not _42702_ (_36539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  nor _42703_ (_36540_, _36522_, _36539_);
  or _42704_ (_38349_, _36540_, _36538_);
  and _42705_ (_36541_, _36522_, _35842_);
  not _42706_ (_36542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  nor _42707_ (_36543_, _36522_, _36542_);
  or _42708_ (_38350_, _36543_, _36541_);
  and _42709_ (_36544_, _36522_, _35846_);
  not _42710_ (_36545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  nor _42711_ (_36546_, _36522_, _36545_);
  or _42712_ (_38351_, _36546_, _36544_);
  and _42713_ (_36547_, _36221_, _36141_);
  and _42714_ (_36548_, _36547_, _35815_);
  not _42715_ (_36549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  nor _42716_ (_36550_, _36547_, _36549_);
  or _42717_ (_38352_, _36550_, _36548_);
  and _42718_ (_36551_, _36547_, _35822_);
  not _42719_ (_36552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  nor _42720_ (_36553_, _36547_, _36552_);
  or _42721_ (_38353_, _36553_, _36551_);
  and _42722_ (_36554_, _36547_, _35826_);
  not _42723_ (_36555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  nor _42724_ (_36556_, _36547_, _36555_);
  or _42725_ (_38354_, _36556_, _36554_);
  and _42726_ (_36557_, _36547_, _35830_);
  not _42727_ (_36558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  nor _42728_ (_36559_, _36547_, _36558_);
  or _42729_ (_38355_, _36559_, _36557_);
  and _42730_ (_36560_, _36547_, _35834_);
  not _42731_ (_36561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  nor _42732_ (_36562_, _36547_, _36561_);
  or _42733_ (_38356_, _36562_, _36560_);
  and _42734_ (_36563_, _36547_, _35838_);
  not _42735_ (_36564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  nor _42736_ (_36565_, _36547_, _36564_);
  or _42737_ (_38357_, _36565_, _36563_);
  and _42738_ (_36566_, _36547_, _35842_);
  not _42739_ (_36567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  nor _42740_ (_36568_, _36547_, _36567_);
  or _42741_ (_38358_, _36568_, _36566_);
  and _42742_ (_36569_, _36547_, _35846_);
  not _42743_ (_36570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  nor _42744_ (_36571_, _36547_, _36570_);
  or _42745_ (_38359_, _36571_, _36569_);
  and _42746_ (_36572_, _36221_, _36167_);
  and _42747_ (_36573_, _36572_, _35815_);
  not _42748_ (_36574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  nor _42749_ (_36575_, _36572_, _36574_);
  or _42750_ (_38368_, _36575_, _36573_);
  and _42751_ (_36576_, _36572_, _35822_);
  not _42752_ (_36577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  nor _42753_ (_36578_, _36572_, _36577_);
  or _42754_ (_38369_, _36578_, _36576_);
  and _42755_ (_36579_, _36572_, _35826_);
  not _42756_ (_36580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  nor _42757_ (_36581_, _36572_, _36580_);
  or _42758_ (_38370_, _36581_, _36579_);
  and _42759_ (_36582_, _36572_, _35830_);
  not _42760_ (_36583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  nor _42761_ (_36584_, _36572_, _36583_);
  or _42762_ (_38371_, _36584_, _36582_);
  and _42763_ (_36585_, _36572_, _35834_);
  not _42764_ (_36586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  nor _42765_ (_36587_, _36572_, _36586_);
  or _42766_ (_38372_, _36587_, _36585_);
  and _42767_ (_36588_, _36572_, _35838_);
  not _42768_ (_36589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  nor _42769_ (_36590_, _36572_, _36589_);
  or _42770_ (_38373_, _36590_, _36588_);
  and _42771_ (_36591_, _36572_, _35842_);
  not _42772_ (_36592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  nor _42773_ (_36593_, _36572_, _36592_);
  or _42774_ (_38374_, _36593_, _36591_);
  and _42775_ (_36594_, _36572_, _35846_);
  not _42776_ (_36595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  nor _42777_ (_36596_, _36572_, _36595_);
  or _42778_ (_38375_, _36596_, _36594_);
  and _42779_ (_36597_, _36221_, _36193_);
  and _42780_ (_36598_, _36597_, _35815_);
  not _42781_ (_36599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  nor _42782_ (_36600_, _36597_, _36599_);
  or _42783_ (_38376_, _36600_, _36598_);
  and _42784_ (_36601_, _36597_, _35822_);
  not _42785_ (_36602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  nor _42786_ (_36603_, _36597_, _36602_);
  or _42787_ (_38377_, _36603_, _36601_);
  and _42788_ (_36604_, _36597_, _35826_);
  not _42789_ (_36605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  nor _42790_ (_36606_, _36597_, _36605_);
  or _42791_ (_38378_, _36606_, _36604_);
  and _42792_ (_36607_, _36597_, _35830_);
  not _42793_ (_36608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  nor _42794_ (_36609_, _36597_, _36608_);
  or _42795_ (_38379_, _36609_, _36607_);
  and _42796_ (_36610_, _36597_, _35834_);
  not _42797_ (_36611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  nor _42798_ (_36612_, _36597_, _36611_);
  or _42799_ (_38380_, _36612_, _36610_);
  and _42800_ (_36613_, _36597_, _35838_);
  not _42801_ (_36614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  nor _42802_ (_36615_, _36597_, _36614_);
  or _42803_ (_38381_, _36615_, _36613_);
  and _42804_ (_36616_, _36597_, _35842_);
  not _42805_ (_36617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  nor _42806_ (_36618_, _36597_, _36617_);
  or _42807_ (_38382_, _36618_, _36616_);
  and _42808_ (_36619_, _36597_, _35846_);
  not _42809_ (_36620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  nor _42810_ (_36621_, _36597_, _36620_);
  or _42811_ (_38383_, _36621_, _36619_);
  and _42812_ (_36622_, _35574_, _34702_);
  and _42813_ (_36623_, _36622_, _36219_);
  and _42814_ (_36624_, _36623_, _35572_);
  and _42815_ (_36625_, _36624_, _35815_);
  not _42816_ (_36626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  nor _42817_ (_36627_, _36624_, _36626_);
  or _42818_ (_38384_, _36627_, _36625_);
  and _42819_ (_36628_, _36624_, _35822_);
  not _42820_ (_36629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  nor _42821_ (_36630_, _36624_, _36629_);
  or _42822_ (_38385_, _36630_, _36628_);
  and _42823_ (_36631_, _36624_, _35826_);
  not _42824_ (_36632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  nor _42825_ (_36633_, _36624_, _36632_);
  or _42826_ (_38386_, _36633_, _36631_);
  and _42827_ (_36634_, _36624_, _35830_);
  not _42828_ (_36635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  nor _42829_ (_36636_, _36624_, _36635_);
  or _42830_ (_38387_, _36636_, _36634_);
  and _42831_ (_36637_, _36624_, _35834_);
  not _42832_ (_36638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  nor _42833_ (_36639_, _36624_, _36638_);
  or _42834_ (_38388_, _36639_, _36637_);
  and _42835_ (_36640_, _36624_, _35838_);
  not _42836_ (_36641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  nor _42837_ (_36642_, _36624_, _36641_);
  or _42838_ (_38389_, _36642_, _36640_);
  and _42839_ (_36643_, _36624_, _35842_);
  not _42840_ (_36644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  nor _42841_ (_36645_, _36624_, _36644_);
  or _42842_ (_38390_, _36645_, _36643_);
  and _42843_ (_36646_, _36624_, _35846_);
  not _42844_ (_36647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  nor _42845_ (_36648_, _36624_, _36647_);
  or _42846_ (_38391_, _36648_, _36646_);
  and _42847_ (_36649_, _36623_, _35817_);
  and _42848_ (_36650_, _36649_, _35815_);
  not _42849_ (_36651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  nor _42850_ (_36652_, _36649_, _36651_);
  or _42851_ (_38392_, _36652_, _36650_);
  and _42852_ (_36653_, _36649_, _35822_);
  not _42853_ (_36654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  nor _42854_ (_36655_, _36649_, _36654_);
  or _42855_ (_38393_, _36655_, _36653_);
  and _42856_ (_36656_, _36649_, _35826_);
  not _42857_ (_36657_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  nor _42858_ (_36658_, _36649_, _36657_);
  or _42859_ (_38394_, _36658_, _36656_);
  and _42860_ (_36659_, _36649_, _35830_);
  not _42861_ (_36660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  nor _42862_ (_36661_, _36649_, _36660_);
  or _42863_ (_38395_, _36661_, _36659_);
  and _42864_ (_36662_, _36649_, _35834_);
  not _42865_ (_36663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  nor _42866_ (_36664_, _36649_, _36663_);
  or _42867_ (_38396_, _36664_, _36662_);
  and _42868_ (_36665_, _36649_, _35838_);
  not _42869_ (_36666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  nor _42870_ (_36667_, _36649_, _36666_);
  or _42871_ (_38397_, _36667_, _36665_);
  and _42872_ (_36668_, _36649_, _35842_);
  not _42873_ (_36669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  nor _42874_ (_36670_, _36649_, _36669_);
  or _42875_ (_38398_, _36670_, _36668_);
  and _42876_ (_36671_, _36649_, _35846_);
  not _42877_ (_36672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  nor _42878_ (_36673_, _36649_, _36672_);
  or _42879_ (_38399_, _36673_, _36671_);
  and _42880_ (_36674_, _36623_, _35851_);
  and _42881_ (_36675_, _36674_, _35815_);
  not _42882_ (_36676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  nor _42883_ (_36677_, _36674_, _36676_);
  or _42884_ (_38400_, _36677_, _36675_);
  and _42885_ (_36678_, _36674_, _35822_);
  not _42886_ (_36679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  nor _42887_ (_36680_, _36674_, _36679_);
  or _42888_ (_38401_, _36680_, _36678_);
  and _42889_ (_36681_, _36674_, _35826_);
  not _42890_ (_36682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  nor _42891_ (_36683_, _36674_, _36682_);
  or _42892_ (_38402_, _36683_, _36681_);
  and _42893_ (_36684_, _36674_, _35830_);
  not _42894_ (_36685_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  nor _42895_ (_36686_, _36674_, _36685_);
  or _42896_ (_38403_, _36686_, _36684_);
  and _42897_ (_36687_, _36674_, _35834_);
  not _42898_ (_36688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  nor _42899_ (_36689_, _36674_, _36688_);
  or _42900_ (_38404_, _36689_, _36687_);
  and _42901_ (_36690_, _36674_, _35838_);
  not _42902_ (_36691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  nor _42903_ (_36692_, _36674_, _36691_);
  or _42904_ (_38405_, _36692_, _36690_);
  and _42905_ (_36693_, _36674_, _35842_);
  not _42906_ (_36694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  nor _42907_ (_36695_, _36674_, _36694_);
  or _42908_ (_38406_, _36695_, _36693_);
  and _42909_ (_36696_, _36674_, _35846_);
  not _42910_ (_36697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  nor _42911_ (_36698_, _36674_, _36697_);
  or _42912_ (_38407_, _36698_, _36696_);
  and _42913_ (_36699_, _36623_, _35878_);
  and _42914_ (_36700_, _36699_, _35815_);
  not _42915_ (_36701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  nor _42916_ (_36702_, _36699_, _36701_);
  or _42917_ (_38408_, _36702_, _36700_);
  and _42918_ (_36703_, _36699_, _35822_);
  not _42919_ (_36704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  nor _42920_ (_36705_, _36699_, _36704_);
  or _42921_ (_38409_, _36705_, _36703_);
  and _42922_ (_36706_, _36699_, _35826_);
  not _42923_ (_36707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  nor _42924_ (_36708_, _36699_, _36707_);
  or _42925_ (_38410_, _36708_, _36706_);
  and _42926_ (_36709_, _36699_, _35830_);
  not _42927_ (_36710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  nor _42928_ (_36711_, _36699_, _36710_);
  or _42929_ (_38411_, _36711_, _36709_);
  and _42930_ (_36712_, _36699_, _35834_);
  not _42931_ (_36713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  nor _42932_ (_36714_, _36699_, _36713_);
  or _42933_ (_38412_, _36714_, _36712_);
  and _42934_ (_36715_, _36699_, _35838_);
  not _42935_ (_36716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  nor _42936_ (_36717_, _36699_, _36716_);
  or _42937_ (_38413_, _36717_, _36715_);
  and _42938_ (_36718_, _36699_, _35842_);
  not _42939_ (_36719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  nor _42940_ (_36720_, _36699_, _36719_);
  or _42941_ (_38414_, _36720_, _36718_);
  and _42942_ (_36721_, _36699_, _35846_);
  not _42943_ (_36722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  nor _42944_ (_36723_, _36699_, _36722_);
  or _42945_ (_38415_, _36723_, _36721_);
  and _42946_ (_36724_, _36623_, _35905_);
  and _42947_ (_36725_, _36724_, _35815_);
  not _42948_ (_36726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  nor _42949_ (_36727_, _36724_, _36726_);
  or _42950_ (_38416_, _36727_, _36725_);
  and _42951_ (_36728_, _36724_, _35822_);
  not _42952_ (_00009_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  nor _42953_ (_00010_, _36724_, _00009_);
  or _42954_ (_38417_, _00010_, _36728_);
  and _42955_ (_00011_, _36724_, _35826_);
  not _42956_ (_00012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  nor _42957_ (_00013_, _36724_, _00012_);
  or _42958_ (_38418_, _00013_, _00011_);
  and _42959_ (_00014_, _36724_, _35830_);
  not _42960_ (_00015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  nor _42961_ (_00016_, _36724_, _00015_);
  or _42962_ (_38419_, _00016_, _00014_);
  and _42963_ (_00017_, _36724_, _35834_);
  not _42964_ (_00018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  nor _42965_ (_00019_, _36724_, _00018_);
  or _42966_ (_38420_, _00019_, _00017_);
  and _42967_ (_00020_, _36724_, _35838_);
  not _42968_ (_00021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  nor _42969_ (_00022_, _36724_, _00021_);
  or _42970_ (_38421_, _00022_, _00020_);
  and _42971_ (_00023_, _36724_, _35842_);
  not _42972_ (_00024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  nor _42973_ (_00025_, _36724_, _00024_);
  or _42974_ (_38422_, _00025_, _00023_);
  and _42975_ (_00026_, _36724_, _35846_);
  not _42976_ (_00027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  nor _42977_ (_00028_, _36724_, _00027_);
  or _42978_ (_38423_, _00028_, _00026_);
  and _42979_ (_00029_, _36623_, _35931_);
  and _42980_ (_00030_, _00029_, _35815_);
  not _42981_ (_00031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  nor _42982_ (_00032_, _00029_, _00031_);
  or _42983_ (_38424_, _00032_, _00030_);
  and _42984_ (_00033_, _00029_, _35822_);
  not _42985_ (_00034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  nor _42986_ (_00035_, _00029_, _00034_);
  or _42987_ (_38425_, _00035_, _00033_);
  and _42988_ (_00036_, _00029_, _35826_);
  not _42989_ (_00037_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  nor _42990_ (_00038_, _00029_, _00037_);
  or _42991_ (_38426_, _00038_, _00036_);
  and _42992_ (_00039_, _00029_, _35830_);
  not _42993_ (_00040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  nor _42994_ (_00041_, _00029_, _00040_);
  or _42995_ (_38427_, _00041_, _00039_);
  and _42996_ (_00042_, _00029_, _35834_);
  not _42997_ (_00043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  nor _42998_ (_00044_, _00029_, _00043_);
  or _42999_ (_38428_, _00044_, _00042_);
  and _43000_ (_00045_, _00029_, _35838_);
  not _43001_ (_00046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  nor _43002_ (_00047_, _00029_, _00046_);
  or _43003_ (_38429_, _00047_, _00045_);
  and _43004_ (_00048_, _00029_, _35842_);
  not _43005_ (_00049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  nor _43006_ (_00050_, _00029_, _00049_);
  or _43007_ (_38430_, _00050_, _00048_);
  and _43008_ (_00051_, _00029_, _35846_);
  not _43009_ (_00052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  nor _43010_ (_00053_, _00029_, _00052_);
  or _43011_ (_38431_, _00053_, _00051_);
  and _43012_ (_00054_, _36623_, _35957_);
  and _43013_ (_00055_, _00054_, _35815_);
  not _43014_ (_00056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  nor _43015_ (_00057_, _00054_, _00056_);
  or _43016_ (_38432_, _00057_, _00055_);
  and _43017_ (_00058_, _00054_, _35822_);
  not _43018_ (_00059_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  nor _43019_ (_00060_, _00054_, _00059_);
  or _43020_ (_38433_, _00060_, _00058_);
  and _43021_ (_00061_, _00054_, _35826_);
  not _43022_ (_00062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  nor _43023_ (_00063_, _00054_, _00062_);
  or _43024_ (_38434_, _00063_, _00061_);
  and _43025_ (_00064_, _00054_, _35830_);
  not _43026_ (_00065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  nor _43027_ (_00066_, _00054_, _00065_);
  or _43028_ (_38435_, _00066_, _00064_);
  and _43029_ (_00067_, _00054_, _35834_);
  not _43030_ (_00068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  nor _43031_ (_00069_, _00054_, _00068_);
  or _43032_ (_38436_, _00069_, _00067_);
  and _43033_ (_00070_, _00054_, _35838_);
  not _43034_ (_00071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  nor _43035_ (_00072_, _00054_, _00071_);
  or _43036_ (_38437_, _00072_, _00070_);
  and _43037_ (_00073_, _00054_, _35842_);
  not _43038_ (_00074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  nor _43039_ (_00075_, _00054_, _00074_);
  or _43040_ (_38438_, _00075_, _00073_);
  and _43041_ (_00076_, _00054_, _35846_);
  not _43042_ (_00077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  nor _43043_ (_00078_, _00054_, _00077_);
  or _43044_ (_38439_, _00078_, _00076_);
  and _43045_ (_00079_, _36623_, _35983_);
  and _43046_ (_00080_, _00079_, _35815_);
  not _43047_ (_00081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  nor _43048_ (_00082_, _00079_, _00081_);
  or _43049_ (_38440_, _00082_, _00080_);
  and _43050_ (_00083_, _00079_, _35822_);
  not _43051_ (_00084_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  nor _43052_ (_00085_, _00079_, _00084_);
  or _43053_ (_38441_, _00085_, _00083_);
  and _43054_ (_00086_, _00079_, _35826_);
  not _43055_ (_00087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  nor _43056_ (_00088_, _00079_, _00087_);
  or _43057_ (_38442_, _00088_, _00086_);
  and _43058_ (_00089_, _00079_, _35830_);
  not _43059_ (_00090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  nor _43060_ (_00091_, _00079_, _00090_);
  or _43061_ (_38443_, _00091_, _00089_);
  and _43062_ (_00092_, _00079_, _35834_);
  not _43063_ (_00093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  nor _43064_ (_00094_, _00079_, _00093_);
  or _43065_ (_38444_, _00094_, _00092_);
  and _43066_ (_00095_, _00079_, _35838_);
  not _43067_ (_00096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  nor _43068_ (_00097_, _00079_, _00096_);
  or _43069_ (_38445_, _00097_, _00095_);
  and _43070_ (_00098_, _00079_, _35842_);
  not _43071_ (_00099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  nor _43072_ (_00100_, _00079_, _00099_);
  or _43073_ (_38446_, _00100_, _00098_);
  and _43074_ (_00101_, _00079_, _35846_);
  not _43075_ (_00102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  nor _43076_ (_00103_, _00079_, _00102_);
  or _43077_ (_38447_, _00103_, _00101_);
  and _43078_ (_00104_, _36623_, _36010_);
  and _43079_ (_00105_, _00104_, _35815_);
  not _43080_ (_00106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  nor _43081_ (_00107_, _00104_, _00106_);
  or _43082_ (_38456_, _00107_, _00105_);
  and _43083_ (_00108_, _00104_, _35822_);
  not _43084_ (_00109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  nor _43085_ (_00110_, _00104_, _00109_);
  or _43086_ (_38457_, _00110_, _00108_);
  and _43087_ (_00111_, _00104_, _35826_);
  not _43088_ (_00112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  nor _43089_ (_00113_, _00104_, _00112_);
  or _43090_ (_38458_, _00113_, _00111_);
  and _43091_ (_00114_, _00104_, _35830_);
  not _43092_ (_00115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  nor _43093_ (_00116_, _00104_, _00115_);
  or _43094_ (_38459_, _00116_, _00114_);
  and _43095_ (_00117_, _00104_, _35834_);
  not _43096_ (_00118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  nor _43097_ (_00119_, _00104_, _00118_);
  or _43098_ (_38460_, _00119_, _00117_);
  and _43099_ (_00120_, _00104_, _35838_);
  not _43100_ (_00121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  nor _43101_ (_00122_, _00104_, _00121_);
  or _43102_ (_38461_, _00122_, _00120_);
  and _43103_ (_00123_, _00104_, _35842_);
  not _43104_ (_00124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  nor _43105_ (_00125_, _00104_, _00124_);
  or _43106_ (_38462_, _00125_, _00123_);
  and _43107_ (_00126_, _00104_, _35846_);
  not _43108_ (_00127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  nor _43109_ (_00128_, _00104_, _00127_);
  or _43110_ (_38463_, _00128_, _00126_);
  and _43111_ (_00129_, _36623_, _36036_);
  and _43112_ (_00130_, _00129_, _35815_);
  not _43113_ (_00131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  nor _43114_ (_00132_, _00129_, _00131_);
  or _43115_ (_38464_, _00132_, _00130_);
  and _43116_ (_00133_, _00129_, _35822_);
  not _43117_ (_00134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  nor _43118_ (_00135_, _00129_, _00134_);
  or _43119_ (_38465_, _00135_, _00133_);
  and _43120_ (_00136_, _00129_, _35826_);
  not _43121_ (_00137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  nor _43122_ (_00138_, _00129_, _00137_);
  or _43123_ (_38466_, _00138_, _00136_);
  and _43124_ (_00139_, _00129_, _35830_);
  not _43125_ (_00140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  nor _43126_ (_00141_, _00129_, _00140_);
  or _43127_ (_38467_, _00141_, _00139_);
  and _43128_ (_00142_, _00129_, _35834_);
  not _43129_ (_00143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  nor _43130_ (_00144_, _00129_, _00143_);
  or _43131_ (_38468_, _00144_, _00142_);
  and _43132_ (_00145_, _00129_, _35838_);
  not _43133_ (_00146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  nor _43134_ (_00147_, _00129_, _00146_);
  or _43135_ (_38469_, _00147_, _00145_);
  and _43136_ (_00148_, _00129_, _35842_);
  not _43137_ (_00149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  nor _43138_ (_00150_, _00129_, _00149_);
  or _43139_ (_38470_, _00150_, _00148_);
  and _43140_ (_00151_, _00129_, _35846_);
  not _43141_ (_00152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  nor _43142_ (_00153_, _00129_, _00152_);
  or _43143_ (_38471_, _00153_, _00151_);
  and _43144_ (_00154_, _36623_, _36062_);
  and _43145_ (_00155_, _00154_, _35815_);
  not _43146_ (_00156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  nor _43147_ (_00157_, _00154_, _00156_);
  or _43148_ (_38472_, _00157_, _00155_);
  and _43149_ (_00158_, _00154_, _35822_);
  not _43150_ (_00159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  nor _43151_ (_00160_, _00154_, _00159_);
  or _43152_ (_38473_, _00160_, _00158_);
  and _43153_ (_00161_, _00154_, _35826_);
  not _43154_ (_00162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  nor _43155_ (_00163_, _00154_, _00162_);
  or _43156_ (_38474_, _00163_, _00161_);
  and _43157_ (_00164_, _00154_, _35830_);
  not _43158_ (_00165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  nor _43159_ (_00166_, _00154_, _00165_);
  or _43160_ (_38475_, _00166_, _00164_);
  and _43161_ (_00167_, _00154_, _35834_);
  not _43162_ (_00168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  nor _43163_ (_00169_, _00154_, _00168_);
  or _43164_ (_38476_, _00169_, _00167_);
  and _43165_ (_00170_, _00154_, _35838_);
  not _43166_ (_00171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  nor _43167_ (_00172_, _00154_, _00171_);
  or _43168_ (_38477_, _00172_, _00170_);
  and _43169_ (_00173_, _00154_, _35842_);
  not _43170_ (_00174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  nor _43171_ (_00175_, _00154_, _00174_);
  or _43172_ (_38478_, _00175_, _00173_);
  and _43173_ (_00176_, _00154_, _35846_);
  not _43174_ (_00177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  nor _43175_ (_00178_, _00154_, _00177_);
  or _43176_ (_38479_, _00178_, _00176_);
  and _43177_ (_00179_, _36623_, _36088_);
  and _43178_ (_00180_, _00179_, _35815_);
  not _43179_ (_00181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  nor _43180_ (_00182_, _00179_, _00181_);
  or _43181_ (_38480_, _00182_, _00180_);
  and _43182_ (_00183_, _00179_, _35822_);
  not _43183_ (_00184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  nor _43184_ (_00185_, _00179_, _00184_);
  or _43185_ (_38481_, _00185_, _00183_);
  and _43186_ (_00186_, _00179_, _35826_);
  not _43187_ (_00187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  nor _43188_ (_00188_, _00179_, _00187_);
  or _43189_ (_38482_, _00188_, _00186_);
  and _43190_ (_00189_, _00179_, _35830_);
  not _43191_ (_00190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  nor _43192_ (_00191_, _00179_, _00190_);
  or _43193_ (_38483_, _00191_, _00189_);
  and _43194_ (_00192_, _00179_, _35834_);
  not _43195_ (_00193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  nor _43196_ (_00194_, _00179_, _00193_);
  or _43197_ (_38484_, _00194_, _00192_);
  and _43198_ (_00195_, _00179_, _35838_);
  not _43199_ (_00196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  nor _43200_ (_00197_, _00179_, _00196_);
  or _43201_ (_38485_, _00197_, _00195_);
  and _43202_ (_00198_, _00179_, _35842_);
  not _43203_ (_00199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  nor _43204_ (_00200_, _00179_, _00199_);
  or _43205_ (_38486_, _00200_, _00198_);
  and _43206_ (_00201_, _00179_, _35846_);
  not _43207_ (_00202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  nor _43208_ (_00203_, _00179_, _00202_);
  or _43209_ (_38487_, _00203_, _00201_);
  and _43210_ (_00204_, _36623_, _36115_);
  and _43211_ (_00205_, _00204_, _35815_);
  not _43212_ (_00206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  nor _43213_ (_00207_, _00204_, _00206_);
  or _43214_ (_38488_, _00207_, _00205_);
  and _43215_ (_00208_, _00204_, _35822_);
  not _43216_ (_00209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  nor _43217_ (_00210_, _00204_, _00209_);
  or _43218_ (_38489_, _00210_, _00208_);
  and _43219_ (_00211_, _00204_, _35826_);
  not _43220_ (_00212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  nor _43221_ (_00213_, _00204_, _00212_);
  or _43222_ (_38490_, _00213_, _00211_);
  and _43223_ (_00214_, _00204_, _35830_);
  not _43224_ (_00215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  nor _43225_ (_00216_, _00204_, _00215_);
  or _43226_ (_38491_, _00216_, _00214_);
  and _43227_ (_00217_, _00204_, _35834_);
  not _43228_ (_00218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  nor _43229_ (_00219_, _00204_, _00218_);
  or _43230_ (_38492_, _00219_, _00217_);
  and _43231_ (_00220_, _00204_, _35838_);
  not _43232_ (_00221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  nor _43233_ (_00222_, _00204_, _00221_);
  or _43234_ (_38493_, _00222_, _00220_);
  and _43235_ (_00223_, _00204_, _35842_);
  not _43236_ (_00224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  nor _43237_ (_00225_, _00204_, _00224_);
  or _43238_ (_38494_, _00225_, _00223_);
  and _43239_ (_00226_, _00204_, _35846_);
  not _43240_ (_00227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  nor _43241_ (_00228_, _00204_, _00227_);
  or _43242_ (_38495_, _00228_, _00226_);
  and _43243_ (_00229_, _36623_, _36141_);
  and _43244_ (_00230_, _00229_, _35815_);
  not _43245_ (_00231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  nor _43246_ (_00232_, _00229_, _00231_);
  or _43247_ (_38496_, _00232_, _00230_);
  and _43248_ (_00233_, _00229_, _35822_);
  not _43249_ (_00234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  nor _43250_ (_00235_, _00229_, _00234_);
  or _43251_ (_38497_, _00235_, _00233_);
  and _43252_ (_00236_, _00229_, _35826_);
  not _43253_ (_00237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  nor _43254_ (_00238_, _00229_, _00237_);
  or _43255_ (_38498_, _00238_, _00236_);
  and _43256_ (_00239_, _00229_, _35830_);
  not _43257_ (_00240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  nor _43258_ (_00241_, _00229_, _00240_);
  or _43259_ (_38499_, _00241_, _00239_);
  and _43260_ (_00242_, _00229_, _35834_);
  not _43261_ (_00243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  nor _43262_ (_00244_, _00229_, _00243_);
  or _43263_ (_38500_, _00244_, _00242_);
  and _43264_ (_00245_, _00229_, _35838_);
  not _43265_ (_00246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  nor _43266_ (_00247_, _00229_, _00246_);
  or _43267_ (_38501_, _00247_, _00245_);
  and _43268_ (_00248_, _00229_, _35842_);
  not _43269_ (_00249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  nor _43270_ (_00250_, _00229_, _00249_);
  or _43271_ (_38502_, _00250_, _00248_);
  and _43272_ (_00251_, _00229_, _35846_);
  not _43273_ (_00252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  nor _43274_ (_00253_, _00229_, _00252_);
  or _43275_ (_38503_, _00253_, _00251_);
  and _43276_ (_00254_, _36623_, _36167_);
  and _43277_ (_00255_, _00254_, _35815_);
  not _43278_ (_00256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  nor _43279_ (_00257_, _00254_, _00256_);
  or _43280_ (_38504_, _00257_, _00255_);
  and _43281_ (_00258_, _00254_, _35822_);
  not _43282_ (_00259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  nor _43283_ (_00260_, _00254_, _00259_);
  or _43284_ (_38505_, _00260_, _00258_);
  and _43285_ (_00261_, _00254_, _35826_);
  not _43286_ (_00262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  nor _43287_ (_00263_, _00254_, _00262_);
  or _43288_ (_38506_, _00263_, _00261_);
  and _43289_ (_00264_, _00254_, _35830_);
  not _43290_ (_00265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  nor _43291_ (_00266_, _00254_, _00265_);
  or _43292_ (_38507_, _00266_, _00264_);
  and _43293_ (_00267_, _00254_, _35834_);
  not _43294_ (_00268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  nor _43295_ (_00269_, _00254_, _00268_);
  or _43296_ (_38508_, _00269_, _00267_);
  and _43297_ (_00270_, _00254_, _35838_);
  not _43298_ (_00271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  nor _43299_ (_00272_, _00254_, _00271_);
  or _43300_ (_38509_, _00272_, _00270_);
  and _43301_ (_00273_, _00254_, _35842_);
  not _43302_ (_00274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  nor _43303_ (_00275_, _00254_, _00274_);
  or _43304_ (_38510_, _00275_, _00273_);
  and _43305_ (_00276_, _00254_, _35846_);
  not _43306_ (_00277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  nor _43307_ (_00278_, _00254_, _00277_);
  or _43308_ (_38511_, _00278_, _00276_);
  and _43309_ (_00279_, _36623_, _36193_);
  and _43310_ (_00280_, _00279_, _35815_);
  not _43311_ (_00281_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  nor _43312_ (_00282_, _00279_, _00281_);
  or _43313_ (_38512_, _00282_, _00280_);
  and _43314_ (_00283_, _00279_, _35822_);
  not _43315_ (_00284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  nor _43316_ (_00285_, _00279_, _00284_);
  or _43317_ (_38513_, _00285_, _00283_);
  and _43318_ (_00286_, _00279_, _35826_);
  not _43319_ (_00287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  nor _43320_ (_00288_, _00279_, _00287_);
  or _43321_ (_38514_, _00288_, _00286_);
  and _43322_ (_00289_, _00279_, _35830_);
  not _43323_ (_00290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  nor _43324_ (_00291_, _00279_, _00290_);
  or _43325_ (_38515_, _00291_, _00289_);
  and _43326_ (_00292_, _00279_, _35834_);
  not _43327_ (_00293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  nor _43328_ (_00294_, _00279_, _00293_);
  or _43329_ (_38516_, _00294_, _00292_);
  and _43330_ (_00295_, _00279_, _35838_);
  not _43331_ (_00296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  nor _43332_ (_00297_, _00279_, _00296_);
  or _43333_ (_38517_, _00297_, _00295_);
  and _43334_ (_00298_, _00279_, _35842_);
  not _43335_ (_00299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  nor _43336_ (_00300_, _00279_, _00299_);
  or _43337_ (_38518_, _00300_, _00298_);
  and _43338_ (_00301_, _00279_, _35846_);
  not _43339_ (_00302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  nor _43340_ (_00303_, _00279_, _00302_);
  or _43341_ (_38519_, _00303_, _00301_);
  and _43342_ (_00304_, _35573_, _34640_);
  and _43343_ (_00305_, _00304_, _36219_);
  and _43344_ (_00306_, _00305_, _35572_);
  and _43345_ (_00307_, _00306_, _35815_);
  not _43346_ (_00308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  nor _43347_ (_00309_, _00306_, _00308_);
  or _43348_ (_38520_, _00309_, _00307_);
  and _43349_ (_00310_, _00306_, _35822_);
  not _43350_ (_00311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  nor _43351_ (_00312_, _00306_, _00311_);
  or _43352_ (_38521_, _00312_, _00310_);
  and _43353_ (_00313_, _00306_, _35826_);
  not _43354_ (_00314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  nor _43355_ (_00315_, _00306_, _00314_);
  or _43356_ (_38522_, _00315_, _00313_);
  and _43357_ (_00316_, _00306_, _35830_);
  not _43358_ (_00317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  nor _43359_ (_00318_, _00306_, _00317_);
  or _43360_ (_38523_, _00318_, _00316_);
  and _43361_ (_00319_, _00306_, _35834_);
  not _43362_ (_00320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  nor _43363_ (_00321_, _00306_, _00320_);
  or _43364_ (_38524_, _00321_, _00319_);
  and _43365_ (_00322_, _00306_, _35838_);
  not _43366_ (_00323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  nor _43367_ (_00324_, _00306_, _00323_);
  or _43368_ (_38525_, _00324_, _00322_);
  and _43369_ (_00325_, _00306_, _35842_);
  not _43370_ (_00326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  nor _43371_ (_00327_, _00306_, _00326_);
  or _43372_ (_38526_, _00327_, _00325_);
  and _43373_ (_00328_, _00306_, _35846_);
  not _43374_ (_00329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  nor _43375_ (_00330_, _00306_, _00329_);
  or _43376_ (_38527_, _00330_, _00328_);
  and _43377_ (_00331_, _00305_, _35817_);
  and _43378_ (_00332_, _00331_, _35815_);
  not _43379_ (_00333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  nor _43380_ (_00334_, _00331_, _00333_);
  or _43381_ (_38528_, _00334_, _00332_);
  and _43382_ (_00335_, _00331_, _35822_);
  not _43383_ (_00336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  nor _43384_ (_00337_, _00331_, _00336_);
  or _43385_ (_38529_, _00337_, _00335_);
  and _43386_ (_00338_, _00331_, _35826_);
  not _43387_ (_00339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  nor _43388_ (_00340_, _00331_, _00339_);
  or _43389_ (_38530_, _00340_, _00338_);
  and _43390_ (_00341_, _00331_, _35830_);
  not _43391_ (_00342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  nor _43392_ (_00343_, _00331_, _00342_);
  or _43393_ (_38531_, _00343_, _00341_);
  and _43394_ (_00344_, _00331_, _35834_);
  not _43395_ (_00345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  nor _43396_ (_00346_, _00331_, _00345_);
  or _43397_ (_38532_, _00346_, _00344_);
  and _43398_ (_00347_, _00331_, _35838_);
  not _43399_ (_00348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  nor _43400_ (_00349_, _00331_, _00348_);
  or _43401_ (_38533_, _00349_, _00347_);
  and _43402_ (_00350_, _00331_, _35842_);
  not _43403_ (_00351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  nor _43404_ (_00352_, _00331_, _00351_);
  or _43405_ (_38534_, _00352_, _00350_);
  and _43406_ (_00353_, _00331_, _35846_);
  not _43407_ (_00354_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  nor _43408_ (_00355_, _00331_, _00354_);
  or _43409_ (_38535_, _00355_, _00353_);
  and _43410_ (_00356_, _00305_, _35851_);
  and _43411_ (_00357_, _00356_, _35815_);
  not _43412_ (_00358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  nor _43413_ (_00359_, _00356_, _00358_);
  or _43414_ (_38544_, _00359_, _00357_);
  and _43415_ (_00360_, _00356_, _35822_);
  not _43416_ (_00361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  nor _43417_ (_00362_, _00356_, _00361_);
  or _43418_ (_38545_, _00362_, _00360_);
  and _43419_ (_00363_, _00356_, _35826_);
  not _43420_ (_00364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  nor _43421_ (_00365_, _00356_, _00364_);
  or _43422_ (_38546_, _00365_, _00363_);
  and _43423_ (_00366_, _00356_, _35830_);
  not _43424_ (_00367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  nor _43425_ (_00368_, _00356_, _00367_);
  or _43426_ (_38547_, _00368_, _00366_);
  and _43427_ (_00369_, _00356_, _35834_);
  not _43428_ (_00370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  nor _43429_ (_00371_, _00356_, _00370_);
  or _43430_ (_38548_, _00371_, _00369_);
  and _43431_ (_00372_, _00356_, _35838_);
  not _43432_ (_00373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  nor _43433_ (_00374_, _00356_, _00373_);
  or _43434_ (_38549_, _00374_, _00372_);
  and _43435_ (_00375_, _00356_, _35842_);
  not _43436_ (_00376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  nor _43437_ (_00377_, _00356_, _00376_);
  or _43438_ (_38550_, _00377_, _00375_);
  and _43439_ (_00378_, _00356_, _35846_);
  not _43440_ (_00379_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  nor _43441_ (_00380_, _00356_, _00379_);
  or _43442_ (_38551_, _00380_, _00378_);
  and _43443_ (_00381_, _00305_, _35878_);
  and _43444_ (_00382_, _00381_, _35815_);
  not _43445_ (_00383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  nor _43446_ (_00384_, _00381_, _00383_);
  or _43447_ (_38552_, _00384_, _00382_);
  and _43448_ (_00385_, _00381_, _35822_);
  not _43449_ (_00386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  nor _43450_ (_00387_, _00381_, _00386_);
  or _43451_ (_38553_, _00387_, _00385_);
  and _43452_ (_00388_, _00381_, _35826_);
  not _43453_ (_00389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  nor _43454_ (_00390_, _00381_, _00389_);
  or _43455_ (_38554_, _00390_, _00388_);
  and _43456_ (_00391_, _00381_, _35830_);
  not _43457_ (_00392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  nor _43458_ (_00393_, _00381_, _00392_);
  or _43459_ (_38555_, _00393_, _00391_);
  and _43460_ (_00394_, _00381_, _35834_);
  not _43461_ (_00395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  nor _43462_ (_00396_, _00381_, _00395_);
  or _43463_ (_38556_, _00396_, _00394_);
  and _43464_ (_00397_, _00381_, _35838_);
  not _43465_ (_00398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  nor _43466_ (_00399_, _00381_, _00398_);
  or _43467_ (_38557_, _00399_, _00397_);
  and _43468_ (_00400_, _00381_, _35842_);
  not _43469_ (_00401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  nor _43470_ (_00402_, _00381_, _00401_);
  or _43471_ (_38558_, _00402_, _00400_);
  and _43472_ (_00403_, _00381_, _35846_);
  not _43473_ (_00404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  nor _43474_ (_00405_, _00381_, _00404_);
  or _43475_ (_38559_, _00405_, _00403_);
  and _43476_ (_00406_, _00305_, _35905_);
  and _43477_ (_00407_, _00406_, _35815_);
  not _43478_ (_00408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  nor _43479_ (_00409_, _00406_, _00408_);
  or _43480_ (_38560_, _00409_, _00407_);
  and _43481_ (_00410_, _00406_, _35822_);
  not _43482_ (_00411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  nor _43483_ (_00412_, _00406_, _00411_);
  or _43484_ (_38561_, _00412_, _00410_);
  and _43485_ (_00413_, _00406_, _35826_);
  not _43486_ (_00414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  nor _43487_ (_00415_, _00406_, _00414_);
  or _43488_ (_38562_, _00415_, _00413_);
  and _43489_ (_00416_, _00406_, _35830_);
  not _43490_ (_00417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  nor _43491_ (_00418_, _00406_, _00417_);
  or _43492_ (_38563_, _00418_, _00416_);
  and _43493_ (_00419_, _00406_, _35834_);
  not _43494_ (_00420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  nor _43495_ (_00421_, _00406_, _00420_);
  or _43496_ (_38564_, _00421_, _00419_);
  and _43497_ (_00422_, _00406_, _35838_);
  not _43498_ (_00423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  nor _43499_ (_00424_, _00406_, _00423_);
  or _43500_ (_38565_, _00424_, _00422_);
  and _43501_ (_00425_, _00406_, _35842_);
  not _43502_ (_00426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  nor _43503_ (_00427_, _00406_, _00426_);
  or _43504_ (_38566_, _00427_, _00425_);
  and _43505_ (_00428_, _00406_, _35846_);
  not _43506_ (_00429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  nor _43507_ (_00430_, _00406_, _00429_);
  or _43508_ (_38567_, _00430_, _00428_);
  and _43509_ (_00431_, _00305_, _35931_);
  and _43510_ (_00432_, _00431_, _35815_);
  not _43511_ (_00433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  nor _43512_ (_00434_, _00431_, _00433_);
  or _43513_ (_38568_, _00434_, _00432_);
  and _43514_ (_00435_, _00431_, _35822_);
  not _43515_ (_00436_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  nor _43516_ (_00437_, _00431_, _00436_);
  or _43517_ (_38569_, _00437_, _00435_);
  and _43518_ (_00438_, _00431_, _35826_);
  not _43519_ (_00439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  nor _43520_ (_00440_, _00431_, _00439_);
  or _43521_ (_38570_, _00440_, _00438_);
  and _43522_ (_00441_, _00431_, _35830_);
  not _43523_ (_00442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  nor _43524_ (_00443_, _00431_, _00442_);
  or _43525_ (_38571_, _00443_, _00441_);
  and _43526_ (_00444_, _00431_, _35834_);
  not _43527_ (_00445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  nor _43528_ (_00446_, _00431_, _00445_);
  or _43529_ (_38572_, _00446_, _00444_);
  and _43530_ (_00447_, _00431_, _35838_);
  not _43531_ (_00448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  nor _43532_ (_00449_, _00431_, _00448_);
  or _43533_ (_38573_, _00449_, _00447_);
  and _43534_ (_00450_, _00431_, _35842_);
  not _43535_ (_00451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  nor _43536_ (_00452_, _00431_, _00451_);
  or _43537_ (_38574_, _00452_, _00450_);
  and _43538_ (_00453_, _00431_, _35846_);
  not _43539_ (_00454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  nor _43540_ (_00455_, _00431_, _00454_);
  or _43541_ (_38575_, _00455_, _00453_);
  and _43542_ (_00456_, _00305_, _35957_);
  and _43543_ (_00457_, _00456_, _35815_);
  not _43544_ (_00458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  nor _43545_ (_00459_, _00456_, _00458_);
  or _43546_ (_38576_, _00459_, _00457_);
  and _43547_ (_00460_, _00456_, _35822_);
  not _43548_ (_00461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  nor _43549_ (_00462_, _00456_, _00461_);
  or _43550_ (_38577_, _00462_, _00460_);
  and _43551_ (_00463_, _00456_, _35826_);
  not _43552_ (_00464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  nor _43553_ (_00465_, _00456_, _00464_);
  or _43554_ (_38578_, _00465_, _00463_);
  and _43555_ (_00466_, _00456_, _35830_);
  not _43556_ (_00467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  nor _43557_ (_00468_, _00456_, _00467_);
  or _43558_ (_38579_, _00468_, _00466_);
  and _43559_ (_00469_, _00456_, _35834_);
  not _43560_ (_00470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  nor _43561_ (_00471_, _00456_, _00470_);
  or _43562_ (_38580_, _00471_, _00469_);
  and _43563_ (_00472_, _00456_, _35838_);
  not _43564_ (_00473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  nor _43565_ (_00474_, _00456_, _00473_);
  or _43566_ (_38581_, _00474_, _00472_);
  and _43567_ (_00475_, _00456_, _35842_);
  not _43568_ (_00476_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  nor _43569_ (_00477_, _00456_, _00476_);
  or _43570_ (_38582_, _00477_, _00475_);
  and _43571_ (_00478_, _00456_, _35846_);
  not _43572_ (_00479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  nor _43573_ (_00480_, _00456_, _00479_);
  or _43574_ (_38583_, _00480_, _00478_);
  and _43575_ (_00481_, _00305_, _35983_);
  and _43576_ (_00482_, _00481_, _35815_);
  not _43577_ (_00483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  nor _43578_ (_00484_, _00481_, _00483_);
  or _43579_ (_38584_, _00484_, _00482_);
  and _43580_ (_00485_, _00481_, _35822_);
  not _43581_ (_00486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  nor _43582_ (_00487_, _00481_, _00486_);
  or _43583_ (_38585_, _00487_, _00485_);
  and _43584_ (_00488_, _00481_, _35826_);
  not _43585_ (_00489_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  nor _43586_ (_00490_, _00481_, _00489_);
  or _43587_ (_38586_, _00490_, _00488_);
  and _43588_ (_00491_, _00481_, _35830_);
  not _43589_ (_00492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  nor _43590_ (_00493_, _00481_, _00492_);
  or _43591_ (_38587_, _00493_, _00491_);
  and _43592_ (_00494_, _00481_, _35834_);
  not _43593_ (_00495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  nor _43594_ (_00496_, _00481_, _00495_);
  or _43595_ (_38588_, _00496_, _00494_);
  and _43596_ (_00497_, _00481_, _35838_);
  not _43597_ (_00498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  nor _43598_ (_00499_, _00481_, _00498_);
  or _43599_ (_38589_, _00499_, _00497_);
  and _43600_ (_00500_, _00481_, _35842_);
  not _43601_ (_00501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  nor _43602_ (_00502_, _00481_, _00501_);
  or _43603_ (_38590_, _00502_, _00500_);
  and _43604_ (_00503_, _00481_, _35846_);
  not _43605_ (_00504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  nor _43606_ (_00505_, _00481_, _00504_);
  or _43607_ (_38591_, _00505_, _00503_);
  and _43608_ (_00506_, _00305_, _36010_);
  and _43609_ (_00507_, _00506_, _35815_);
  not _43610_ (_00508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  nor _43611_ (_00509_, _00506_, _00508_);
  or _43612_ (_38592_, _00509_, _00507_);
  and _43613_ (_00510_, _00506_, _35822_);
  not _43614_ (_00511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  nor _43615_ (_00512_, _00506_, _00511_);
  or _43616_ (_38593_, _00512_, _00510_);
  and _43617_ (_00513_, _00506_, _35826_);
  not _43618_ (_00514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  nor _43619_ (_00515_, _00506_, _00514_);
  or _43620_ (_38594_, _00515_, _00513_);
  and _43621_ (_00516_, _00506_, _35830_);
  not _43622_ (_00517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  nor _43623_ (_00518_, _00506_, _00517_);
  or _43624_ (_38595_, _00518_, _00516_);
  and _43625_ (_00519_, _00506_, _35834_);
  not _43626_ (_00520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  nor _43627_ (_00521_, _00506_, _00520_);
  or _43628_ (_38596_, _00521_, _00519_);
  and _43629_ (_00522_, _00506_, _35838_);
  not _43630_ (_00523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  nor _43631_ (_00524_, _00506_, _00523_);
  or _43632_ (_38597_, _00524_, _00522_);
  and _43633_ (_00525_, _00506_, _35842_);
  not _43634_ (_00526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  nor _43635_ (_00527_, _00506_, _00526_);
  or _43636_ (_38598_, _00527_, _00525_);
  and _43637_ (_00528_, _00506_, _35846_);
  not _43638_ (_00529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  nor _43639_ (_00530_, _00506_, _00529_);
  or _43640_ (_38599_, _00530_, _00528_);
  and _43641_ (_00531_, _00305_, _36036_);
  and _43642_ (_00532_, _00531_, _35815_);
  not _43643_ (_00533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  nor _43644_ (_00534_, _00531_, _00533_);
  or _43645_ (_38600_, _00534_, _00532_);
  and _43646_ (_00535_, _00531_, _35822_);
  not _43647_ (_00536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  nor _43648_ (_00537_, _00531_, _00536_);
  or _43649_ (_38601_, _00537_, _00535_);
  and _43650_ (_00538_, _00531_, _35826_);
  not _43651_ (_00539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  nor _43652_ (_00540_, _00531_, _00539_);
  or _43653_ (_38602_, _00540_, _00538_);
  and _43654_ (_00541_, _00531_, _35830_);
  not _43655_ (_00542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  nor _43656_ (_00543_, _00531_, _00542_);
  or _43657_ (_38603_, _00543_, _00541_);
  and _43658_ (_00544_, _00531_, _35834_);
  not _43659_ (_00545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  nor _43660_ (_00546_, _00531_, _00545_);
  or _43661_ (_38604_, _00546_, _00544_);
  and _43662_ (_00547_, _00531_, _35838_);
  not _43663_ (_00548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  nor _43664_ (_00549_, _00531_, _00548_);
  or _43665_ (_38605_, _00549_, _00547_);
  and _43666_ (_00550_, _00531_, _35842_);
  not _43667_ (_00551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  nor _43668_ (_00552_, _00531_, _00551_);
  or _43669_ (_38606_, _00552_, _00550_);
  and _43670_ (_00553_, _00531_, _35846_);
  not _43671_ (_00554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  nor _43672_ (_00555_, _00531_, _00554_);
  or _43673_ (_38607_, _00555_, _00553_);
  and _43674_ (_00556_, _00305_, _36062_);
  and _43675_ (_00557_, _00556_, _35815_);
  not _43676_ (_00558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  nor _43677_ (_00559_, _00556_, _00558_);
  or _43678_ (_38608_, _00559_, _00557_);
  and _43679_ (_00560_, _00556_, _35822_);
  not _43680_ (_00561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  nor _43681_ (_00562_, _00556_, _00561_);
  or _43682_ (_38609_, _00562_, _00560_);
  and _43683_ (_00563_, _00556_, _35826_);
  not _43684_ (_00564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  nor _43685_ (_00565_, _00556_, _00564_);
  or _43686_ (_38610_, _00565_, _00563_);
  and _43687_ (_00566_, _00556_, _35830_);
  not _43688_ (_00567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  nor _43689_ (_00568_, _00556_, _00567_);
  or _43690_ (_38611_, _00568_, _00566_);
  and _43691_ (_00569_, _00556_, _35834_);
  not _43692_ (_00570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  nor _43693_ (_00571_, _00556_, _00570_);
  or _43694_ (_38612_, _00571_, _00569_);
  and _43695_ (_00572_, _00556_, _35838_);
  not _43696_ (_00573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  nor _43697_ (_00574_, _00556_, _00573_);
  or _43698_ (_38613_, _00574_, _00572_);
  and _43699_ (_00575_, _00556_, _35842_);
  not _43700_ (_00576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  nor _43701_ (_00577_, _00556_, _00576_);
  or _43702_ (_38614_, _00577_, _00575_);
  and _43703_ (_00578_, _00556_, _35846_);
  not _43704_ (_00579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  nor _43705_ (_00580_, _00556_, _00579_);
  or _43706_ (_38615_, _00580_, _00578_);
  and _43707_ (_00581_, _00305_, _36088_);
  and _43708_ (_00582_, _00581_, _35815_);
  not _43709_ (_00583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  nor _43710_ (_00584_, _00581_, _00583_);
  or _43711_ (_38616_, _00584_, _00582_);
  and _43712_ (_00585_, _00581_, _35822_);
  not _43713_ (_00586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  nor _43714_ (_00587_, _00581_, _00586_);
  or _43715_ (_38617_, _00587_, _00585_);
  and _43716_ (_00588_, _00581_, _35826_);
  not _43717_ (_00589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  nor _43718_ (_00590_, _00581_, _00589_);
  or _43719_ (_38618_, _00590_, _00588_);
  and _43720_ (_00591_, _00581_, _35830_);
  not _43721_ (_00592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  nor _43722_ (_00593_, _00581_, _00592_);
  or _43723_ (_38619_, _00593_, _00591_);
  and _43724_ (_00594_, _00581_, _35834_);
  not _43725_ (_00595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  nor _43726_ (_00596_, _00581_, _00595_);
  or _43727_ (_38620_, _00596_, _00594_);
  and _43728_ (_00597_, _00581_, _35838_);
  not _43729_ (_00598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  nor _43730_ (_00599_, _00581_, _00598_);
  or _43731_ (_38621_, _00599_, _00597_);
  and _43732_ (_00600_, _00581_, _35842_);
  not _43733_ (_00601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  nor _43734_ (_00602_, _00581_, _00601_);
  or _43735_ (_38622_, _00602_, _00600_);
  and _43736_ (_00603_, _00581_, _35846_);
  not _43737_ (_00604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  nor _43738_ (_00605_, _00581_, _00604_);
  or _43739_ (_38623_, _00605_, _00603_);
  and _43740_ (_00606_, _00305_, _36115_);
  and _43741_ (_00607_, _00606_, _35815_);
  not _43742_ (_00608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  nor _43743_ (_00609_, _00606_, _00608_);
  or _43744_ (_38632_, _00609_, _00607_);
  and _43745_ (_00610_, _00606_, _35822_);
  not _43746_ (_00611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  nor _43747_ (_00612_, _00606_, _00611_);
  or _43748_ (_38633_, _00612_, _00610_);
  and _43749_ (_00613_, _00606_, _35826_);
  not _43750_ (_00614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  nor _43751_ (_00615_, _00606_, _00614_);
  or _43752_ (_38634_, _00615_, _00613_);
  and _43753_ (_00616_, _00606_, _35830_);
  not _43754_ (_00617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  nor _43755_ (_00618_, _00606_, _00617_);
  or _43756_ (_38635_, _00618_, _00616_);
  and _43757_ (_00619_, _00606_, _35834_);
  not _43758_ (_00620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  nor _43759_ (_00621_, _00606_, _00620_);
  or _43760_ (_38636_, _00621_, _00619_);
  and _43761_ (_00622_, _00606_, _35838_);
  not _43762_ (_00623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  nor _43763_ (_00624_, _00606_, _00623_);
  or _43764_ (_38637_, _00624_, _00622_);
  and _43765_ (_00625_, _00606_, _35842_);
  not _43766_ (_00626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  nor _43767_ (_00627_, _00606_, _00626_);
  or _43768_ (_38638_, _00627_, _00625_);
  and _43769_ (_00628_, _00606_, _35846_);
  not _43770_ (_00629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  nor _43771_ (_00630_, _00606_, _00629_);
  or _43772_ (_38639_, _00630_, _00628_);
  and _43773_ (_00631_, _00305_, _36141_);
  and _43774_ (_00632_, _00631_, _35815_);
  not _43775_ (_00633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  nor _43776_ (_00634_, _00631_, _00633_);
  or _43777_ (_38640_, _00634_, _00632_);
  and _43778_ (_00635_, _00631_, _35822_);
  not _43779_ (_00636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  nor _43780_ (_00637_, _00631_, _00636_);
  or _43781_ (_38641_, _00637_, _00635_);
  and _43782_ (_00638_, _00631_, _35826_);
  not _43783_ (_00639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  nor _43784_ (_00640_, _00631_, _00639_);
  or _43785_ (_38642_, _00640_, _00638_);
  and _43786_ (_00641_, _00631_, _35830_);
  not _43787_ (_00642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  nor _43788_ (_00643_, _00631_, _00642_);
  or _43789_ (_38643_, _00643_, _00641_);
  and _43790_ (_00644_, _00631_, _35834_);
  not _43791_ (_00645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  nor _43792_ (_00646_, _00631_, _00645_);
  or _43793_ (_38644_, _00646_, _00644_);
  and _43794_ (_00647_, _00631_, _35838_);
  not _43795_ (_00648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  nor _43796_ (_00649_, _00631_, _00648_);
  or _43797_ (_38645_, _00649_, _00647_);
  and _43798_ (_00650_, _00631_, _35842_);
  not _43799_ (_00651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  nor _43800_ (_00652_, _00631_, _00651_);
  or _43801_ (_38646_, _00652_, _00650_);
  and _43802_ (_00653_, _00631_, _35846_);
  not _43803_ (_00654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  nor _43804_ (_00655_, _00631_, _00654_);
  or _43805_ (_38647_, _00655_, _00653_);
  and _43806_ (_00656_, _00305_, _36167_);
  and _43807_ (_00657_, _00656_, _35815_);
  not _43808_ (_00658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  nor _43809_ (_00659_, _00656_, _00658_);
  or _43810_ (_38648_, _00659_, _00657_);
  and _43811_ (_00660_, _00656_, _35822_);
  not _43812_ (_00661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  nor _43813_ (_00662_, _00656_, _00661_);
  or _43814_ (_38649_, _00662_, _00660_);
  and _43815_ (_00663_, _00656_, _35826_);
  not _43816_ (_00664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  nor _43817_ (_00665_, _00656_, _00664_);
  or _43818_ (_38650_, _00665_, _00663_);
  and _43819_ (_00666_, _00656_, _35830_);
  not _43820_ (_00667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  nor _43821_ (_00668_, _00656_, _00667_);
  or _43822_ (_38651_, _00668_, _00666_);
  and _43823_ (_00669_, _00656_, _35834_);
  not _43824_ (_00670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  nor _43825_ (_00671_, _00656_, _00670_);
  or _43826_ (_38652_, _00671_, _00669_);
  and _43827_ (_00672_, _00656_, _35838_);
  not _43828_ (_00673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  nor _43829_ (_00674_, _00656_, _00673_);
  or _43830_ (_38653_, _00674_, _00672_);
  and _43831_ (_00675_, _00656_, _35842_);
  not _43832_ (_00676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  nor _43833_ (_00677_, _00656_, _00676_);
  or _43834_ (_38654_, _00677_, _00675_);
  and _43835_ (_00678_, _00656_, _35846_);
  not _43836_ (_00679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  nor _43837_ (_00680_, _00656_, _00679_);
  or _43838_ (_38655_, _00680_, _00678_);
  and _43839_ (_00681_, _00305_, _36193_);
  and _43840_ (_00682_, _00681_, _35815_);
  not _43841_ (_00683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  nor _43842_ (_00684_, _00681_, _00683_);
  or _43843_ (_38656_, _00684_, _00682_);
  and _43844_ (_00685_, _00681_, _35822_);
  not _43845_ (_00686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  nor _43846_ (_00687_, _00681_, _00686_);
  or _43847_ (_38657_, _00687_, _00685_);
  and _43848_ (_00688_, _00681_, _35826_);
  not _43849_ (_00689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  nor _43850_ (_00690_, _00681_, _00689_);
  or _43851_ (_38658_, _00690_, _00688_);
  and _43852_ (_00691_, _00681_, _35830_);
  not _43853_ (_00692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  nor _43854_ (_00693_, _00681_, _00692_);
  or _43855_ (_38659_, _00693_, _00691_);
  and _43856_ (_00694_, _00681_, _35834_);
  not _43857_ (_00695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  nor _43858_ (_00696_, _00681_, _00695_);
  or _43859_ (_38660_, _00696_, _00694_);
  and _43860_ (_00697_, _00681_, _35838_);
  not _43861_ (_00698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  nor _43862_ (_00699_, _00681_, _00698_);
  or _43863_ (_38661_, _00699_, _00697_);
  and _43864_ (_00700_, _00681_, _35842_);
  not _43865_ (_00701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  nor _43866_ (_00702_, _00681_, _00701_);
  or _43867_ (_38662_, _00702_, _00700_);
  and _43868_ (_00703_, _00681_, _35846_);
  not _43869_ (_00704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  nor _43870_ (_00705_, _00681_, _00704_);
  or _43871_ (_38663_, _00705_, _00703_);
  and _43872_ (_00706_, _33659_, _33618_);
  and _43873_ (_00707_, _00706_, _34693_);
  and _43874_ (_00708_, _00707_, _35575_);
  and _43875_ (_00709_, _00708_, _35572_);
  and _43876_ (_00710_, _00709_, _35815_);
  not _43877_ (_00711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  nor _43878_ (_00712_, _00709_, _00711_);
  or _43879_ (_38664_, _00712_, _00710_);
  and _43880_ (_00713_, _00709_, _35822_);
  not _43881_ (_00714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  nor _43882_ (_00715_, _00709_, _00714_);
  or _43883_ (_38665_, _00715_, _00713_);
  and _43884_ (_00716_, _00709_, _35826_);
  not _43885_ (_00717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  nor _43886_ (_00718_, _00709_, _00717_);
  or _43887_ (_38666_, _00718_, _00716_);
  and _43888_ (_00719_, _00709_, _35830_);
  not _43889_ (_00720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  nor _43890_ (_00721_, _00709_, _00720_);
  or _43891_ (_38667_, _00721_, _00719_);
  and _43892_ (_00722_, _00709_, _35834_);
  not _43893_ (_00723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  nor _43894_ (_00724_, _00709_, _00723_);
  or _43895_ (_38668_, _00724_, _00722_);
  and _43896_ (_00725_, _00709_, _35838_);
  not _43897_ (_00726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  nor _43898_ (_00727_, _00709_, _00726_);
  or _43899_ (_38669_, _00727_, _00725_);
  and _43900_ (_00728_, _00709_, _35842_);
  not _43901_ (_00729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  nor _43902_ (_00730_, _00709_, _00729_);
  or _43903_ (_38670_, _00730_, _00728_);
  and _43904_ (_00731_, _00709_, _35846_);
  not _43905_ (_00732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  nor _43906_ (_00733_, _00709_, _00732_);
  or _43907_ (_38671_, _00733_, _00731_);
  and _43908_ (_00734_, _00708_, _35817_);
  and _43909_ (_00735_, _00734_, _35815_);
  not _43910_ (_00736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  nor _43911_ (_00737_, _00734_, _00736_);
  or _43912_ (_38672_, _00737_, _00735_);
  and _43913_ (_00738_, _00734_, _35822_);
  not _43914_ (_00739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  nor _43915_ (_00740_, _00734_, _00739_);
  or _43916_ (_38673_, _00740_, _00738_);
  and _43917_ (_00741_, _00734_, _35826_);
  not _43918_ (_00742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  nor _43919_ (_00743_, _00734_, _00742_);
  or _43920_ (_38674_, _00743_, _00741_);
  and _43921_ (_00744_, _00734_, _35830_);
  not _43922_ (_00745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  nor _43923_ (_00746_, _00734_, _00745_);
  or _43924_ (_38675_, _00746_, _00744_);
  and _43925_ (_00747_, _00734_, _35834_);
  not _43926_ (_00748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  nor _43927_ (_00749_, _00734_, _00748_);
  or _43928_ (_38676_, _00749_, _00747_);
  and _43929_ (_00750_, _00734_, _35838_);
  not _43930_ (_00751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  nor _43931_ (_00752_, _00734_, _00751_);
  or _43932_ (_38677_, _00752_, _00750_);
  and _43933_ (_00753_, _00734_, _35842_);
  not _43934_ (_00754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  nor _43935_ (_00755_, _00734_, _00754_);
  or _43936_ (_38678_, _00755_, _00753_);
  and _43937_ (_00756_, _00734_, _35846_);
  not _43938_ (_00757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  nor _43939_ (_00758_, _00734_, _00757_);
  or _43940_ (_38679_, _00758_, _00756_);
  and _43941_ (_00759_, _00708_, _35851_);
  and _43942_ (_00760_, _00759_, _35815_);
  not _43943_ (_00761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  nor _43944_ (_00762_, _00759_, _00761_);
  or _43945_ (_38680_, _00762_, _00760_);
  and _43946_ (_00763_, _00759_, _35822_);
  not _43947_ (_00764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  nor _43948_ (_00765_, _00759_, _00764_);
  or _43949_ (_38681_, _00765_, _00763_);
  and _43950_ (_00766_, _00759_, _35826_);
  not _43951_ (_00767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  nor _43952_ (_00768_, _00759_, _00767_);
  or _43953_ (_38682_, _00768_, _00766_);
  and _43954_ (_00769_, _00759_, _35830_);
  not _43955_ (_00770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  nor _43956_ (_00771_, _00759_, _00770_);
  or _43957_ (_38683_, _00771_, _00769_);
  and _43958_ (_00772_, _00759_, _35834_);
  not _43959_ (_00773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  nor _43960_ (_00774_, _00759_, _00773_);
  or _43961_ (_38684_, _00774_, _00772_);
  and _43962_ (_00775_, _00759_, _35838_);
  not _43963_ (_00776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  nor _43964_ (_00777_, _00759_, _00776_);
  or _43965_ (_38685_, _00777_, _00775_);
  and _43966_ (_00778_, _00759_, _35842_);
  not _43967_ (_00779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  nor _43968_ (_00780_, _00759_, _00779_);
  or _43969_ (_38686_, _00780_, _00778_);
  and _43970_ (_00781_, _00759_, _35846_);
  not _43971_ (_00782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  nor _43972_ (_00783_, _00759_, _00782_);
  or _43973_ (_38687_, _00783_, _00781_);
  and _43974_ (_00784_, _00708_, _35878_);
  and _43975_ (_00785_, _00784_, _35815_);
  not _43976_ (_00786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  nor _43977_ (_00787_, _00784_, _00786_);
  or _43978_ (_38688_, _00787_, _00785_);
  and _43979_ (_00788_, _00784_, _35822_);
  not _43980_ (_00789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  nor _43981_ (_00790_, _00784_, _00789_);
  or _43982_ (_38689_, _00790_, _00788_);
  and _43983_ (_00791_, _00784_, _35826_);
  not _43984_ (_00792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  nor _43985_ (_00793_, _00784_, _00792_);
  or _43986_ (_38690_, _00793_, _00791_);
  and _43987_ (_00794_, _00784_, _35830_);
  not _43988_ (_00795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  nor _43989_ (_00796_, _00784_, _00795_);
  or _43990_ (_38691_, _00796_, _00794_);
  and _43991_ (_00797_, _00784_, _35834_);
  not _43992_ (_00798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  nor _43993_ (_00799_, _00784_, _00798_);
  or _43994_ (_38692_, _00799_, _00797_);
  and _43995_ (_00800_, _00784_, _35838_);
  not _43996_ (_00801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  nor _43997_ (_00802_, _00784_, _00801_);
  or _43998_ (_38693_, _00802_, _00800_);
  and _43999_ (_00803_, _00784_, _35842_);
  not _44000_ (_00804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  nor _44001_ (_00805_, _00784_, _00804_);
  or _44002_ (_38694_, _00805_, _00803_);
  and _44003_ (_00806_, _00784_, _35846_);
  not _44004_ (_00807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  nor _44005_ (_00808_, _00784_, _00807_);
  or _44006_ (_38695_, _00808_, _00806_);
  and _44007_ (_00809_, _00708_, _35905_);
  and _44008_ (_00810_, _00809_, _35815_);
  not _44009_ (_00811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  nor _44010_ (_00812_, _00809_, _00811_);
  or _44011_ (_38696_, _00812_, _00810_);
  and _44012_ (_00813_, _00809_, _35822_);
  not _44013_ (_00814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  nor _44014_ (_00815_, _00809_, _00814_);
  or _44015_ (_38697_, _00815_, _00813_);
  and _44016_ (_00816_, _00809_, _35826_);
  not _44017_ (_00817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  nor _44018_ (_00818_, _00809_, _00817_);
  or _44019_ (_38698_, _00818_, _00816_);
  and _44020_ (_00819_, _00809_, _35830_);
  not _44021_ (_00820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  nor _44022_ (_00821_, _00809_, _00820_);
  or _44023_ (_38699_, _00821_, _00819_);
  and _44024_ (_00822_, _00809_, _35834_);
  not _44025_ (_00823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  nor _44026_ (_00824_, _00809_, _00823_);
  or _44027_ (_38700_, _00824_, _00822_);
  and _44028_ (_00825_, _00809_, _35838_);
  not _44029_ (_00826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  nor _44030_ (_00827_, _00809_, _00826_);
  or _44031_ (_38701_, _00827_, _00825_);
  and _44032_ (_00828_, _00809_, _35842_);
  not _44033_ (_00829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  nor _44034_ (_00830_, _00809_, _00829_);
  or _44035_ (_38702_, _00830_, _00828_);
  and _44036_ (_00831_, _00809_, _35846_);
  not _44037_ (_00832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  nor _44038_ (_00833_, _00809_, _00832_);
  or _44039_ (_38703_, _00833_, _00831_);
  and _44040_ (_00834_, _00708_, _35931_);
  and _44041_ (_00835_, _00834_, _35815_);
  not _44042_ (_00836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  nor _44043_ (_00837_, _00834_, _00836_);
  or _44044_ (_38704_, _00837_, _00835_);
  and _44045_ (_00838_, _00834_, _35822_);
  not _44046_ (_00839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  nor _44047_ (_00840_, _00834_, _00839_);
  or _44048_ (_38705_, _00840_, _00838_);
  and _44049_ (_00841_, _00834_, _35826_);
  not _44050_ (_00842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  nor _44051_ (_00843_, _00834_, _00842_);
  or _44052_ (_38706_, _00843_, _00841_);
  and _44053_ (_00844_, _00834_, _35830_);
  not _44054_ (_00845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  nor _44055_ (_00846_, _00834_, _00845_);
  or _44056_ (_38707_, _00846_, _00844_);
  and _44057_ (_00847_, _00834_, _35834_);
  not _44058_ (_00848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  nor _44059_ (_00849_, _00834_, _00848_);
  or _44060_ (_38708_, _00849_, _00847_);
  and _44061_ (_00850_, _00834_, _35838_);
  not _44062_ (_00851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  nor _44063_ (_00852_, _00834_, _00851_);
  or _44064_ (_38709_, _00852_, _00850_);
  and _44065_ (_00853_, _00834_, _35842_);
  not _44066_ (_00854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  nor _44067_ (_00855_, _00834_, _00854_);
  or _44068_ (_38710_, _00855_, _00853_);
  and _44069_ (_00856_, _00834_, _35846_);
  not _44070_ (_00857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  nor _44071_ (_00858_, _00834_, _00857_);
  or _44072_ (_38711_, _00858_, _00856_);
  and _44073_ (_00859_, _00708_, _35957_);
  and _44074_ (_00860_, _00859_, _35815_);
  not _44075_ (_00861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  nor _44076_ (_00862_, _00859_, _00861_);
  or _44077_ (_38720_, _00862_, _00860_);
  and _44078_ (_00863_, _00859_, _35822_);
  not _44079_ (_00864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  nor _44080_ (_00865_, _00859_, _00864_);
  or _44081_ (_38721_, _00865_, _00863_);
  and _44082_ (_00866_, _00859_, _35826_);
  not _44083_ (_00867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  nor _44084_ (_00868_, _00859_, _00867_);
  or _44085_ (_38722_, _00868_, _00866_);
  and _44086_ (_00869_, _00859_, _35830_);
  not _44087_ (_00870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  nor _44088_ (_00871_, _00859_, _00870_);
  or _44089_ (_38723_, _00871_, _00869_);
  and _44090_ (_00872_, _00859_, _35834_);
  not _44091_ (_00873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  nor _44092_ (_00874_, _00859_, _00873_);
  or _44093_ (_38724_, _00874_, _00872_);
  and _44094_ (_00875_, _00859_, _35838_);
  not _44095_ (_00876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  nor _44096_ (_00877_, _00859_, _00876_);
  or _44097_ (_38725_, _00877_, _00875_);
  and _44098_ (_00878_, _00859_, _35842_);
  not _44099_ (_00879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  nor _44100_ (_00880_, _00859_, _00879_);
  or _44101_ (_38726_, _00880_, _00878_);
  and _44102_ (_00881_, _00859_, _35846_);
  not _44103_ (_00882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  nor _44104_ (_00883_, _00859_, _00882_);
  or _44105_ (_38727_, _00883_, _00881_);
  and _44106_ (_00884_, _00708_, _35983_);
  and _44107_ (_00885_, _00884_, _35815_);
  not _44108_ (_00886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  nor _44109_ (_00887_, _00884_, _00886_);
  or _44110_ (_38728_, _00887_, _00885_);
  and _44111_ (_00888_, _00884_, _35822_);
  not _44112_ (_00889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  nor _44113_ (_00890_, _00884_, _00889_);
  or _44114_ (_38729_, _00890_, _00888_);
  and _44115_ (_00891_, _00884_, _35826_);
  not _44116_ (_00892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  nor _44117_ (_00893_, _00884_, _00892_);
  or _44118_ (_38730_, _00893_, _00891_);
  and _44119_ (_00894_, _00884_, _35830_);
  not _44120_ (_00895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  nor _44121_ (_00896_, _00884_, _00895_);
  or _44122_ (_38731_, _00896_, _00894_);
  and _44123_ (_00897_, _00884_, _35834_);
  not _44124_ (_00898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  nor _44125_ (_00899_, _00884_, _00898_);
  or _44126_ (_38732_, _00899_, _00897_);
  and _44127_ (_00900_, _00884_, _35838_);
  not _44128_ (_00901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  nor _44129_ (_00902_, _00884_, _00901_);
  or _44130_ (_38733_, _00902_, _00900_);
  and _44131_ (_00903_, _00884_, _35842_);
  not _44132_ (_00904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  nor _44133_ (_00905_, _00884_, _00904_);
  or _44134_ (_38734_, _00905_, _00903_);
  and _44135_ (_00906_, _00884_, _35846_);
  not _44136_ (_00907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  nor _44137_ (_00908_, _00884_, _00907_);
  or _44138_ (_38735_, _00908_, _00906_);
  and _44139_ (_00909_, _00708_, _36010_);
  and _44140_ (_00910_, _00909_, _35815_);
  not _44141_ (_00911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  nor _44142_ (_00912_, _00909_, _00911_);
  or _44143_ (_38736_, _00912_, _00910_);
  and _44144_ (_00913_, _00909_, _35822_);
  not _44145_ (_00914_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  nor _44146_ (_00915_, _00909_, _00914_);
  or _44147_ (_38737_, _00915_, _00913_);
  and _44148_ (_00916_, _00909_, _35826_);
  not _44149_ (_00917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  nor _44150_ (_00918_, _00909_, _00917_);
  or _44151_ (_38738_, _00918_, _00916_);
  and _44152_ (_00919_, _00909_, _35830_);
  not _44153_ (_00920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  nor _44154_ (_00921_, _00909_, _00920_);
  or _44155_ (_38739_, _00921_, _00919_);
  and _44156_ (_00922_, _00909_, _35834_);
  not _44157_ (_00923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  nor _44158_ (_00924_, _00909_, _00923_);
  or _44159_ (_38740_, _00924_, _00922_);
  and _44160_ (_00925_, _00909_, _35838_);
  not _44161_ (_00926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  nor _44162_ (_00927_, _00909_, _00926_);
  or _44163_ (_38741_, _00927_, _00925_);
  and _44164_ (_00928_, _00909_, _35842_);
  not _44165_ (_00929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  nor _44166_ (_00930_, _00909_, _00929_);
  or _44167_ (_38742_, _00930_, _00928_);
  and _44168_ (_00931_, _00909_, _35846_);
  not _44169_ (_00932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  nor _44170_ (_00933_, _00909_, _00932_);
  or _44171_ (_38743_, _00933_, _00931_);
  and _44172_ (_00934_, _00708_, _36036_);
  and _44173_ (_00935_, _00934_, _35815_);
  not _44174_ (_00936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  nor _44175_ (_00937_, _00934_, _00936_);
  or _44176_ (_38744_, _00937_, _00935_);
  and _44177_ (_00938_, _00934_, _35822_);
  not _44178_ (_00939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  nor _44179_ (_00940_, _00934_, _00939_);
  or _44180_ (_38745_, _00940_, _00938_);
  and _44181_ (_00941_, _00934_, _35826_);
  not _44182_ (_00942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  nor _44183_ (_00943_, _00934_, _00942_);
  or _44184_ (_38746_, _00943_, _00941_);
  and _44185_ (_00944_, _00934_, _35830_);
  not _44186_ (_00945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  nor _44187_ (_00946_, _00934_, _00945_);
  or _44188_ (_38747_, _00946_, _00944_);
  and _44189_ (_00947_, _00934_, _35834_);
  not _44190_ (_00948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  nor _44191_ (_00949_, _00934_, _00948_);
  or _44192_ (_38748_, _00949_, _00947_);
  and _44193_ (_00950_, _00934_, _35838_);
  not _44194_ (_00951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  nor _44195_ (_00952_, _00934_, _00951_);
  or _44196_ (_38749_, _00952_, _00950_);
  and _44197_ (_00953_, _00934_, _35842_);
  not _44198_ (_00954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  nor _44199_ (_00955_, _00934_, _00954_);
  or _44200_ (_38750_, _00955_, _00953_);
  and _44201_ (_00956_, _00934_, _35846_);
  not _44202_ (_00957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  nor _44203_ (_00958_, _00934_, _00957_);
  or _44204_ (_38751_, _00958_, _00956_);
  and _44205_ (_00959_, _00708_, _36062_);
  and _44206_ (_00960_, _00959_, _35815_);
  not _44207_ (_00961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  nor _44208_ (_00962_, _00959_, _00961_);
  or _44209_ (_38752_, _00962_, _00960_);
  and _44210_ (_00963_, _00959_, _35822_);
  not _44211_ (_00964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  nor _44212_ (_00965_, _00959_, _00964_);
  or _44213_ (_38753_, _00965_, _00963_);
  and _44214_ (_00966_, _00959_, _35826_);
  not _44215_ (_00967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  nor _44216_ (_00968_, _00959_, _00967_);
  or _44217_ (_38754_, _00968_, _00966_);
  and _44218_ (_00969_, _00959_, _35830_);
  not _44219_ (_00970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  nor _44220_ (_00971_, _00959_, _00970_);
  or _44221_ (_38755_, _00971_, _00969_);
  and _44222_ (_00972_, _00959_, _35834_);
  not _44223_ (_00973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  nor _44224_ (_00974_, _00959_, _00973_);
  or _44225_ (_38756_, _00974_, _00972_);
  and _44226_ (_00975_, _00959_, _35838_);
  not _44227_ (_00976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  nor _44228_ (_00977_, _00959_, _00976_);
  or _44229_ (_38757_, _00977_, _00975_);
  and _44230_ (_00978_, _00959_, _35842_);
  not _44231_ (_00979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  nor _44232_ (_00980_, _00959_, _00979_);
  or _44233_ (_38758_, _00980_, _00978_);
  and _44234_ (_00981_, _00959_, _35846_);
  not _44235_ (_00982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  nor _44236_ (_00983_, _00959_, _00982_);
  or _44237_ (_38759_, _00983_, _00981_);
  and _44238_ (_00984_, _00708_, _36088_);
  and _44239_ (_00985_, _00984_, _35815_);
  not _44240_ (_00986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  nor _44241_ (_00987_, _00984_, _00986_);
  or _44242_ (_38760_, _00987_, _00985_);
  and _44243_ (_00988_, _00984_, _35822_);
  not _44244_ (_00989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  nor _44245_ (_00990_, _00984_, _00989_);
  or _44246_ (_38761_, _00990_, _00988_);
  and _44247_ (_00991_, _00984_, _35826_);
  not _44248_ (_00992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  nor _44249_ (_00993_, _00984_, _00992_);
  or _44250_ (_38762_, _00993_, _00991_);
  and _44251_ (_00994_, _00984_, _35830_);
  not _44252_ (_00995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  nor _44253_ (_00996_, _00984_, _00995_);
  or _44254_ (_38763_, _00996_, _00994_);
  and _44255_ (_00997_, _00984_, _35834_);
  not _44256_ (_00998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  nor _44257_ (_00999_, _00984_, _00998_);
  or _44258_ (_38764_, _00999_, _00997_);
  and _44259_ (_01000_, _00984_, _35838_);
  not _44260_ (_01001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  nor _44261_ (_01002_, _00984_, _01001_);
  or _44262_ (_38765_, _01002_, _01000_);
  and _44263_ (_01003_, _00984_, _35842_);
  not _44264_ (_01004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  nor _44265_ (_01005_, _00984_, _01004_);
  or _44266_ (_38766_, _01005_, _01003_);
  and _44267_ (_01006_, _00984_, _35846_);
  not _44268_ (_01007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  nor _44269_ (_01008_, _00984_, _01007_);
  or _44270_ (_38767_, _01008_, _01006_);
  and _44271_ (_01009_, _00708_, _36115_);
  and _44272_ (_01010_, _01009_, _35815_);
  not _44273_ (_01011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  nor _44274_ (_01012_, _01009_, _01011_);
  or _44275_ (_38768_, _01012_, _01010_);
  and _44276_ (_01013_, _01009_, _35822_);
  not _44277_ (_01014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  nor _44278_ (_01015_, _01009_, _01014_);
  or _44279_ (_38769_, _01015_, _01013_);
  and _44280_ (_01016_, _01009_, _35826_);
  not _44281_ (_01017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  nor _44282_ (_01018_, _01009_, _01017_);
  or _44283_ (_38770_, _01018_, _01016_);
  and _44284_ (_01019_, _01009_, _35830_);
  not _44285_ (_01020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  nor _44286_ (_01021_, _01009_, _01020_);
  or _44287_ (_38771_, _01021_, _01019_);
  and _44288_ (_01022_, _01009_, _35834_);
  not _44289_ (_01023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  nor _44290_ (_01024_, _01009_, _01023_);
  or _44291_ (_38772_, _01024_, _01022_);
  and _44292_ (_01025_, _01009_, _35838_);
  not _44293_ (_01026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  nor _44294_ (_01027_, _01009_, _01026_);
  or _44295_ (_38773_, _01027_, _01025_);
  and _44296_ (_01028_, _01009_, _35842_);
  not _44297_ (_01029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  nor _44298_ (_01030_, _01009_, _01029_);
  or _44299_ (_38774_, _01030_, _01028_);
  and _44300_ (_01031_, _01009_, _35846_);
  not _44301_ (_01032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  nor _44302_ (_01033_, _01009_, _01032_);
  or _44303_ (_38775_, _01033_, _01031_);
  and _44304_ (_01034_, _00708_, _36141_);
  and _44305_ (_01035_, _01034_, _35815_);
  not _44306_ (_01036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  nor _44307_ (_01037_, _01034_, _01036_);
  or _44308_ (_38776_, _01037_, _01035_);
  and _44309_ (_01038_, _01034_, _35822_);
  not _44310_ (_01039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  nor _44311_ (_01040_, _01034_, _01039_);
  or _44312_ (_38777_, _01040_, _01038_);
  and _44313_ (_01041_, _01034_, _35826_);
  not _44314_ (_01042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  nor _44315_ (_01043_, _01034_, _01042_);
  or _44316_ (_38778_, _01043_, _01041_);
  and _44317_ (_01044_, _01034_, _35830_);
  not _44318_ (_01045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  nor _44319_ (_01046_, _01034_, _01045_);
  or _44320_ (_38779_, _01046_, _01044_);
  and _44321_ (_01047_, _01034_, _35834_);
  not _44322_ (_01048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  nor _44323_ (_01049_, _01034_, _01048_);
  or _44324_ (_38780_, _01049_, _01047_);
  and _44325_ (_01050_, _01034_, _35838_);
  not _44326_ (_01051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  nor _44327_ (_01052_, _01034_, _01051_);
  or _44328_ (_38781_, _01052_, _01050_);
  and _44329_ (_01053_, _01034_, _35842_);
  not _44330_ (_01054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  nor _44331_ (_01055_, _01034_, _01054_);
  or _44332_ (_38782_, _01055_, _01053_);
  and _44333_ (_01056_, _01034_, _35846_);
  not _44334_ (_01057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  nor _44335_ (_01058_, _01034_, _01057_);
  or _44336_ (_38783_, _01058_, _01056_);
  and _44337_ (_01059_, _00708_, _36167_);
  and _44338_ (_01060_, _01059_, _35815_);
  not _44339_ (_01061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  nor _44340_ (_01062_, _01059_, _01061_);
  or _44341_ (_38784_, _01062_, _01060_);
  and _44342_ (_01063_, _01059_, _35822_);
  not _44343_ (_01064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  nor _44344_ (_01065_, _01059_, _01064_);
  or _44345_ (_38785_, _01065_, _01063_);
  and _44346_ (_01066_, _01059_, _35826_);
  not _44347_ (_01067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  nor _44348_ (_01068_, _01059_, _01067_);
  or _44349_ (_38786_, _01068_, _01066_);
  and _44350_ (_01069_, _01059_, _35830_);
  not _44351_ (_01070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  nor _44352_ (_01071_, _01059_, _01070_);
  or _44353_ (_38787_, _01071_, _01069_);
  and _44354_ (_01072_, _01059_, _35834_);
  not _44355_ (_01073_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  nor _44356_ (_01074_, _01059_, _01073_);
  or _44357_ (_38788_, _01074_, _01072_);
  and _44358_ (_01075_, _01059_, _35838_);
  not _44359_ (_01076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  nor _44360_ (_01077_, _01059_, _01076_);
  or _44361_ (_38789_, _01077_, _01075_);
  and _44362_ (_01078_, _01059_, _35842_);
  not _44363_ (_01079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  nor _44364_ (_01080_, _01059_, _01079_);
  or _44365_ (_38790_, _01080_, _01078_);
  and _44366_ (_01081_, _01059_, _35846_);
  not _44367_ (_01082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  nor _44368_ (_01083_, _01059_, _01082_);
  or _44369_ (_38791_, _01083_, _01081_);
  and _44370_ (_01084_, _00708_, _36193_);
  and _44371_ (_01085_, _01084_, _35815_);
  not _44372_ (_01086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  nor _44373_ (_01087_, _01084_, _01086_);
  or _44374_ (_38792_, _01087_, _01085_);
  and _44375_ (_01088_, _01084_, _35822_);
  not _44376_ (_01089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  nor _44377_ (_01090_, _01084_, _01089_);
  or _44378_ (_38793_, _01090_, _01088_);
  and _44379_ (_01091_, _01084_, _35826_);
  not _44380_ (_01092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  nor _44381_ (_01093_, _01084_, _01092_);
  or _44382_ (_38794_, _01093_, _01091_);
  and _44383_ (_01094_, _01084_, _35830_);
  not _44384_ (_01095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  nor _44385_ (_01096_, _01084_, _01095_);
  or _44386_ (_38795_, _01096_, _01094_);
  and _44387_ (_01097_, _01084_, _35834_);
  not _44388_ (_01098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  nor _44389_ (_01099_, _01084_, _01098_);
  or _44390_ (_38796_, _01099_, _01097_);
  and _44391_ (_01100_, _01084_, _35838_);
  not _44392_ (_01101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  nor _44393_ (_01102_, _01084_, _01101_);
  or _44394_ (_38797_, _01102_, _01100_);
  and _44395_ (_01103_, _01084_, _35842_);
  not _44396_ (_01104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  nor _44397_ (_01105_, _01084_, _01104_);
  or _44398_ (_38798_, _01105_, _01103_);
  and _44399_ (_01106_, _01084_, _35846_);
  not _44400_ (_01107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  nor _44401_ (_01108_, _01084_, _01107_);
  or _44402_ (_38799_, _01108_, _01106_);
  and _44403_ (_01109_, _00707_, _36220_);
  and _44404_ (_01110_, _01109_, _35572_);
  and _44405_ (_01111_, _01110_, _35815_);
  not _44406_ (_01112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  nor _44407_ (_01113_, _01110_, _01112_);
  or _44408_ (_38808_, _01113_, _01111_);
  and _44409_ (_01114_, _01110_, _35822_);
  not _44410_ (_01115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  nor _44411_ (_01116_, _01110_, _01115_);
  or _44412_ (_38809_, _01116_, _01114_);
  and _44413_ (_01117_, _01110_, _35826_);
  not _44414_ (_01118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  nor _44415_ (_01119_, _01110_, _01118_);
  or _44416_ (_38810_, _01119_, _01117_);
  and _44417_ (_01120_, _01110_, _35830_);
  not _44418_ (_01121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  nor _44419_ (_01122_, _01110_, _01121_);
  or _44420_ (_38811_, _01122_, _01120_);
  and _44421_ (_01123_, _01110_, _35834_);
  not _44422_ (_01124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  nor _44423_ (_01125_, _01110_, _01124_);
  or _44424_ (_38812_, _01125_, _01123_);
  and _44425_ (_01126_, _01110_, _35838_);
  not _44426_ (_01127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  nor _44427_ (_01128_, _01110_, _01127_);
  or _44428_ (_38813_, _01128_, _01126_);
  and _44429_ (_01129_, _01110_, _35842_);
  not _44430_ (_01130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  nor _44431_ (_01131_, _01110_, _01130_);
  or _44432_ (_38814_, _01131_, _01129_);
  and _44433_ (_01132_, _01110_, _35846_);
  not _44434_ (_01133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  nor _44435_ (_01134_, _01110_, _01133_);
  or _44436_ (_38815_, _01134_, _01132_);
  and _44437_ (_01135_, _01109_, _35817_);
  and _44438_ (_01136_, _01135_, _35815_);
  not _44439_ (_01137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  nor _44440_ (_01138_, _01135_, _01137_);
  or _44441_ (_38816_, _01138_, _01136_);
  and _44442_ (_01139_, _01135_, _35822_);
  not _44443_ (_01140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  nor _44444_ (_01141_, _01135_, _01140_);
  or _44445_ (_38817_, _01141_, _01139_);
  and _44446_ (_01142_, _01135_, _35826_);
  not _44447_ (_01143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  nor _44448_ (_01144_, _01135_, _01143_);
  or _44449_ (_38818_, _01144_, _01142_);
  and _44450_ (_01145_, _01135_, _35830_);
  not _44451_ (_01146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  nor _44452_ (_01147_, _01135_, _01146_);
  or _44453_ (_38819_, _01147_, _01145_);
  and _44454_ (_01148_, _01135_, _35834_);
  not _44455_ (_01149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  nor _44456_ (_01150_, _01135_, _01149_);
  or _44457_ (_38820_, _01150_, _01148_);
  and _44458_ (_01151_, _01135_, _35838_);
  not _44459_ (_01152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  nor _44460_ (_01153_, _01135_, _01152_);
  or _44461_ (_38821_, _01153_, _01151_);
  and _44462_ (_01154_, _01135_, _35842_);
  not _44463_ (_01155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  nor _44464_ (_01156_, _01135_, _01155_);
  or _44465_ (_38822_, _01156_, _01154_);
  and _44466_ (_01157_, _01135_, _35846_);
  not _44467_ (_01158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  nor _44468_ (_01159_, _01135_, _01158_);
  or _44469_ (_38823_, _01159_, _01157_);
  and _44470_ (_01160_, _01109_, _35851_);
  and _44471_ (_01161_, _01160_, _35815_);
  not _44472_ (_01162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  nor _44473_ (_01163_, _01160_, _01162_);
  or _44474_ (_38824_, _01163_, _01161_);
  and _44475_ (_01164_, _01160_, _35822_);
  not _44476_ (_01165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  nor _44477_ (_01166_, _01160_, _01165_);
  or _44478_ (_38825_, _01166_, _01164_);
  and _44479_ (_01167_, _01160_, _35826_);
  not _44480_ (_01168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  nor _44481_ (_01169_, _01160_, _01168_);
  or _44482_ (_38826_, _01169_, _01167_);
  and _44483_ (_01170_, _01160_, _35830_);
  not _44484_ (_01171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  nor _44485_ (_01172_, _01160_, _01171_);
  or _44486_ (_38827_, _01172_, _01170_);
  and _44487_ (_01173_, _01160_, _35834_);
  not _44488_ (_01174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  nor _44489_ (_01175_, _01160_, _01174_);
  or _44490_ (_38828_, _01175_, _01173_);
  and _44491_ (_01176_, _01160_, _35838_);
  not _44492_ (_01177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  nor _44493_ (_01178_, _01160_, _01177_);
  or _44494_ (_38829_, _01178_, _01176_);
  and _44495_ (_01179_, _01160_, _35842_);
  not _44496_ (_01180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  nor _44497_ (_01181_, _01160_, _01180_);
  or _44498_ (_38830_, _01181_, _01179_);
  and _44499_ (_01182_, _01160_, _35846_);
  not _44500_ (_01183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  nor _44501_ (_01184_, _01160_, _01183_);
  or _44502_ (_38831_, _01184_, _01182_);
  and _44503_ (_01185_, _01109_, _35878_);
  and _44504_ (_01186_, _01185_, _35815_);
  not _44505_ (_01187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  nor _44506_ (_01188_, _01185_, _01187_);
  or _44507_ (_38832_, _01188_, _01186_);
  and _44508_ (_01189_, _01185_, _35822_);
  not _44509_ (_01190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  nor _44510_ (_01191_, _01185_, _01190_);
  or _44511_ (_38833_, _01191_, _01189_);
  and _44512_ (_01192_, _01185_, _35826_);
  not _44513_ (_01193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  nor _44514_ (_01194_, _01185_, _01193_);
  or _44515_ (_38834_, _01194_, _01192_);
  and _44516_ (_01195_, _01185_, _35830_);
  not _44517_ (_01196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  nor _44518_ (_01197_, _01185_, _01196_);
  or _44519_ (_38835_, _01197_, _01195_);
  and _44520_ (_01198_, _01185_, _35834_);
  not _44521_ (_01199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  nor _44522_ (_01200_, _01185_, _01199_);
  or _44523_ (_38836_, _01200_, _01198_);
  and _44524_ (_01201_, _01185_, _35838_);
  not _44525_ (_01202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  nor _44526_ (_01203_, _01185_, _01202_);
  or _44527_ (_38837_, _01203_, _01201_);
  and _44528_ (_01204_, _01185_, _35842_);
  not _44529_ (_01205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  nor _44530_ (_01206_, _01185_, _01205_);
  or _44531_ (_38838_, _01206_, _01204_);
  and _44532_ (_01207_, _01185_, _35846_);
  not _44533_ (_01208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  nor _44534_ (_01209_, _01185_, _01208_);
  or _44535_ (_38839_, _01209_, _01207_);
  and _44536_ (_01210_, _01109_, _35905_);
  and _44537_ (_01211_, _01210_, _35815_);
  not _44538_ (_01212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  nor _44539_ (_01213_, _01210_, _01212_);
  or _44540_ (_38840_, _01213_, _01211_);
  and _44541_ (_01214_, _01210_, _35822_);
  not _44542_ (_01215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  nor _44543_ (_01216_, _01210_, _01215_);
  or _44544_ (_38841_, _01216_, _01214_);
  and _44545_ (_01217_, _01210_, _35826_);
  not _44546_ (_01218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  nor _44547_ (_01219_, _01210_, _01218_);
  or _44548_ (_38842_, _01219_, _01217_);
  and _44549_ (_01220_, _01210_, _35830_);
  not _44550_ (_01221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  nor _44551_ (_01222_, _01210_, _01221_);
  or _44552_ (_38843_, _01222_, _01220_);
  and _44553_ (_01223_, _01210_, _35834_);
  not _44554_ (_01224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  nor _44555_ (_01225_, _01210_, _01224_);
  or _44556_ (_38844_, _01225_, _01223_);
  and _44557_ (_01226_, _01210_, _35838_);
  not _44558_ (_01227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  nor _44559_ (_01228_, _01210_, _01227_);
  or _44560_ (_38845_, _01228_, _01226_);
  and _44561_ (_01229_, _01210_, _35842_);
  not _44562_ (_01230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  nor _44563_ (_01231_, _01210_, _01230_);
  or _44564_ (_38846_, _01231_, _01229_);
  and _44565_ (_01232_, _01210_, _35846_);
  not _44566_ (_01233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  nor _44567_ (_01234_, _01210_, _01233_);
  or _44568_ (_38847_, _01234_, _01232_);
  and _44569_ (_01235_, _01109_, _35931_);
  and _44570_ (_01236_, _01235_, _35815_);
  not _44571_ (_01237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  nor _44572_ (_01238_, _01235_, _01237_);
  or _44573_ (_38848_, _01238_, _01236_);
  and _44574_ (_01239_, _01235_, _35822_);
  not _44575_ (_01240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  nor _44576_ (_01241_, _01235_, _01240_);
  or _44577_ (_38849_, _01241_, _01239_);
  and _44578_ (_01242_, _01235_, _35826_);
  not _44579_ (_01243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  nor _44580_ (_01244_, _01235_, _01243_);
  or _44581_ (_38850_, _01244_, _01242_);
  and _44582_ (_01245_, _01235_, _35830_);
  not _44583_ (_01246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  nor _44584_ (_01247_, _01235_, _01246_);
  or _44585_ (_38851_, _01247_, _01245_);
  and _44586_ (_01248_, _01235_, _35834_);
  not _44587_ (_01249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  nor _44588_ (_01250_, _01235_, _01249_);
  or _44589_ (_38852_, _01250_, _01248_);
  and _44590_ (_01251_, _01235_, _35838_);
  not _44591_ (_01252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  nor _44592_ (_01253_, _01235_, _01252_);
  or _44593_ (_38853_, _01253_, _01251_);
  and _44594_ (_01254_, _01235_, _35842_);
  not _44595_ (_01255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  nor _44596_ (_01256_, _01235_, _01255_);
  or _44597_ (_38854_, _01256_, _01254_);
  and _44598_ (_01257_, _01235_, _35846_);
  not _44599_ (_01258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  nor _44600_ (_01259_, _01235_, _01258_);
  or _44601_ (_38855_, _01259_, _01257_);
  and _44602_ (_01260_, _01109_, _35957_);
  and _44603_ (_01261_, _01260_, _35815_);
  not _44604_ (_01262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  nor _44605_ (_01263_, _01260_, _01262_);
  or _44606_ (_38856_, _01263_, _01261_);
  and _44607_ (_01264_, _01260_, _35822_);
  not _44608_ (_01265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  nor _44609_ (_01266_, _01260_, _01265_);
  or _44610_ (_38857_, _01266_, _01264_);
  and _44611_ (_01267_, _01260_, _35826_);
  not _44612_ (_01268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  nor _44613_ (_01269_, _01260_, _01268_);
  or _44614_ (_38858_, _01269_, _01267_);
  and _44615_ (_01270_, _01260_, _35830_);
  not _44616_ (_01271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  nor _44617_ (_01272_, _01260_, _01271_);
  or _44618_ (_38859_, _01272_, _01270_);
  and _44619_ (_01273_, _01260_, _35834_);
  not _44620_ (_01274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  nor _44621_ (_01275_, _01260_, _01274_);
  or _44622_ (_38860_, _01275_, _01273_);
  and _44623_ (_01276_, _01260_, _35838_);
  not _44624_ (_01277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  nor _44625_ (_01278_, _01260_, _01277_);
  or _44626_ (_38861_, _01278_, _01276_);
  and _44627_ (_01279_, _01260_, _35842_);
  not _44628_ (_01280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  nor _44629_ (_01281_, _01260_, _01280_);
  or _44630_ (_38862_, _01281_, _01279_);
  and _44631_ (_01282_, _01260_, _35846_);
  not _44632_ (_01283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  nor _44633_ (_01284_, _01260_, _01283_);
  or _44634_ (_38863_, _01284_, _01282_);
  and _44635_ (_01285_, _01109_, _35983_);
  and _44636_ (_01286_, _01285_, _35815_);
  not _44637_ (_01287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  nor _44638_ (_01288_, _01285_, _01287_);
  or _44639_ (_38864_, _01288_, _01286_);
  and _44640_ (_01289_, _01285_, _35822_);
  not _44641_ (_01290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  nor _44642_ (_01291_, _01285_, _01290_);
  or _44643_ (_38865_, _01291_, _01289_);
  and _44644_ (_01292_, _01285_, _35826_);
  not _44645_ (_01293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  nor _44646_ (_01294_, _01285_, _01293_);
  or _44647_ (_38866_, _01294_, _01292_);
  and _44648_ (_01295_, _01285_, _35830_);
  not _44649_ (_01296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  nor _44650_ (_01297_, _01285_, _01296_);
  or _44651_ (_38867_, _01297_, _01295_);
  and _44652_ (_01298_, _01285_, _35834_);
  not _44653_ (_01299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  nor _44654_ (_01300_, _01285_, _01299_);
  or _44655_ (_38868_, _01300_, _01298_);
  and _44656_ (_01301_, _01285_, _35838_);
  not _44657_ (_01302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  nor _44658_ (_01303_, _01285_, _01302_);
  or _44659_ (_38869_, _01303_, _01301_);
  and _44660_ (_01304_, _01285_, _35842_);
  not _44661_ (_01305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  nor _44662_ (_01306_, _01285_, _01305_);
  or _44663_ (_38870_, _01306_, _01304_);
  and _44664_ (_01307_, _01285_, _35846_);
  not _44665_ (_01308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  nor _44666_ (_01309_, _01285_, _01308_);
  or _44667_ (_38871_, _01309_, _01307_);
  and _44668_ (_01310_, _01109_, _36010_);
  and _44669_ (_01311_, _01310_, _35815_);
  not _44670_ (_01312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  nor _44671_ (_01313_, _01310_, _01312_);
  or _44672_ (_38872_, _01313_, _01311_);
  and _44673_ (_01314_, _01310_, _35822_);
  not _44674_ (_01315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  nor _44675_ (_01316_, _01310_, _01315_);
  or _44676_ (_38873_, _01316_, _01314_);
  and _44677_ (_01317_, _01310_, _35826_);
  not _44678_ (_01318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  nor _44679_ (_01319_, _01310_, _01318_);
  or _44680_ (_38874_, _01319_, _01317_);
  and _44681_ (_01320_, _01310_, _35830_);
  not _44682_ (_01321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  nor _44683_ (_01322_, _01310_, _01321_);
  or _44684_ (_38875_, _01322_, _01320_);
  and _44685_ (_01323_, _01310_, _35834_);
  not _44686_ (_01324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  nor _44687_ (_01325_, _01310_, _01324_);
  or _44688_ (_38876_, _01325_, _01323_);
  and _44689_ (_01326_, _01310_, _35838_);
  not _44690_ (_01327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  nor _44691_ (_01328_, _01310_, _01327_);
  or _44692_ (_38877_, _01328_, _01326_);
  and _44693_ (_01329_, _01310_, _35842_);
  not _44694_ (_01330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  nor _44695_ (_01331_, _01310_, _01330_);
  or _44696_ (_38878_, _01331_, _01329_);
  and _44697_ (_01332_, _01310_, _35846_);
  not _44698_ (_01333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  nor _44699_ (_01334_, _01310_, _01333_);
  or _44700_ (_38879_, _01334_, _01332_);
  and _44701_ (_01335_, _01109_, _36036_);
  and _44702_ (_01336_, _01335_, _35815_);
  not _44703_ (_01337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  nor _44704_ (_01338_, _01335_, _01337_);
  or _44705_ (_38880_, _01338_, _01336_);
  and _44706_ (_01339_, _01335_, _35822_);
  not _44707_ (_01340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  nor _44708_ (_01341_, _01335_, _01340_);
  or _44709_ (_38881_, _01341_, _01339_);
  and _44710_ (_01342_, _01335_, _35826_);
  not _44711_ (_01343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  nor _44712_ (_01344_, _01335_, _01343_);
  or _44713_ (_38882_, _01344_, _01342_);
  and _44714_ (_01345_, _01335_, _35830_);
  not _44715_ (_01346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  nor _44716_ (_01347_, _01335_, _01346_);
  or _44717_ (_38883_, _01347_, _01345_);
  and _44718_ (_01348_, _01335_, _35834_);
  not _44719_ (_01349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  nor _44720_ (_01350_, _01335_, _01349_);
  or _44721_ (_38884_, _01350_, _01348_);
  and _44722_ (_01351_, _01335_, _35838_);
  not _44723_ (_01352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  nor _44724_ (_01353_, _01335_, _01352_);
  or _44725_ (_38885_, _01353_, _01351_);
  and _44726_ (_01354_, _01335_, _35842_);
  not _44727_ (_01355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  nor _44728_ (_01356_, _01335_, _01355_);
  or _44729_ (_38886_, _01356_, _01354_);
  and _44730_ (_01357_, _01335_, _35846_);
  not _44731_ (_01358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  nor _44732_ (_01359_, _01335_, _01358_);
  or _44733_ (_38887_, _01359_, _01357_);
  and _44734_ (_01360_, _01109_, _36062_);
  and _44735_ (_01361_, _01360_, _35815_);
  not _44736_ (_01362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  nor _44737_ (_01363_, _01360_, _01362_);
  or _44738_ (_38896_, _01363_, _01361_);
  and _44739_ (_01364_, _01360_, _35822_);
  not _44740_ (_01365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  nor _44741_ (_01366_, _01360_, _01365_);
  or _44742_ (_38897_, _01366_, _01364_);
  and _44743_ (_01367_, _01360_, _35826_);
  not _44744_ (_01368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  nor _44745_ (_01369_, _01360_, _01368_);
  or _44746_ (_38898_, _01369_, _01367_);
  and _44747_ (_01370_, _01360_, _35830_);
  not _44748_ (_01371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  nor _44749_ (_01372_, _01360_, _01371_);
  or _44750_ (_38899_, _01372_, _01370_);
  and _44751_ (_01373_, _01360_, _35834_);
  not _44752_ (_01374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  nor _44753_ (_01375_, _01360_, _01374_);
  or _44754_ (_38900_, _01375_, _01373_);
  and _44755_ (_01376_, _01360_, _35838_);
  not _44756_ (_01377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  nor _44757_ (_01378_, _01360_, _01377_);
  or _44758_ (_38901_, _01378_, _01376_);
  and _44759_ (_01379_, _01360_, _35842_);
  not _44760_ (_01380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  nor _44761_ (_01381_, _01360_, _01380_);
  or _44762_ (_38902_, _01381_, _01379_);
  and _44763_ (_01382_, _01360_, _35846_);
  not _44764_ (_01383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  nor _44765_ (_01384_, _01360_, _01383_);
  or _44766_ (_38903_, _01384_, _01382_);
  and _44767_ (_01385_, _01109_, _36088_);
  and _44768_ (_01386_, _01385_, _35815_);
  not _44769_ (_01387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  nor _44770_ (_01388_, _01385_, _01387_);
  or _44771_ (_38904_, _01388_, _01386_);
  and _44772_ (_01389_, _01385_, _35822_);
  not _44773_ (_01390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  nor _44774_ (_01391_, _01385_, _01390_);
  or _44775_ (_38905_, _01391_, _01389_);
  and _44776_ (_01392_, _01385_, _35826_);
  not _44777_ (_01393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  nor _44778_ (_01394_, _01385_, _01393_);
  or _44779_ (_38906_, _01394_, _01392_);
  and _44780_ (_01395_, _01385_, _35830_);
  not _44781_ (_01396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  nor _44782_ (_01397_, _01385_, _01396_);
  or _44783_ (_38907_, _01397_, _01395_);
  and _44784_ (_01398_, _01385_, _35834_);
  not _44785_ (_01399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  nor _44786_ (_01400_, _01385_, _01399_);
  or _44787_ (_38908_, _01400_, _01398_);
  and _44788_ (_01401_, _01385_, _35838_);
  not _44789_ (_01402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  nor _44790_ (_01403_, _01385_, _01402_);
  or _44791_ (_38909_, _01403_, _01401_);
  and _44792_ (_01404_, _01385_, _35842_);
  not _44793_ (_01405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  nor _44794_ (_01406_, _01385_, _01405_);
  or _44795_ (_38910_, _01406_, _01404_);
  and _44796_ (_01407_, _01385_, _35846_);
  not _44797_ (_01408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  nor _44798_ (_01409_, _01385_, _01408_);
  or _44799_ (_38911_, _01409_, _01407_);
  and _44800_ (_01410_, _01109_, _36115_);
  and _44801_ (_01411_, _01410_, _35815_);
  not _44802_ (_01412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  nor _44803_ (_01413_, _01410_, _01412_);
  or _44804_ (_38912_, _01413_, _01411_);
  and _44805_ (_01414_, _01410_, _35822_);
  not _44806_ (_01415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  nor _44807_ (_01416_, _01410_, _01415_);
  or _44808_ (_38913_, _01416_, _01414_);
  and _44809_ (_01417_, _01410_, _35826_);
  not _44810_ (_01418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  nor _44811_ (_01419_, _01410_, _01418_);
  or _44812_ (_38914_, _01419_, _01417_);
  and _44813_ (_01420_, _01410_, _35830_);
  not _44814_ (_01421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  nor _44815_ (_01422_, _01410_, _01421_);
  or _44816_ (_38915_, _01422_, _01420_);
  and _44817_ (_01423_, _01410_, _35834_);
  not _44818_ (_01424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  nor _44819_ (_01425_, _01410_, _01424_);
  or _44820_ (_38916_, _01425_, _01423_);
  and _44821_ (_01426_, _01410_, _35838_);
  not _44822_ (_01427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  nor _44823_ (_01428_, _01410_, _01427_);
  or _44824_ (_38917_, _01428_, _01426_);
  and _44825_ (_01429_, _01410_, _35842_);
  not _44826_ (_01430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  nor _44827_ (_01431_, _01410_, _01430_);
  or _44828_ (_38918_, _01431_, _01429_);
  and _44829_ (_01432_, _01410_, _35846_);
  not _44830_ (_01433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  nor _44831_ (_01434_, _01410_, _01433_);
  or _44832_ (_38919_, _01434_, _01432_);
  and _44833_ (_01435_, _01109_, _36141_);
  and _44834_ (_01436_, _01435_, _35815_);
  not _44835_ (_01437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  nor _44836_ (_01438_, _01435_, _01437_);
  or _44837_ (_38920_, _01438_, _01436_);
  and _44838_ (_01439_, _01435_, _35822_);
  not _44839_ (_01440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  nor _44840_ (_01441_, _01435_, _01440_);
  or _44841_ (_38921_, _01441_, _01439_);
  and _44842_ (_01442_, _01435_, _35826_);
  not _44843_ (_01443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  nor _44844_ (_01444_, _01435_, _01443_);
  or _44845_ (_38922_, _01444_, _01442_);
  and _44846_ (_01445_, _01435_, _35830_);
  not _44847_ (_01446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  nor _44848_ (_01447_, _01435_, _01446_);
  or _44849_ (_38923_, _01447_, _01445_);
  and _44850_ (_01448_, _01435_, _35834_);
  not _44851_ (_01449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  nor _44852_ (_01450_, _01435_, _01449_);
  or _44853_ (_38924_, _01450_, _01448_);
  and _44854_ (_01451_, _01435_, _35838_);
  not _44855_ (_01452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  nor _44856_ (_01453_, _01435_, _01452_);
  or _44857_ (_38925_, _01453_, _01451_);
  and _44858_ (_01454_, _01435_, _35842_);
  not _44859_ (_01455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  nor _44860_ (_01456_, _01435_, _01455_);
  or _44861_ (_38926_, _01456_, _01454_);
  and _44862_ (_01457_, _01435_, _35846_);
  not _44863_ (_01458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  nor _44864_ (_01459_, _01435_, _01458_);
  or _44865_ (_38927_, _01459_, _01457_);
  and _44866_ (_01460_, _01109_, _36167_);
  and _44867_ (_01461_, _01460_, _35815_);
  not _44868_ (_01462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  nor _44869_ (_01463_, _01460_, _01462_);
  or _44870_ (_38928_, _01463_, _01461_);
  and _44871_ (_01464_, _01460_, _35822_);
  not _44872_ (_01465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  nor _44873_ (_01466_, _01460_, _01465_);
  or _44874_ (_38929_, _01466_, _01464_);
  and _44875_ (_01467_, _01460_, _35826_);
  not _44876_ (_01468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  nor _44877_ (_01469_, _01460_, _01468_);
  or _44878_ (_38930_, _01469_, _01467_);
  and _44879_ (_01470_, _01460_, _35830_);
  not _44880_ (_01471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  nor _44881_ (_01472_, _01460_, _01471_);
  or _44882_ (_38931_, _01472_, _01470_);
  and _44883_ (_01473_, _01460_, _35834_);
  not _44884_ (_01474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  nor _44885_ (_01475_, _01460_, _01474_);
  or _44886_ (_38932_, _01475_, _01473_);
  and _44887_ (_01476_, _01460_, _35838_);
  not _44888_ (_01477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  nor _44889_ (_01478_, _01460_, _01477_);
  or _44890_ (_38933_, _01478_, _01476_);
  and _44891_ (_01479_, _01460_, _35842_);
  not _44892_ (_01480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  nor _44893_ (_01481_, _01460_, _01480_);
  or _44894_ (_38934_, _01481_, _01479_);
  and _44895_ (_01482_, _01460_, _35846_);
  not _44896_ (_01483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  nor _44897_ (_01484_, _01460_, _01483_);
  or _44898_ (_38935_, _01484_, _01482_);
  and _44899_ (_01485_, _01109_, _36193_);
  and _44900_ (_01486_, _01485_, _35815_);
  not _44901_ (_01487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  nor _44902_ (_01488_, _01485_, _01487_);
  or _44903_ (_38936_, _01488_, _01486_);
  and _44904_ (_01489_, _01485_, _35822_);
  not _44905_ (_01490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  nor _44906_ (_01491_, _01485_, _01490_);
  or _44907_ (_38937_, _01491_, _01489_);
  and _44908_ (_01492_, _01485_, _35826_);
  not _44909_ (_01493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  nor _44910_ (_01494_, _01485_, _01493_);
  or _44911_ (_38938_, _01494_, _01492_);
  and _44912_ (_01495_, _01485_, _35830_);
  not _44913_ (_01496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  nor _44914_ (_01497_, _01485_, _01496_);
  or _44915_ (_38939_, _01497_, _01495_);
  and _44916_ (_01498_, _01485_, _35834_);
  not _44917_ (_01499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  nor _44918_ (_01500_, _01485_, _01499_);
  or _44919_ (_38940_, _01500_, _01498_);
  and _44920_ (_01501_, _01485_, _35838_);
  not _44921_ (_01502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  nor _44922_ (_01503_, _01485_, _01502_);
  or _44923_ (_38941_, _01503_, _01501_);
  and _44924_ (_01504_, _01485_, _35842_);
  not _44925_ (_01505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  nor _44926_ (_01506_, _01485_, _01505_);
  or _44927_ (_38942_, _01506_, _01504_);
  and _44928_ (_01507_, _01485_, _35846_);
  not _44929_ (_01508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  nor _44930_ (_01509_, _01485_, _01508_);
  or _44931_ (_38943_, _01509_, _01507_);
  and _44932_ (_01510_, _00707_, _36622_);
  and _44933_ (_01511_, _01510_, _35572_);
  and _44934_ (_01512_, _01511_, _35815_);
  not _44935_ (_01513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  nor _44936_ (_01514_, _01511_, _01513_);
  or _44937_ (_38944_, _01514_, _01512_);
  and _44938_ (_01515_, _01511_, _35822_);
  not _44939_ (_01516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  nor _44940_ (_01517_, _01511_, _01516_);
  or _44941_ (_38945_, _01517_, _01515_);
  and _44942_ (_01518_, _01511_, _35826_);
  not _44943_ (_01519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  nor _44944_ (_01520_, _01511_, _01519_);
  or _44945_ (_38946_, _01520_, _01518_);
  and _44946_ (_01521_, _01511_, _35830_);
  not _44947_ (_01522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  nor _44948_ (_01523_, _01511_, _01522_);
  or _44949_ (_38947_, _01523_, _01521_);
  and _44950_ (_01524_, _01511_, _35834_);
  not _44951_ (_01525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  nor _44952_ (_01526_, _01511_, _01525_);
  or _44953_ (_38948_, _01526_, _01524_);
  and _44954_ (_01527_, _01511_, _35838_);
  not _44955_ (_01528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  nor _44956_ (_01529_, _01511_, _01528_);
  or _44957_ (_38949_, _01529_, _01527_);
  and _44958_ (_01530_, _01511_, _35842_);
  not _44959_ (_01531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  nor _44960_ (_01532_, _01511_, _01531_);
  or _44961_ (_38950_, _01532_, _01530_);
  and _44962_ (_01533_, _01511_, _35846_);
  not _44963_ (_01534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  nor _44964_ (_01535_, _01511_, _01534_);
  or _44965_ (_38951_, _01535_, _01533_);
  and _44966_ (_01536_, _01510_, _35817_);
  and _44967_ (_01537_, _01536_, _35815_);
  not _44968_ (_01538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  nor _44969_ (_01539_, _01536_, _01538_);
  or _44970_ (_38952_, _01539_, _01537_);
  and _44971_ (_01540_, _01536_, _35822_);
  not _44972_ (_01541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  nor _44973_ (_01542_, _01536_, _01541_);
  or _44974_ (_38953_, _01542_, _01540_);
  and _44975_ (_01543_, _01536_, _35826_);
  not _44976_ (_01544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  nor _44977_ (_01545_, _01536_, _01544_);
  or _44978_ (_38954_, _01545_, _01543_);
  and _44979_ (_01546_, _01536_, _35830_);
  not _44980_ (_01547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  nor _44981_ (_01548_, _01536_, _01547_);
  or _44982_ (_38955_, _01548_, _01546_);
  and _44983_ (_01549_, _01536_, _35834_);
  not _44984_ (_01550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  nor _44985_ (_01551_, _01536_, _01550_);
  or _44986_ (_38956_, _01551_, _01549_);
  and _44987_ (_01552_, _01536_, _35838_);
  not _44988_ (_01553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  nor _44989_ (_01554_, _01536_, _01553_);
  or _44990_ (_38957_, _01554_, _01552_);
  and _44991_ (_01555_, _01536_, _35842_);
  not _44992_ (_01556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  nor _44993_ (_01557_, _01536_, _01556_);
  or _44994_ (_38958_, _01557_, _01555_);
  and _44995_ (_01558_, _01536_, _35846_);
  not _44996_ (_01559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  nor _44997_ (_01560_, _01536_, _01559_);
  or _44998_ (_38959_, _01560_, _01558_);
  and _44999_ (_01561_, _01510_, _35851_);
  and _45000_ (_01562_, _01561_, _35815_);
  not _45001_ (_01563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  nor _45002_ (_01564_, _01561_, _01563_);
  or _45003_ (_38960_, _01564_, _01562_);
  and _45004_ (_01565_, _01561_, _35822_);
  not _45005_ (_01566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  nor _45006_ (_01567_, _01561_, _01566_);
  or _45007_ (_38961_, _01567_, _01565_);
  and _45008_ (_01568_, _01561_, _35826_);
  not _45009_ (_01569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  nor _45010_ (_01570_, _01561_, _01569_);
  or _45011_ (_38962_, _01570_, _01568_);
  and _45012_ (_01571_, _01561_, _35830_);
  not _45013_ (_01572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  nor _45014_ (_01573_, _01561_, _01572_);
  or _45015_ (_38963_, _01573_, _01571_);
  and _45016_ (_01574_, _01561_, _35834_);
  not _45017_ (_01575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  nor _45018_ (_01576_, _01561_, _01575_);
  or _45019_ (_38964_, _01576_, _01574_);
  and _45020_ (_01577_, _01561_, _35838_);
  not _45021_ (_01578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  nor _45022_ (_01579_, _01561_, _01578_);
  or _45023_ (_38965_, _01579_, _01577_);
  and _45024_ (_01580_, _01561_, _35842_);
  not _45025_ (_01581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  nor _45026_ (_01582_, _01561_, _01581_);
  or _45027_ (_38966_, _01582_, _01580_);
  and _45028_ (_01583_, _01561_, _35846_);
  not _45029_ (_01584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  nor _45030_ (_01585_, _01561_, _01584_);
  or _45031_ (_38967_, _01585_, _01583_);
  and _45032_ (_01586_, _01510_, _35878_);
  and _45033_ (_01587_, _01586_, _35815_);
  not _45034_ (_01588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  nor _45035_ (_01589_, _01586_, _01588_);
  or _45036_ (_38968_, _01589_, _01587_);
  and _45037_ (_01590_, _01586_, _35822_);
  not _45038_ (_01591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  nor _45039_ (_01592_, _01586_, _01591_);
  or _45040_ (_38969_, _01592_, _01590_);
  and _45041_ (_01593_, _01586_, _35826_);
  not _45042_ (_01594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  nor _45043_ (_01595_, _01586_, _01594_);
  or _45044_ (_38970_, _01595_, _01593_);
  and _45045_ (_01596_, _01586_, _35830_);
  not _45046_ (_01597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  nor _45047_ (_01598_, _01586_, _01597_);
  or _45048_ (_38971_, _01598_, _01596_);
  and _45049_ (_01599_, _01586_, _35834_);
  not _45050_ (_01600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  nor _45051_ (_01601_, _01586_, _01600_);
  or _45052_ (_38972_, _01601_, _01599_);
  and _45053_ (_01602_, _01586_, _35838_);
  not _45054_ (_01603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  nor _45055_ (_01604_, _01586_, _01603_);
  or _45056_ (_38973_, _01604_, _01602_);
  and _45057_ (_01605_, _01586_, _35842_);
  not _45058_ (_01606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  nor _45059_ (_01607_, _01586_, _01606_);
  or _45060_ (_38974_, _01607_, _01605_);
  and _45061_ (_01608_, _01586_, _35846_);
  not _45062_ (_01609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  nor _45063_ (_01610_, _01586_, _01609_);
  or _45064_ (_38975_, _01610_, _01608_);
  and _45065_ (_01611_, _01510_, _35905_);
  and _45066_ (_01612_, _01611_, _35815_);
  not _45067_ (_01613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  nor _45068_ (_01614_, _01611_, _01613_);
  or _45069_ (_36936_, _01614_, _01612_);
  and _45070_ (_01615_, _01611_, _35822_);
  not _45071_ (_01616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  nor _45072_ (_01617_, _01611_, _01616_);
  or _45073_ (_36937_, _01617_, _01615_);
  and _45074_ (_01618_, _01611_, _35826_);
  not _45075_ (_01619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  nor _45076_ (_01620_, _01611_, _01619_);
  or _45077_ (_36938_, _01620_, _01618_);
  and _45078_ (_01621_, _01611_, _35830_);
  not _45079_ (_01622_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  nor _45080_ (_01623_, _01611_, _01622_);
  or _45081_ (_36939_, _01623_, _01621_);
  and _45082_ (_01624_, _01611_, _35834_);
  not _45083_ (_01625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  nor _45084_ (_01626_, _01611_, _01625_);
  or _45085_ (_36940_, _01626_, _01624_);
  and _45086_ (_01627_, _01611_, _35838_);
  not _45087_ (_01628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  nor _45088_ (_01629_, _01611_, _01628_);
  or _45089_ (_36941_, _01629_, _01627_);
  and _45090_ (_01630_, _01611_, _35842_);
  not _45091_ (_01631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  nor _45092_ (_01632_, _01611_, _01631_);
  or _45093_ (_36942_, _01632_, _01630_);
  and _45094_ (_01633_, _01611_, _35846_);
  not _45095_ (_01634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  nor _45096_ (_01635_, _01611_, _01634_);
  or _45097_ (_36943_, _01635_, _01633_);
  and _45098_ (_01636_, _01510_, _35931_);
  and _45099_ (_01637_, _01636_, _35815_);
  not _45100_ (_01638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  nor _45101_ (_01639_, _01636_, _01638_);
  or _45102_ (_36944_, _01639_, _01637_);
  and _45103_ (_01640_, _01636_, _35822_);
  not _45104_ (_01641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  nor _45105_ (_01642_, _01636_, _01641_);
  or _45106_ (_36945_, _01642_, _01640_);
  and _45107_ (_01643_, _01636_, _35826_);
  not _45108_ (_01644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  nor _45109_ (_01645_, _01636_, _01644_);
  or _45110_ (_36946_, _01645_, _01643_);
  and _45111_ (_01646_, _01636_, _35830_);
  not _45112_ (_01647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  nor _45113_ (_01648_, _01636_, _01647_);
  or _45114_ (_36947_, _01648_, _01646_);
  and _45115_ (_01649_, _01636_, _35834_);
  not _45116_ (_01650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  nor _45117_ (_01651_, _01636_, _01650_);
  or _45118_ (_36948_, _01651_, _01649_);
  and _45119_ (_01652_, _01636_, _35838_);
  not _45120_ (_01653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  nor _45121_ (_01654_, _01636_, _01653_);
  or _45122_ (_36949_, _01654_, _01652_);
  and _45123_ (_01655_, _01636_, _35842_);
  not _45124_ (_01656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  nor _45125_ (_01657_, _01636_, _01656_);
  or _45126_ (_36950_, _01657_, _01655_);
  and _45127_ (_01658_, _01636_, _35846_);
  not _45128_ (_01659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  nor _45129_ (_01660_, _01636_, _01659_);
  or _45130_ (_36951_, _01660_, _01658_);
  and _45131_ (_01661_, _01510_, _35957_);
  and _45132_ (_01662_, _01661_, _35815_);
  not _45133_ (_01663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  nor _45134_ (_01664_, _01661_, _01663_);
  or _45135_ (_36952_, _01664_, _01662_);
  and _45136_ (_01665_, _01661_, _35822_);
  not _45137_ (_01666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  nor _45138_ (_01667_, _01661_, _01666_);
  or _45139_ (_36953_, _01667_, _01665_);
  and _45140_ (_01668_, _01661_, _35826_);
  not _45141_ (_01669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  nor _45142_ (_01670_, _01661_, _01669_);
  or _45143_ (_36954_, _01670_, _01668_);
  and _45144_ (_01671_, _01661_, _35830_);
  not _45145_ (_01672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  nor _45146_ (_01673_, _01661_, _01672_);
  or _45147_ (_36955_, _01673_, _01671_);
  and _45148_ (_01674_, _01661_, _35834_);
  not _45149_ (_01675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  nor _45150_ (_01676_, _01661_, _01675_);
  or _45151_ (_36956_, _01676_, _01674_);
  and _45152_ (_01677_, _01661_, _35838_);
  not _45153_ (_01678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  nor _45154_ (_01679_, _01661_, _01678_);
  or _45155_ (_36957_, _01679_, _01677_);
  and _45156_ (_01680_, _01661_, _35842_);
  not _45157_ (_01681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  nor _45158_ (_01682_, _01661_, _01681_);
  or _45159_ (_36958_, _01682_, _01680_);
  and _45160_ (_01683_, _01661_, _35846_);
  not _45161_ (_01684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  nor _45162_ (_01685_, _01661_, _01684_);
  or _45163_ (_36959_, _01685_, _01683_);
  and _45164_ (_01686_, _01510_, _35983_);
  and _45165_ (_01687_, _01686_, _35815_);
  not _45166_ (_01688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  nor _45167_ (_01689_, _01686_, _01688_);
  or _45168_ (_36960_, _01689_, _01687_);
  and _45169_ (_01690_, _01686_, _35822_);
  not _45170_ (_01691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  nor _45171_ (_01692_, _01686_, _01691_);
  or _45172_ (_36961_, _01692_, _01690_);
  and _45173_ (_01693_, _01686_, _35826_);
  not _45174_ (_01694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  nor _45175_ (_01695_, _01686_, _01694_);
  or _45176_ (_36962_, _01695_, _01693_);
  and _45177_ (_01696_, _01686_, _35830_);
  not _45178_ (_01697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  nor _45179_ (_01698_, _01686_, _01697_);
  or _45180_ (_36963_, _01698_, _01696_);
  and _45181_ (_01699_, _01686_, _35834_);
  not _45182_ (_01700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  nor _45183_ (_01701_, _01686_, _01700_);
  or _45184_ (_36964_, _01701_, _01699_);
  and _45185_ (_01702_, _01686_, _35838_);
  not _45186_ (_01703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  nor _45187_ (_01704_, _01686_, _01703_);
  or _45188_ (_36965_, _01704_, _01702_);
  and _45189_ (_01705_, _01686_, _35842_);
  not _45190_ (_01706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  nor _45191_ (_01707_, _01686_, _01706_);
  or _45192_ (_36966_, _01707_, _01705_);
  and _45193_ (_01708_, _01686_, _35846_);
  not _45194_ (_01709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  nor _45195_ (_01710_, _01686_, _01709_);
  or _45196_ (_36967_, _01710_, _01708_);
  and _45197_ (_01711_, _01510_, _36010_);
  and _45198_ (_01712_, _01711_, _35815_);
  not _45199_ (_01713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  nor _45200_ (_01714_, _01711_, _01713_);
  or _45201_ (_36968_, _01714_, _01712_);
  and _45202_ (_01715_, _01711_, _35822_);
  not _45203_ (_01716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  nor _45204_ (_01717_, _01711_, _01716_);
  or _45205_ (_36969_, _01717_, _01715_);
  and _45206_ (_01718_, _01711_, _35826_);
  not _45207_ (_01719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  nor _45208_ (_01720_, _01711_, _01719_);
  or _45209_ (_36970_, _01720_, _01718_);
  and _45210_ (_01721_, _01711_, _35830_);
  not _45211_ (_01722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  nor _45212_ (_01723_, _01711_, _01722_);
  or _45213_ (_36971_, _01723_, _01721_);
  and _45214_ (_01724_, _01711_, _35834_);
  not _45215_ (_01725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  nor _45216_ (_01726_, _01711_, _01725_);
  or _45217_ (_36972_, _01726_, _01724_);
  and _45218_ (_01727_, _01711_, _35838_);
  not _45219_ (_01728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  nor _45220_ (_01729_, _01711_, _01728_);
  or _45221_ (_36973_, _01729_, _01727_);
  and _45222_ (_01730_, _01711_, _35842_);
  not _45223_ (_01731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  nor _45224_ (_01732_, _01711_, _01731_);
  or _45225_ (_36974_, _01732_, _01730_);
  and _45226_ (_01733_, _01711_, _35846_);
  not _45227_ (_01734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  nor _45228_ (_01735_, _01711_, _01734_);
  or _45229_ (_36975_, _01735_, _01733_);
  and _45230_ (_01736_, _01510_, _36036_);
  and _45231_ (_01737_, _01736_, _35815_);
  not _45232_ (_01738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  nor _45233_ (_01739_, _01736_, _01738_);
  or _45234_ (_36976_, _01739_, _01737_);
  and _45235_ (_01740_, _01736_, _35822_);
  not _45236_ (_01741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  nor _45237_ (_01742_, _01736_, _01741_);
  or _45238_ (_36977_, _01742_, _01740_);
  and _45239_ (_01743_, _01736_, _35826_);
  not _45240_ (_01744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  nor _45241_ (_01745_, _01736_, _01744_);
  or _45242_ (_36978_, _01745_, _01743_);
  and _45243_ (_01746_, _01736_, _35830_);
  not _45244_ (_01747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  nor _45245_ (_01748_, _01736_, _01747_);
  or _45246_ (_36979_, _01748_, _01746_);
  and _45247_ (_01749_, _01736_, _35834_);
  not _45248_ (_01750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  nor _45249_ (_01751_, _01736_, _01750_);
  or _45250_ (_36980_, _01751_, _01749_);
  and _45251_ (_01752_, _01736_, _35838_);
  not _45252_ (_01753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  nor _45253_ (_01754_, _01736_, _01753_);
  or _45254_ (_36981_, _01754_, _01752_);
  and _45255_ (_01755_, _01736_, _35842_);
  not _45256_ (_01756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  nor _45257_ (_01757_, _01736_, _01756_);
  or _45258_ (_36982_, _01757_, _01755_);
  and _45259_ (_01758_, _01736_, _35846_);
  not _45260_ (_01759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  nor _45261_ (_01760_, _01736_, _01759_);
  or _45262_ (_36983_, _01760_, _01758_);
  and _45263_ (_01761_, _01510_, _36062_);
  and _45264_ (_01762_, _01761_, _35815_);
  not _45265_ (_01763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  nor _45266_ (_01764_, _01761_, _01763_);
  or _45267_ (_36984_, _01764_, _01762_);
  and _45268_ (_01765_, _01761_, _35822_);
  not _45269_ (_01766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  nor _45270_ (_01767_, _01761_, _01766_);
  or _45271_ (_36985_, _01767_, _01765_);
  and _45272_ (_01768_, _01761_, _35826_);
  not _45273_ (_01769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  nor _45274_ (_01770_, _01761_, _01769_);
  or _45275_ (_36986_, _01770_, _01768_);
  and _45276_ (_01771_, _01761_, _35830_);
  not _45277_ (_01772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  nor _45278_ (_01773_, _01761_, _01772_);
  or _45279_ (_36987_, _01773_, _01771_);
  and _45280_ (_01774_, _01761_, _35834_);
  not _45281_ (_01775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  nor _45282_ (_01776_, _01761_, _01775_);
  or _45283_ (_36988_, _01776_, _01774_);
  and _45284_ (_01777_, _01761_, _35838_);
  not _45285_ (_01778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  nor _45286_ (_01779_, _01761_, _01778_);
  or _45287_ (_36989_, _01779_, _01777_);
  and _45288_ (_01780_, _01761_, _35842_);
  not _45289_ (_01781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  nor _45290_ (_01782_, _01761_, _01781_);
  or _45291_ (_36990_, _01782_, _01780_);
  and _45292_ (_01783_, _01761_, _35846_);
  not _45293_ (_01784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  nor _45294_ (_01785_, _01761_, _01784_);
  or _45295_ (_36991_, _01785_, _01783_);
  and _45296_ (_01786_, _01510_, _36088_);
  and _45297_ (_01787_, _01786_, _35815_);
  not _45298_ (_01788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  nor _45299_ (_01789_, _01786_, _01788_);
  or _45300_ (_36992_, _01789_, _01787_);
  and _45301_ (_01790_, _01786_, _35822_);
  not _45302_ (_01791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  nor _45303_ (_01792_, _01786_, _01791_);
  or _45304_ (_36993_, _01792_, _01790_);
  and _45305_ (_01793_, _01786_, _35826_);
  not _45306_ (_01794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  nor _45307_ (_01795_, _01786_, _01794_);
  or _45308_ (_36994_, _01795_, _01793_);
  and _45309_ (_01796_, _01786_, _35830_);
  not _45310_ (_01797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  nor _45311_ (_01798_, _01786_, _01797_);
  or _45312_ (_36995_, _01798_, _01796_);
  and _45313_ (_01799_, _01786_, _35834_);
  not _45314_ (_01800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  nor _45315_ (_01801_, _01786_, _01800_);
  or _45316_ (_36996_, _01801_, _01799_);
  and _45317_ (_01802_, _01786_, _35838_);
  not _45318_ (_01803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  nor _45319_ (_01804_, _01786_, _01803_);
  or _45320_ (_36997_, _01804_, _01802_);
  and _45321_ (_01805_, _01786_, _35842_);
  not _45322_ (_01806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  nor _45323_ (_01807_, _01786_, _01806_);
  or _45324_ (_36998_, _01807_, _01805_);
  and _45325_ (_01808_, _01786_, _35846_);
  not _45326_ (_01809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  nor _45327_ (_01810_, _01786_, _01809_);
  or _45328_ (_36999_, _01810_, _01808_);
  and _45329_ (_01811_, _01510_, _36115_);
  and _45330_ (_01812_, _01811_, _35815_);
  not _45331_ (_01813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  nor _45332_ (_01814_, _01811_, _01813_);
  or _45333_ (_37000_, _01814_, _01812_);
  and _45334_ (_01815_, _01811_, _35822_);
  not _45335_ (_01816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  nor _45336_ (_01817_, _01811_, _01816_);
  or _45337_ (_37001_, _01817_, _01815_);
  and _45338_ (_01818_, _01811_, _35826_);
  not _45339_ (_01819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  nor _45340_ (_01820_, _01811_, _01819_);
  or _45341_ (_37002_, _01820_, _01818_);
  and _45342_ (_01821_, _01811_, _35830_);
  not _45343_ (_01822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  nor _45344_ (_01823_, _01811_, _01822_);
  or _45345_ (_37003_, _01823_, _01821_);
  and _45346_ (_01824_, _01811_, _35834_);
  not _45347_ (_01825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  nor _45348_ (_01826_, _01811_, _01825_);
  or _45349_ (_37004_, _01826_, _01824_);
  and _45350_ (_01827_, _01811_, _35838_);
  not _45351_ (_01828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  nor _45352_ (_01829_, _01811_, _01828_);
  or _45353_ (_37005_, _01829_, _01827_);
  and _45354_ (_01830_, _01811_, _35842_);
  not _45355_ (_01831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  nor _45356_ (_01832_, _01811_, _01831_);
  or _45357_ (_37006_, _01832_, _01830_);
  and _45358_ (_01833_, _01811_, _35846_);
  not _45359_ (_01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  nor _45360_ (_01835_, _01811_, _01834_);
  or _45361_ (_37007_, _01835_, _01833_);
  and _45362_ (_01836_, _01510_, _36141_);
  and _45363_ (_01837_, _01836_, _35815_);
  not _45364_ (_01838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  nor _45365_ (_01839_, _01836_, _01838_);
  or _45366_ (_37008_, _01839_, _01837_);
  and _45367_ (_01840_, _01836_, _35822_);
  not _45368_ (_01841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  nor _45369_ (_01842_, _01836_, _01841_);
  or _45370_ (_37009_, _01842_, _01840_);
  and _45371_ (_01843_, _01836_, _35826_);
  not _45372_ (_01844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  nor _45373_ (_01845_, _01836_, _01844_);
  or _45374_ (_37010_, _01845_, _01843_);
  and _45375_ (_01846_, _01836_, _35830_);
  not _45376_ (_01847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  nor _45377_ (_01848_, _01836_, _01847_);
  or _45378_ (_37011_, _01848_, _01846_);
  and _45379_ (_01849_, _01836_, _35834_);
  not _45380_ (_01850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  nor _45381_ (_01851_, _01836_, _01850_);
  or _45382_ (_37012_, _01851_, _01849_);
  and _45383_ (_01852_, _01836_, _35838_);
  not _45384_ (_01853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  nor _45385_ (_01854_, _01836_, _01853_);
  or _45386_ (_37013_, _01854_, _01852_);
  and _45387_ (_01855_, _01836_, _35842_);
  not _45388_ (_01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  nor _45389_ (_01857_, _01836_, _01856_);
  or _45390_ (_37014_, _01857_, _01855_);
  and _45391_ (_01858_, _01836_, _35846_);
  not _45392_ (_01859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  nor _45393_ (_01860_, _01836_, _01859_);
  or _45394_ (_37015_, _01860_, _01858_);
  and _45395_ (_01861_, _01510_, _36167_);
  and _45396_ (_01862_, _01861_, _35815_);
  not _45397_ (_01863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  nor _45398_ (_01864_, _01861_, _01863_);
  or _45399_ (_37024_, _01864_, _01862_);
  and _45400_ (_01865_, _01861_, _35822_);
  not _45401_ (_01866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  nor _45402_ (_01867_, _01861_, _01866_);
  or _45403_ (_37025_, _01867_, _01865_);
  and _45404_ (_01868_, _01861_, _35826_);
  not _45405_ (_01869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  nor _45406_ (_01870_, _01861_, _01869_);
  or _45407_ (_37026_, _01870_, _01868_);
  and _45408_ (_01871_, _01861_, _35830_);
  not _45409_ (_01872_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  nor _45410_ (_01873_, _01861_, _01872_);
  or _45411_ (_37027_, _01873_, _01871_);
  and _45412_ (_01874_, _01861_, _35834_);
  not _45413_ (_01875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  nor _45414_ (_01876_, _01861_, _01875_);
  or _45415_ (_37028_, _01876_, _01874_);
  and _45416_ (_01877_, _01861_, _35838_);
  not _45417_ (_01878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  nor _45418_ (_01879_, _01861_, _01878_);
  or _45419_ (_37029_, _01879_, _01877_);
  and _45420_ (_01880_, _01861_, _35842_);
  not _45421_ (_01881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  nor _45422_ (_01882_, _01861_, _01881_);
  or _45423_ (_37030_, _01882_, _01880_);
  and _45424_ (_01883_, _01861_, _35846_);
  not _45425_ (_01884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  nor _45426_ (_01885_, _01861_, _01884_);
  or _45427_ (_37031_, _01885_, _01883_);
  and _45428_ (_01886_, _01510_, _36193_);
  and _45429_ (_01887_, _01886_, _35815_);
  not _45430_ (_01888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  nor _45431_ (_01889_, _01886_, _01888_);
  or _45432_ (_37032_, _01889_, _01887_);
  and _45433_ (_01890_, _01886_, _35822_);
  not _45434_ (_01891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  nor _45435_ (_01892_, _01886_, _01891_);
  or _45436_ (_37033_, _01892_, _01890_);
  and _45437_ (_01893_, _01886_, _35826_);
  not _45438_ (_01894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  nor _45439_ (_01895_, _01886_, _01894_);
  or _45440_ (_37034_, _01895_, _01893_);
  and _45441_ (_01896_, _01886_, _35830_);
  not _45442_ (_01897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  nor _45443_ (_01898_, _01886_, _01897_);
  or _45444_ (_37035_, _01898_, _01896_);
  and _45445_ (_01899_, _01886_, _35834_);
  not _45446_ (_01900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  nor _45447_ (_01901_, _01886_, _01900_);
  or _45448_ (_37036_, _01901_, _01899_);
  and _45449_ (_01902_, _01886_, _35838_);
  not _45450_ (_01903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  nor _45451_ (_01904_, _01886_, _01903_);
  or _45452_ (_37037_, _01904_, _01902_);
  and _45453_ (_01905_, _01886_, _35842_);
  not _45454_ (_01906_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  nor _45455_ (_01907_, _01886_, _01906_);
  or _45456_ (_37038_, _01907_, _01905_);
  and _45457_ (_01908_, _01886_, _35846_);
  not _45458_ (_01909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  nor _45459_ (_01910_, _01886_, _01909_);
  or _45460_ (_37039_, _01910_, _01908_);
  and _45461_ (_01911_, _00707_, _00304_);
  and _45462_ (_01912_, _01911_, _35572_);
  and _45463_ (_01913_, _01912_, _35815_);
  not _45464_ (_01914_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  nor _45465_ (_01915_, _01912_, _01914_);
  or _45466_ (_37040_, _01915_, _01913_);
  and _45467_ (_01916_, _01912_, _35822_);
  not _45468_ (_01917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  nor _45469_ (_01918_, _01912_, _01917_);
  or _45470_ (_37041_, _01918_, _01916_);
  and _45471_ (_01919_, _01912_, _35826_);
  not _45472_ (_01920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  nor _45473_ (_01921_, _01912_, _01920_);
  or _45474_ (_37042_, _01921_, _01919_);
  and _45475_ (_01922_, _01912_, _35830_);
  not _45476_ (_01923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  nor _45477_ (_01924_, _01912_, _01923_);
  or _45478_ (_37043_, _01924_, _01922_);
  and _45479_ (_01925_, _01912_, _35834_);
  not _45480_ (_01926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  nor _45481_ (_01927_, _01912_, _01926_);
  or _45482_ (_37044_, _01927_, _01925_);
  and _45483_ (_01928_, _01912_, _35838_);
  not _45484_ (_01929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  nor _45485_ (_01930_, _01912_, _01929_);
  or _45486_ (_37045_, _01930_, _01928_);
  and _45487_ (_01931_, _01912_, _35842_);
  not _45488_ (_01932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  nor _45489_ (_01933_, _01912_, _01932_);
  or _45490_ (_37046_, _01933_, _01931_);
  and _45491_ (_01934_, _01912_, _35846_);
  not _45492_ (_01935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  nor _45493_ (_01936_, _01912_, _01935_);
  or _45494_ (_37047_, _01936_, _01934_);
  and _45495_ (_01937_, _01911_, _35817_);
  and _45496_ (_01938_, _01937_, _35815_);
  not _45497_ (_01939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  nor _45498_ (_01940_, _01937_, _01939_);
  or _45499_ (_37048_, _01940_, _01938_);
  and _45500_ (_01941_, _01937_, _35822_);
  not _45501_ (_01942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  nor _45502_ (_01943_, _01937_, _01942_);
  or _45503_ (_37049_, _01943_, _01941_);
  and _45504_ (_01944_, _01937_, _35826_);
  not _45505_ (_01945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  nor _45506_ (_01946_, _01937_, _01945_);
  or _45507_ (_37050_, _01946_, _01944_);
  and _45508_ (_01947_, _01937_, _35830_);
  not _45509_ (_01948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  nor _45510_ (_01949_, _01937_, _01948_);
  or _45511_ (_37051_, _01949_, _01947_);
  and _45512_ (_01950_, _01937_, _35834_);
  not _45513_ (_01951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  nor _45514_ (_01952_, _01937_, _01951_);
  or _45515_ (_37052_, _01952_, _01950_);
  and _45516_ (_01953_, _01937_, _35838_);
  not _45517_ (_01954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  nor _45518_ (_01955_, _01937_, _01954_);
  or _45519_ (_37053_, _01955_, _01953_);
  and _45520_ (_01956_, _01937_, _35842_);
  not _45521_ (_01957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  nor _45522_ (_01958_, _01937_, _01957_);
  or _45523_ (_37054_, _01958_, _01956_);
  and _45524_ (_01959_, _01937_, _35846_);
  not _45525_ (_01960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  nor _45526_ (_01961_, _01937_, _01960_);
  or _45527_ (_37055_, _01961_, _01959_);
  and _45528_ (_01962_, _01911_, _35851_);
  and _45529_ (_01963_, _01962_, _35815_);
  not _45530_ (_01964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  nor _45531_ (_01965_, _01962_, _01964_);
  or _45532_ (_37056_, _01965_, _01963_);
  and _45533_ (_01966_, _01962_, _35822_);
  not _45534_ (_01967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  nor _45535_ (_01968_, _01962_, _01967_);
  or _45536_ (_37057_, _01968_, _01966_);
  and _45537_ (_01969_, _01962_, _35826_);
  not _45538_ (_01970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  nor _45539_ (_01971_, _01962_, _01970_);
  or _45540_ (_37058_, _01971_, _01969_);
  and _45541_ (_01972_, _01962_, _35830_);
  not _45542_ (_01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  nor _45543_ (_01974_, _01962_, _01973_);
  or _45544_ (_37059_, _01974_, _01972_);
  and _45545_ (_01975_, _01962_, _35834_);
  not _45546_ (_01976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  nor _45547_ (_01977_, _01962_, _01976_);
  or _45548_ (_37060_, _01977_, _01975_);
  and _45549_ (_01978_, _01962_, _35838_);
  not _45550_ (_01979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  nor _45551_ (_01980_, _01962_, _01979_);
  or _45552_ (_37061_, _01980_, _01978_);
  and _45553_ (_01981_, _01962_, _35842_);
  not _45554_ (_01982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  nor _45555_ (_01983_, _01962_, _01982_);
  or _45556_ (_37062_, _01983_, _01981_);
  and _45557_ (_01984_, _01962_, _35846_);
  not _45558_ (_01985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  nor _45559_ (_01986_, _01962_, _01985_);
  or _45560_ (_37063_, _01986_, _01984_);
  and _45561_ (_01987_, _01911_, _35878_);
  and _45562_ (_01988_, _01987_, _35815_);
  not _45563_ (_01989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  nor _45564_ (_01990_, _01987_, _01989_);
  or _45565_ (_37064_, _01990_, _01988_);
  and _45566_ (_01991_, _01987_, _35822_);
  not _45567_ (_01992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  nor _45568_ (_01993_, _01987_, _01992_);
  or _45569_ (_37065_, _01993_, _01991_);
  and _45570_ (_01994_, _01987_, _35826_);
  not _45571_ (_01995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  nor _45572_ (_01996_, _01987_, _01995_);
  or _45573_ (_37066_, _01996_, _01994_);
  and _45574_ (_01997_, _01987_, _35830_);
  not _45575_ (_01998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  nor _45576_ (_01999_, _01987_, _01998_);
  or _45577_ (_37067_, _01999_, _01997_);
  and _45578_ (_02000_, _01987_, _35834_);
  not _45579_ (_02001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  nor _45580_ (_02002_, _01987_, _02001_);
  or _45581_ (_37068_, _02002_, _02000_);
  and _45582_ (_02003_, _01987_, _35838_);
  not _45583_ (_02004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  nor _45584_ (_02005_, _01987_, _02004_);
  or _45585_ (_37069_, _02005_, _02003_);
  and _45586_ (_02006_, _01987_, _35842_);
  not _45587_ (_02007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  nor _45588_ (_02008_, _01987_, _02007_);
  or _45589_ (_37070_, _02008_, _02006_);
  and _45590_ (_02009_, _01987_, _35846_);
  not _45591_ (_02010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  nor _45592_ (_02011_, _01987_, _02010_);
  or _45593_ (_37071_, _02011_, _02009_);
  and _45594_ (_02012_, _01911_, _35905_);
  and _45595_ (_02013_, _02012_, _35815_);
  not _45596_ (_02014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  nor _45597_ (_02015_, _02012_, _02014_);
  or _45598_ (_37072_, _02015_, _02013_);
  and _45599_ (_02016_, _02012_, _35822_);
  not _45600_ (_02017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  nor _45601_ (_02018_, _02012_, _02017_);
  or _45602_ (_37073_, _02018_, _02016_);
  and _45603_ (_02019_, _02012_, _35826_);
  not _45604_ (_02020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  nor _45605_ (_02021_, _02012_, _02020_);
  or _45606_ (_37074_, _02021_, _02019_);
  and _45607_ (_02022_, _02012_, _35830_);
  not _45608_ (_02023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  nor _45609_ (_02024_, _02012_, _02023_);
  or _45610_ (_37075_, _02024_, _02022_);
  and _45611_ (_02025_, _02012_, _35834_);
  not _45612_ (_02026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  nor _45613_ (_02027_, _02012_, _02026_);
  or _45614_ (_37076_, _02027_, _02025_);
  and _45615_ (_02028_, _02012_, _35838_);
  not _45616_ (_02029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  nor _45617_ (_02030_, _02012_, _02029_);
  or _45618_ (_37077_, _02030_, _02028_);
  and _45619_ (_02031_, _02012_, _35842_);
  not _45620_ (_02032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  nor _45621_ (_02033_, _02012_, _02032_);
  or _45622_ (_37078_, _02033_, _02031_);
  and _45623_ (_02034_, _02012_, _35846_);
  not _45624_ (_02035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  nor _45625_ (_02036_, _02012_, _02035_);
  or _45626_ (_37079_, _02036_, _02034_);
  and _45627_ (_02037_, _01911_, _35931_);
  and _45628_ (_02038_, _02037_, _35815_);
  not _45629_ (_02039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  nor _45630_ (_02040_, _02037_, _02039_);
  or _45631_ (_37080_, _02040_, _02038_);
  and _45632_ (_02041_, _02037_, _35822_);
  not _45633_ (_02042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  nor _45634_ (_02043_, _02037_, _02042_);
  or _45635_ (_37081_, _02043_, _02041_);
  and _45636_ (_02044_, _02037_, _35826_);
  not _45637_ (_02045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  nor _45638_ (_02046_, _02037_, _02045_);
  or _45639_ (_37082_, _02046_, _02044_);
  and _45640_ (_02047_, _02037_, _35830_);
  not _45641_ (_02048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  nor _45642_ (_02049_, _02037_, _02048_);
  or _45643_ (_37083_, _02049_, _02047_);
  and _45644_ (_02050_, _02037_, _35834_);
  not _45645_ (_02051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  nor _45646_ (_02052_, _02037_, _02051_);
  or _45647_ (_37084_, _02052_, _02050_);
  and _45648_ (_02053_, _02037_, _35838_);
  not _45649_ (_02054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  nor _45650_ (_02055_, _02037_, _02054_);
  or _45651_ (_37085_, _02055_, _02053_);
  and _45652_ (_02056_, _02037_, _35842_);
  not _45653_ (_02057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  nor _45654_ (_02058_, _02037_, _02057_);
  or _45655_ (_37086_, _02058_, _02056_);
  and _45656_ (_02059_, _02037_, _35846_);
  not _45657_ (_02060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  nor _45658_ (_02061_, _02037_, _02060_);
  or _45659_ (_37087_, _02061_, _02059_);
  and _45660_ (_02062_, _01911_, _35957_);
  and _45661_ (_02063_, _02062_, _35815_);
  not _45662_ (_02064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  nor _45663_ (_02065_, _02062_, _02064_);
  or _45664_ (_37088_, _02065_, _02063_);
  and _45665_ (_02066_, _02062_, _35822_);
  not _45666_ (_02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  nor _45667_ (_02068_, _02062_, _02067_);
  or _45668_ (_37089_, _02068_, _02066_);
  and _45669_ (_02069_, _02062_, _35826_);
  not _45670_ (_02070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  nor _45671_ (_02071_, _02062_, _02070_);
  or _45672_ (_37090_, _02071_, _02069_);
  and _45673_ (_02072_, _02062_, _35830_);
  not _45674_ (_02073_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  nor _45675_ (_02074_, _02062_, _02073_);
  or _45676_ (_37091_, _02074_, _02072_);
  and _45677_ (_02075_, _02062_, _35834_);
  not _45678_ (_02076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  nor _45679_ (_02077_, _02062_, _02076_);
  or _45680_ (_37092_, _02077_, _02075_);
  and _45681_ (_02078_, _02062_, _35838_);
  not _45682_ (_02079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  nor _45683_ (_02080_, _02062_, _02079_);
  or _45684_ (_37093_, _02080_, _02078_);
  and _45685_ (_02081_, _02062_, _35842_);
  not _45686_ (_02082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  nor _45687_ (_02083_, _02062_, _02082_);
  or _45688_ (_37094_, _02083_, _02081_);
  and _45689_ (_02084_, _02062_, _35846_);
  not _45690_ (_02085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  nor _45691_ (_02086_, _02062_, _02085_);
  or _45692_ (_37095_, _02086_, _02084_);
  and _45693_ (_02087_, _01911_, _35983_);
  and _45694_ (_02088_, _02087_, _35815_);
  not _45695_ (_02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  nor _45696_ (_02090_, _02087_, _02089_);
  or _45697_ (_37096_, _02090_, _02088_);
  and _45698_ (_02091_, _02087_, _35822_);
  not _45699_ (_02092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  nor _45700_ (_02093_, _02087_, _02092_);
  or _45701_ (_37097_, _02093_, _02091_);
  and _45702_ (_02094_, _02087_, _35826_);
  not _45703_ (_02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  nor _45704_ (_02096_, _02087_, _02095_);
  or _45705_ (_37098_, _02096_, _02094_);
  and _45706_ (_02097_, _02087_, _35830_);
  not _45707_ (_02098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  nor _45708_ (_02099_, _02087_, _02098_);
  or _45709_ (_37099_, _02099_, _02097_);
  and _45710_ (_02100_, _02087_, _35834_);
  not _45711_ (_02101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  nor _45712_ (_02102_, _02087_, _02101_);
  or _45713_ (_37100_, _02102_, _02100_);
  and _45714_ (_02103_, _02087_, _35838_);
  not _45715_ (_02104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  nor _45716_ (_02105_, _02087_, _02104_);
  or _45717_ (_37101_, _02105_, _02103_);
  and _45718_ (_02106_, _02087_, _35842_);
  not _45719_ (_02107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  nor _45720_ (_02108_, _02087_, _02107_);
  or _45721_ (_37102_, _02108_, _02106_);
  and _45722_ (_02109_, _02087_, _35846_);
  not _45723_ (_02110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  nor _45724_ (_02111_, _02087_, _02110_);
  or _45725_ (_37103_, _02111_, _02109_);
  and _45726_ (_02112_, _01911_, _36010_);
  and _45727_ (_02113_, _02112_, _35815_);
  not _45728_ (_02114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  nor _45729_ (_02115_, _02112_, _02114_);
  or _45730_ (_37112_, _02115_, _02113_);
  and _45731_ (_02116_, _02112_, _35822_);
  not _45732_ (_02117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  nor _45733_ (_02118_, _02112_, _02117_);
  or _45734_ (_37113_, _02118_, _02116_);
  and _45735_ (_02119_, _02112_, _35826_);
  not _45736_ (_02120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  nor _45737_ (_02121_, _02112_, _02120_);
  or _45738_ (_37114_, _02121_, _02119_);
  and _45739_ (_02122_, _02112_, _35830_);
  not _45740_ (_02123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  nor _45741_ (_02124_, _02112_, _02123_);
  or _45742_ (_37115_, _02124_, _02122_);
  and _45743_ (_02125_, _02112_, _35834_);
  not _45744_ (_02126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  nor _45745_ (_02127_, _02112_, _02126_);
  or _45746_ (_37116_, _02127_, _02125_);
  and _45747_ (_02128_, _02112_, _35838_);
  not _45748_ (_02129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  nor _45749_ (_02130_, _02112_, _02129_);
  or _45750_ (_37117_, _02130_, _02128_);
  and _45751_ (_02131_, _02112_, _35842_);
  not _45752_ (_02132_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  nor _45753_ (_02133_, _02112_, _02132_);
  or _45754_ (_37118_, _02133_, _02131_);
  and _45755_ (_02134_, _02112_, _35846_);
  not _45756_ (_02135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  nor _45757_ (_02136_, _02112_, _02135_);
  or _45758_ (_37119_, _02136_, _02134_);
  and _45759_ (_02137_, _01911_, _36036_);
  and _45760_ (_02138_, _02137_, _35815_);
  not _45761_ (_02139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  nor _45762_ (_02140_, _02137_, _02139_);
  or _45763_ (_37120_, _02140_, _02138_);
  and _45764_ (_02141_, _02137_, _35822_);
  not _45765_ (_02142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  nor _45766_ (_02143_, _02137_, _02142_);
  or _45767_ (_37121_, _02143_, _02141_);
  and _45768_ (_02144_, _02137_, _35826_);
  not _45769_ (_02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  nor _45770_ (_02146_, _02137_, _02145_);
  or _45771_ (_37122_, _02146_, _02144_);
  and _45772_ (_02147_, _02137_, _35830_);
  not _45773_ (_02148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  nor _45774_ (_02149_, _02137_, _02148_);
  or _45775_ (_37123_, _02149_, _02147_);
  and _45776_ (_02150_, _02137_, _35834_);
  not _45777_ (_02151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  nor _45778_ (_02152_, _02137_, _02151_);
  or _45779_ (_37124_, _02152_, _02150_);
  and _45780_ (_02153_, _02137_, _35838_);
  not _45781_ (_02154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  nor _45782_ (_02155_, _02137_, _02154_);
  or _45783_ (_37125_, _02155_, _02153_);
  and _45784_ (_02156_, _02137_, _35842_);
  not _45785_ (_02157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  nor _45786_ (_02158_, _02137_, _02157_);
  or _45787_ (_37126_, _02158_, _02156_);
  and _45788_ (_02159_, _02137_, _35846_);
  not _45789_ (_02160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  nor _45790_ (_02161_, _02137_, _02160_);
  or _45791_ (_37127_, _02161_, _02159_);
  and _45792_ (_02162_, _01911_, _36062_);
  and _45793_ (_02163_, _02162_, _35815_);
  not _45794_ (_02164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  nor _45795_ (_02165_, _02162_, _02164_);
  or _45796_ (_37128_, _02165_, _02163_);
  and _45797_ (_02166_, _02162_, _35822_);
  not _45798_ (_02167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  nor _45799_ (_02168_, _02162_, _02167_);
  or _45800_ (_37129_, _02168_, _02166_);
  and _45801_ (_02169_, _02162_, _35826_);
  not _45802_ (_02170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  nor _45803_ (_02171_, _02162_, _02170_);
  or _45804_ (_37130_, _02171_, _02169_);
  and _45805_ (_02172_, _02162_, _35830_);
  not _45806_ (_02173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  nor _45807_ (_02174_, _02162_, _02173_);
  or _45808_ (_37131_, _02174_, _02172_);
  and _45809_ (_02175_, _02162_, _35834_);
  not _45810_ (_02176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  nor _45811_ (_02177_, _02162_, _02176_);
  or _45812_ (_37132_, _02177_, _02175_);
  and _45813_ (_02178_, _02162_, _35838_);
  not _45814_ (_02179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  nor _45815_ (_02180_, _02162_, _02179_);
  or _45816_ (_37133_, _02180_, _02178_);
  and _45817_ (_02181_, _02162_, _35842_);
  not _45818_ (_02182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  nor _45819_ (_02183_, _02162_, _02182_);
  or _45820_ (_37134_, _02183_, _02181_);
  and _45821_ (_02184_, _02162_, _35846_);
  not _45822_ (_02185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  nor _45823_ (_02186_, _02162_, _02185_);
  or _45824_ (_37135_, _02186_, _02184_);
  and _45825_ (_02187_, _01911_, _36088_);
  and _45826_ (_02188_, _02187_, _35815_);
  not _45827_ (_02189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  nor _45828_ (_02190_, _02187_, _02189_);
  or _45829_ (_37136_, _02190_, _02188_);
  and _45830_ (_02191_, _02187_, _35822_);
  not _45831_ (_02192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  nor _45832_ (_02193_, _02187_, _02192_);
  or _45833_ (_37137_, _02193_, _02191_);
  and _45834_ (_02194_, _02187_, _35826_);
  not _45835_ (_02195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  nor _45836_ (_02196_, _02187_, _02195_);
  or _45837_ (_37138_, _02196_, _02194_);
  and _45838_ (_02197_, _02187_, _35830_);
  not _45839_ (_02198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  nor _45840_ (_02199_, _02187_, _02198_);
  or _45841_ (_37139_, _02199_, _02197_);
  and _45842_ (_02200_, _02187_, _35834_);
  not _45843_ (_02201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  nor _45844_ (_02202_, _02187_, _02201_);
  or _45845_ (_37140_, _02202_, _02200_);
  and _45846_ (_02203_, _02187_, _35838_);
  not _45847_ (_02204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  nor _45848_ (_02205_, _02187_, _02204_);
  or _45849_ (_37141_, _02205_, _02203_);
  and _45850_ (_02206_, _02187_, _35842_);
  not _45851_ (_02207_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  nor _45852_ (_02208_, _02187_, _02207_);
  or _45853_ (_37142_, _02208_, _02206_);
  and _45854_ (_02209_, _02187_, _35846_);
  not _45855_ (_02210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  nor _45856_ (_02211_, _02187_, _02210_);
  or _45857_ (_37143_, _02211_, _02209_);
  and _45858_ (_02212_, _01911_, _36115_);
  and _45859_ (_02213_, _02212_, _35815_);
  not _45860_ (_02214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  nor _45861_ (_02215_, _02212_, _02214_);
  or _45862_ (_37144_, _02215_, _02213_);
  and _45863_ (_02216_, _02212_, _35822_);
  not _45864_ (_02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  nor _45865_ (_02218_, _02212_, _02217_);
  or _45866_ (_37145_, _02218_, _02216_);
  and _45867_ (_02219_, _02212_, _35826_);
  not _45868_ (_02220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  nor _45869_ (_02221_, _02212_, _02220_);
  or _45870_ (_37146_, _02221_, _02219_);
  and _45871_ (_02222_, _02212_, _35830_);
  not _45872_ (_02223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  nor _45873_ (_02224_, _02212_, _02223_);
  or _45874_ (_37147_, _02224_, _02222_);
  and _45875_ (_02225_, _02212_, _35834_);
  not _45876_ (_02226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  nor _45877_ (_02227_, _02212_, _02226_);
  or _45878_ (_37148_, _02227_, _02225_);
  and _45879_ (_02228_, _02212_, _35838_);
  not _45880_ (_02229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  nor _45881_ (_02230_, _02212_, _02229_);
  or _45882_ (_37149_, _02230_, _02228_);
  and _45883_ (_02231_, _02212_, _35842_);
  not _45884_ (_02232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  nor _45885_ (_02233_, _02212_, _02232_);
  or _45886_ (_37150_, _02233_, _02231_);
  and _45887_ (_02234_, _02212_, _35846_);
  not _45888_ (_02235_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  nor _45889_ (_02236_, _02212_, _02235_);
  or _45890_ (_37151_, _02236_, _02234_);
  and _45891_ (_02237_, _01911_, _36141_);
  and _45892_ (_02238_, _02237_, _35815_);
  not _45893_ (_02239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  nor _45894_ (_02240_, _02237_, _02239_);
  or _45895_ (_37152_, _02240_, _02238_);
  and _45896_ (_02241_, _02237_, _35822_);
  not _45897_ (_02242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  nor _45898_ (_02243_, _02237_, _02242_);
  or _45899_ (_37153_, _02243_, _02241_);
  and _45900_ (_02244_, _02237_, _35826_);
  not _45901_ (_02245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  nor _45902_ (_02246_, _02237_, _02245_);
  or _45903_ (_37154_, _02246_, _02244_);
  and _45904_ (_02247_, _02237_, _35830_);
  not _45905_ (_02248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  nor _45906_ (_02249_, _02237_, _02248_);
  or _45907_ (_37155_, _02249_, _02247_);
  and _45908_ (_02250_, _02237_, _35834_);
  not _45909_ (_02251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  nor _45910_ (_02252_, _02237_, _02251_);
  or _45911_ (_37156_, _02252_, _02250_);
  and _45912_ (_02253_, _02237_, _35838_);
  not _45913_ (_02254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  nor _45914_ (_02255_, _02237_, _02254_);
  or _45915_ (_37157_, _02255_, _02253_);
  and _45916_ (_02256_, _02237_, _35842_);
  not _45917_ (_02257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  nor _45918_ (_02258_, _02237_, _02257_);
  or _45919_ (_37158_, _02258_, _02256_);
  and _45920_ (_02259_, _02237_, _35846_);
  not _45921_ (_02260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  nor _45922_ (_02261_, _02237_, _02260_);
  or _45923_ (_37159_, _02261_, _02259_);
  and _45924_ (_02262_, _01911_, _36167_);
  and _45925_ (_02263_, _02262_, _35815_);
  not _45926_ (_02264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  nor _45927_ (_02265_, _02262_, _02264_);
  or _45928_ (_37160_, _02265_, _02263_);
  and _45929_ (_02266_, _02262_, _35822_);
  not _45930_ (_02267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  nor _45931_ (_02268_, _02262_, _02267_);
  or _45932_ (_37161_, _02268_, _02266_);
  and _45933_ (_02269_, _02262_, _35826_);
  not _45934_ (_02270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  nor _45935_ (_02271_, _02262_, _02270_);
  or _45936_ (_37162_, _02271_, _02269_);
  and _45937_ (_02272_, _02262_, _35830_);
  not _45938_ (_02273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  nor _45939_ (_02274_, _02262_, _02273_);
  or _45940_ (_37163_, _02274_, _02272_);
  and _45941_ (_02275_, _02262_, _35834_);
  not _45942_ (_02276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  nor _45943_ (_02277_, _02262_, _02276_);
  or _45944_ (_37164_, _02277_, _02275_);
  and _45945_ (_02278_, _02262_, _35838_);
  not _45946_ (_02279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  nor _45947_ (_02280_, _02262_, _02279_);
  or _45948_ (_37165_, _02280_, _02278_);
  and _45949_ (_02281_, _02262_, _35842_);
  not _45950_ (_02282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  nor _45951_ (_02283_, _02262_, _02282_);
  or _45952_ (_37166_, _02283_, _02281_);
  and _45953_ (_02284_, _02262_, _35846_);
  not _45954_ (_02285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  nor _45955_ (_02286_, _02262_, _02285_);
  or _45956_ (_37167_, _02286_, _02284_);
  and _45957_ (_02287_, _01911_, _36193_);
  and _45958_ (_02288_, _02287_, _35815_);
  not _45959_ (_02289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  nor _45960_ (_02290_, _02287_, _02289_);
  or _45961_ (_37168_, _02290_, _02288_);
  and _45962_ (_02291_, _02287_, _35822_);
  not _45963_ (_02292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  nor _45964_ (_02293_, _02287_, _02292_);
  or _45965_ (_37169_, _02293_, _02291_);
  and _45966_ (_02294_, _02287_, _35826_);
  not _45967_ (_02295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  nor _45968_ (_02296_, _02287_, _02295_);
  or _45969_ (_37170_, _02296_, _02294_);
  and _45970_ (_02297_, _02287_, _35830_);
  not _45971_ (_02298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  nor _45972_ (_02299_, _02287_, _02298_);
  or _45973_ (_37171_, _02299_, _02297_);
  and _45974_ (_02300_, _02287_, _35834_);
  not _45975_ (_02301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  nor _45976_ (_02302_, _02287_, _02301_);
  or _45977_ (_37172_, _02302_, _02300_);
  and _45978_ (_02303_, _02287_, _35838_);
  not _45979_ (_02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  nor _45980_ (_02305_, _02287_, _02304_);
  or _45981_ (_37173_, _02305_, _02303_);
  and _45982_ (_02306_, _02287_, _35842_);
  not _45983_ (_02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  nor _45984_ (_02308_, _02287_, _02307_);
  or _45985_ (_37174_, _02308_, _02306_);
  and _45986_ (_02309_, _02287_, _35846_);
  not _45987_ (_02310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  nor _45988_ (_02311_, _02287_, _02310_);
  or _45989_ (_37175_, _02311_, _02309_);
  and _45990_ (_02312_, _34784_, _33632_);
  and _45991_ (_02313_, _02312_, _35575_);
  and _45992_ (_02314_, _02313_, _35572_);
  and _45993_ (_02315_, _02314_, _35815_);
  not _45994_ (_02316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  nor _45995_ (_02317_, _02314_, _02316_);
  or _45996_ (_37176_, _02317_, _02315_);
  and _45997_ (_02318_, _02314_, _35822_);
  not _45998_ (_02319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  nor _45999_ (_02320_, _02314_, _02319_);
  or _46000_ (_37177_, _02320_, _02318_);
  and _46001_ (_02321_, _02314_, _35826_);
  not _46002_ (_02322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  nor _46003_ (_02323_, _02314_, _02322_);
  or _46004_ (_37178_, _02323_, _02321_);
  and _46005_ (_02324_, _02314_, _35830_);
  not _46006_ (_02325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  nor _46007_ (_02326_, _02314_, _02325_);
  or _46008_ (_37179_, _02326_, _02324_);
  and _46009_ (_02327_, _02314_, _35834_);
  not _46010_ (_02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  nor _46011_ (_02329_, _02314_, _02328_);
  or _46012_ (_37180_, _02329_, _02327_);
  and _46013_ (_02330_, _02314_, _35838_);
  not _46014_ (_02331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  nor _46015_ (_02332_, _02314_, _02331_);
  or _46016_ (_37181_, _02332_, _02330_);
  and _46017_ (_02333_, _02314_, _35842_);
  not _46018_ (_02334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  nor _46019_ (_02335_, _02314_, _02334_);
  or _46020_ (_37182_, _02335_, _02333_);
  and _46021_ (_02336_, _02314_, _35846_);
  not _46022_ (_02337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  nor _46023_ (_02338_, _02314_, _02337_);
  or _46024_ (_37183_, _02338_, _02336_);
  and _46025_ (_02339_, _02313_, _35817_);
  and _46026_ (_02340_, _02339_, _35815_);
  not _46027_ (_02341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  nor _46028_ (_02342_, _02339_, _02341_);
  or _46029_ (_37184_, _02342_, _02340_);
  and _46030_ (_02343_, _02339_, _35822_);
  not _46031_ (_02344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  nor _46032_ (_02345_, _02339_, _02344_);
  or _46033_ (_37185_, _02345_, _02343_);
  and _46034_ (_02346_, _02339_, _35826_);
  not _46035_ (_02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  nor _46036_ (_02348_, _02339_, _02347_);
  or _46037_ (_37186_, _02348_, _02346_);
  and _46038_ (_02349_, _02339_, _35830_);
  not _46039_ (_02350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  nor _46040_ (_02351_, _02339_, _02350_);
  or _46041_ (_37187_, _02351_, _02349_);
  and _46042_ (_02352_, _02339_, _35834_);
  not _46043_ (_02353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  nor _46044_ (_02354_, _02339_, _02353_);
  or _46045_ (_37188_, _02354_, _02352_);
  and _46046_ (_02355_, _02339_, _35838_);
  not _46047_ (_02356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  nor _46048_ (_02357_, _02339_, _02356_);
  or _46049_ (_37189_, _02357_, _02355_);
  and _46050_ (_02358_, _02339_, _35842_);
  not _46051_ (_02359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  nor _46052_ (_02360_, _02339_, _02359_);
  or _46053_ (_37190_, _02360_, _02358_);
  and _46054_ (_02361_, _02339_, _35846_);
  not _46055_ (_02362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  nor _46056_ (_02363_, _02339_, _02362_);
  or _46057_ (_37191_, _02363_, _02361_);
  and _46058_ (_02364_, _02313_, _35851_);
  and _46059_ (_02365_, _02364_, _35815_);
  not _46060_ (_02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  nor _46061_ (_02367_, _02364_, _02366_);
  or _46062_ (_37200_, _02367_, _02365_);
  and _46063_ (_02368_, _02364_, _35822_);
  not _46064_ (_02369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  nor _46065_ (_02370_, _02364_, _02369_);
  or _46066_ (_37201_, _02370_, _02368_);
  and _46067_ (_02371_, _02364_, _35826_);
  not _46068_ (_02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  nor _46069_ (_02373_, _02364_, _02372_);
  or _46070_ (_37202_, _02373_, _02371_);
  and _46071_ (_02374_, _02364_, _35830_);
  not _46072_ (_02375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  nor _46073_ (_02376_, _02364_, _02375_);
  or _46074_ (_37203_, _02376_, _02374_);
  and _46075_ (_02377_, _02364_, _35834_);
  not _46076_ (_02378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  nor _46077_ (_02379_, _02364_, _02378_);
  or _46078_ (_37204_, _02379_, _02377_);
  and _46079_ (_02380_, _02364_, _35838_);
  not _46080_ (_02381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  nor _46081_ (_02382_, _02364_, _02381_);
  or _46082_ (_37205_, _02382_, _02380_);
  and _46083_ (_02383_, _02364_, _35842_);
  not _46084_ (_02384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  nor _46085_ (_02385_, _02364_, _02384_);
  or _46086_ (_37206_, _02385_, _02383_);
  and _46087_ (_02386_, _02364_, _35846_);
  not _46088_ (_02387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  nor _46089_ (_02388_, _02364_, _02387_);
  or _46090_ (_37207_, _02388_, _02386_);
  and _46091_ (_02389_, _02313_, _35878_);
  and _46092_ (_02390_, _02389_, _35815_);
  not _46093_ (_02391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  nor _46094_ (_02392_, _02389_, _02391_);
  or _46095_ (_37208_, _02392_, _02390_);
  and _46096_ (_02393_, _02389_, _35822_);
  not _46097_ (_02394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  nor _46098_ (_02395_, _02389_, _02394_);
  or _46099_ (_37209_, _02395_, _02393_);
  and _46100_ (_02396_, _02389_, _35826_);
  not _46101_ (_02397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  nor _46102_ (_02398_, _02389_, _02397_);
  or _46103_ (_37210_, _02398_, _02396_);
  and _46104_ (_02399_, _02389_, _35830_);
  not _46105_ (_02400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  nor _46106_ (_02401_, _02389_, _02400_);
  or _46107_ (_37211_, _02401_, _02399_);
  and _46108_ (_02402_, _02389_, _35834_);
  not _46109_ (_02403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  nor _46110_ (_02404_, _02389_, _02403_);
  or _46111_ (_37212_, _02404_, _02402_);
  and _46112_ (_02405_, _02389_, _35838_);
  not _46113_ (_02406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  nor _46114_ (_02407_, _02389_, _02406_);
  or _46115_ (_37213_, _02407_, _02405_);
  and _46116_ (_02408_, _02389_, _35842_);
  not _46117_ (_02409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  nor _46118_ (_02410_, _02389_, _02409_);
  or _46119_ (_37214_, _02410_, _02408_);
  and _46120_ (_02411_, _02389_, _35846_);
  not _46121_ (_02412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  nor _46122_ (_02413_, _02389_, _02412_);
  or _46123_ (_37215_, _02413_, _02411_);
  and _46124_ (_02414_, _02313_, _35905_);
  and _46125_ (_02415_, _02414_, _35815_);
  not _46126_ (_02416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  nor _46127_ (_02417_, _02414_, _02416_);
  or _46128_ (_37216_, _02417_, _02415_);
  and _46129_ (_02418_, _02414_, _35822_);
  not _46130_ (_02419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  nor _46131_ (_02420_, _02414_, _02419_);
  or _46132_ (_37217_, _02420_, _02418_);
  and _46133_ (_02421_, _02414_, _35826_);
  not _46134_ (_02422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  nor _46135_ (_02423_, _02414_, _02422_);
  or _46136_ (_37218_, _02423_, _02421_);
  and _46137_ (_02424_, _02414_, _35830_);
  not _46138_ (_02425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  nor _46139_ (_02426_, _02414_, _02425_);
  or _46140_ (_37219_, _02426_, _02424_);
  and _46141_ (_02427_, _02414_, _35834_);
  not _46142_ (_02428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  nor _46143_ (_02429_, _02414_, _02428_);
  or _46144_ (_37220_, _02429_, _02427_);
  and _46145_ (_02430_, _02414_, _35838_);
  not _46146_ (_02431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  nor _46147_ (_02432_, _02414_, _02431_);
  or _46148_ (_37221_, _02432_, _02430_);
  and _46149_ (_02433_, _02414_, _35842_);
  not _46150_ (_02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  nor _46151_ (_02435_, _02414_, _02434_);
  or _46152_ (_37222_, _02435_, _02433_);
  and _46153_ (_02436_, _02414_, _35846_);
  not _46154_ (_02437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  nor _46155_ (_02438_, _02414_, _02437_);
  or _46156_ (_37223_, _02438_, _02436_);
  and _46157_ (_02439_, _02313_, _35931_);
  and _46158_ (_02440_, _02439_, _35815_);
  not _46159_ (_02441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  nor _46160_ (_02442_, _02439_, _02441_);
  or _46161_ (_37224_, _02442_, _02440_);
  and _46162_ (_02443_, _02439_, _35822_);
  not _46163_ (_02444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  nor _46164_ (_02445_, _02439_, _02444_);
  or _46165_ (_37225_, _02445_, _02443_);
  and _46166_ (_02446_, _02439_, _35826_);
  not _46167_ (_02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  nor _46168_ (_02448_, _02439_, _02447_);
  or _46169_ (_37226_, _02448_, _02446_);
  and _46170_ (_02449_, _02439_, _35830_);
  not _46171_ (_02450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  nor _46172_ (_02451_, _02439_, _02450_);
  or _46173_ (_37227_, _02451_, _02449_);
  and _46174_ (_02452_, _02439_, _35834_);
  not _46175_ (_02453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  nor _46176_ (_02454_, _02439_, _02453_);
  or _46177_ (_37228_, _02454_, _02452_);
  and _46178_ (_02455_, _02439_, _35838_);
  not _46179_ (_02456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  nor _46180_ (_02457_, _02439_, _02456_);
  or _46181_ (_37229_, _02457_, _02455_);
  and _46182_ (_02458_, _02439_, _35842_);
  not _46183_ (_02459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  nor _46184_ (_02460_, _02439_, _02459_);
  or _46185_ (_37230_, _02460_, _02458_);
  and _46186_ (_02461_, _02439_, _35846_);
  not _46187_ (_02462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  nor _46188_ (_02463_, _02439_, _02462_);
  or _46189_ (_37231_, _02463_, _02461_);
  and _46190_ (_02464_, _02313_, _35957_);
  and _46191_ (_02465_, _02464_, _35815_);
  not _46192_ (_02466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  nor _46193_ (_02467_, _02464_, _02466_);
  or _46194_ (_37232_, _02467_, _02465_);
  and _46195_ (_02468_, _02464_, _35822_);
  not _46196_ (_02469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  nor _46197_ (_02470_, _02464_, _02469_);
  or _46198_ (_37233_, _02470_, _02468_);
  and _46199_ (_02471_, _02464_, _35826_);
  not _46200_ (_02472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  nor _46201_ (_02473_, _02464_, _02472_);
  or _46202_ (_37234_, _02473_, _02471_);
  and _46203_ (_02474_, _02464_, _35830_);
  not _46204_ (_02475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  nor _46205_ (_02476_, _02464_, _02475_);
  or _46206_ (_37235_, _02476_, _02474_);
  and _46207_ (_02477_, _02464_, _35834_);
  not _46208_ (_02478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  nor _46209_ (_02479_, _02464_, _02478_);
  or _46210_ (_37236_, _02479_, _02477_);
  and _46211_ (_02480_, _02464_, _35838_);
  not _46212_ (_02481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  nor _46213_ (_02482_, _02464_, _02481_);
  or _46214_ (_37237_, _02482_, _02480_);
  and _46215_ (_02483_, _02464_, _35842_);
  not _46216_ (_02484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  nor _46217_ (_02485_, _02464_, _02484_);
  or _46218_ (_37238_, _02485_, _02483_);
  and _46219_ (_02486_, _02464_, _35846_);
  not _46220_ (_02487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  nor _46221_ (_02488_, _02464_, _02487_);
  or _46222_ (_37239_, _02488_, _02486_);
  and _46223_ (_02489_, _02313_, _35983_);
  and _46224_ (_02490_, _02489_, _35815_);
  not _46225_ (_02491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  nor _46226_ (_02492_, _02489_, _02491_);
  or _46227_ (_37240_, _02492_, _02490_);
  and _46228_ (_02493_, _02489_, _35822_);
  not _46229_ (_02494_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  nor _46230_ (_02495_, _02489_, _02494_);
  or _46231_ (_37241_, _02495_, _02493_);
  and _46232_ (_02496_, _02489_, _35826_);
  not _46233_ (_02497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  nor _46234_ (_02498_, _02489_, _02497_);
  or _46235_ (_37242_, _02498_, _02496_);
  and _46236_ (_02499_, _02489_, _35830_);
  not _46237_ (_02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  nor _46238_ (_02501_, _02489_, _02500_);
  or _46239_ (_37243_, _02501_, _02499_);
  and _46240_ (_02502_, _02489_, _35834_);
  not _46241_ (_02503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  nor _46242_ (_02504_, _02489_, _02503_);
  or _46243_ (_37244_, _02504_, _02502_);
  and _46244_ (_02505_, _02489_, _35838_);
  not _46245_ (_02506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  nor _46246_ (_02507_, _02489_, _02506_);
  or _46247_ (_37245_, _02507_, _02505_);
  and _46248_ (_02508_, _02489_, _35842_);
  not _46249_ (_02509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  nor _46250_ (_02510_, _02489_, _02509_);
  or _46251_ (_37246_, _02510_, _02508_);
  and _46252_ (_02511_, _02489_, _35846_);
  not _46253_ (_02512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  nor _46254_ (_02513_, _02489_, _02512_);
  or _46255_ (_37247_, _02513_, _02511_);
  and _46256_ (_02514_, _02313_, _36010_);
  and _46257_ (_02515_, _02514_, _35815_);
  not _46258_ (_02516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  nor _46259_ (_02517_, _02514_, _02516_);
  or _46260_ (_37248_, _02517_, _02515_);
  and _46261_ (_02518_, _02514_, _35822_);
  not _46262_ (_02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  nor _46263_ (_02520_, _02514_, _02519_);
  or _46264_ (_37249_, _02520_, _02518_);
  and _46265_ (_02521_, _02514_, _35826_);
  not _46266_ (_02522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  nor _46267_ (_02523_, _02514_, _02522_);
  or _46268_ (_37250_, _02523_, _02521_);
  and _46269_ (_02524_, _02514_, _35830_);
  not _46270_ (_02525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  nor _46271_ (_02526_, _02514_, _02525_);
  or _46272_ (_37251_, _02526_, _02524_);
  and _46273_ (_02527_, _02514_, _35834_);
  not _46274_ (_02528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  nor _46275_ (_02529_, _02514_, _02528_);
  or _46276_ (_37252_, _02529_, _02527_);
  and _46277_ (_02530_, _02514_, _35838_);
  not _46278_ (_02531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  nor _46279_ (_02532_, _02514_, _02531_);
  or _46280_ (_37253_, _02532_, _02530_);
  and _46281_ (_02533_, _02514_, _35842_);
  not _46282_ (_02534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  nor _46283_ (_02535_, _02514_, _02534_);
  or _46284_ (_37254_, _02535_, _02533_);
  and _46285_ (_02536_, _02514_, _35846_);
  not _46286_ (_02537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  nor _46287_ (_02538_, _02514_, _02537_);
  or _46288_ (_37255_, _02538_, _02536_);
  and _46289_ (_02539_, _02313_, _36036_);
  and _46290_ (_02540_, _02539_, _35815_);
  not _46291_ (_02541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  nor _46292_ (_02542_, _02539_, _02541_);
  or _46293_ (_37256_, _02542_, _02540_);
  and _46294_ (_02543_, _02539_, _35822_);
  not _46295_ (_02544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  nor _46296_ (_02545_, _02539_, _02544_);
  or _46297_ (_37257_, _02545_, _02543_);
  and _46298_ (_02546_, _02539_, _35826_);
  not _46299_ (_02547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  nor _46300_ (_02548_, _02539_, _02547_);
  or _46301_ (_37258_, _02548_, _02546_);
  and _46302_ (_02549_, _02539_, _35830_);
  not _46303_ (_02550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  nor _46304_ (_02551_, _02539_, _02550_);
  or _46305_ (_37259_, _02551_, _02549_);
  and _46306_ (_02552_, _02539_, _35834_);
  not _46307_ (_02553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  nor _46308_ (_02554_, _02539_, _02553_);
  or _46309_ (_37260_, _02554_, _02552_);
  and _46310_ (_02555_, _02539_, _35838_);
  not _46311_ (_02556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  nor _46312_ (_02557_, _02539_, _02556_);
  or _46313_ (_37261_, _02557_, _02555_);
  and _46314_ (_02558_, _02539_, _35842_);
  not _46315_ (_02559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  nor _46316_ (_02560_, _02539_, _02559_);
  or _46317_ (_37262_, _02560_, _02558_);
  and _46318_ (_02561_, _02539_, _35846_);
  not _46319_ (_02562_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  nor _46320_ (_02563_, _02539_, _02562_);
  or _46321_ (_37263_, _02563_, _02561_);
  and _46322_ (_02564_, _02313_, _36062_);
  and _46323_ (_02565_, _02564_, _35815_);
  not _46324_ (_02566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  nor _46325_ (_02567_, _02564_, _02566_);
  or _46326_ (_37264_, _02567_, _02565_);
  and _46327_ (_02568_, _02564_, _35822_);
  not _46328_ (_02569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  nor _46329_ (_02570_, _02564_, _02569_);
  or _46330_ (_37265_, _02570_, _02568_);
  and _46331_ (_02571_, _02564_, _35826_);
  not _46332_ (_02572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  nor _46333_ (_02573_, _02564_, _02572_);
  or _46334_ (_37266_, _02573_, _02571_);
  and _46335_ (_02574_, _02564_, _35830_);
  not _46336_ (_02575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  nor _46337_ (_02576_, _02564_, _02575_);
  or _46338_ (_37267_, _02576_, _02574_);
  and _46339_ (_02577_, _02564_, _35834_);
  not _46340_ (_02578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  nor _46341_ (_02579_, _02564_, _02578_);
  or _46342_ (_37268_, _02579_, _02577_);
  and _46343_ (_02580_, _02564_, _35838_);
  not _46344_ (_02581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  nor _46345_ (_02582_, _02564_, _02581_);
  or _46346_ (_37269_, _02582_, _02580_);
  and _46347_ (_02583_, _02564_, _35842_);
  not _46348_ (_02584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  nor _46349_ (_02585_, _02564_, _02584_);
  or _46350_ (_37270_, _02585_, _02583_);
  and _46351_ (_02586_, _02564_, _35846_);
  not _46352_ (_02587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  nor _46353_ (_02588_, _02564_, _02587_);
  or _46354_ (_37271_, _02588_, _02586_);
  and _46355_ (_02589_, _02313_, _36088_);
  and _46356_ (_02590_, _02589_, _35815_);
  not _46357_ (_02591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  nor _46358_ (_02592_, _02589_, _02591_);
  or _46359_ (_37272_, _02592_, _02590_);
  and _46360_ (_02593_, _02589_, _35822_);
  not _46361_ (_02594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  nor _46362_ (_02595_, _02589_, _02594_);
  or _46363_ (_37273_, _02595_, _02593_);
  and _46364_ (_02596_, _02589_, _35826_);
  not _46365_ (_02597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  nor _46366_ (_02598_, _02589_, _02597_);
  or _46367_ (_37274_, _02598_, _02596_);
  and _46368_ (_02599_, _02589_, _35830_);
  not _46369_ (_02600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  nor _46370_ (_02601_, _02589_, _02600_);
  or _46371_ (_37275_, _02601_, _02599_);
  and _46372_ (_02602_, _02589_, _35834_);
  not _46373_ (_02603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  nor _46374_ (_02604_, _02589_, _02603_);
  or _46375_ (_37276_, _02604_, _02602_);
  and _46376_ (_02605_, _02589_, _35838_);
  not _46377_ (_02606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  nor _46378_ (_02607_, _02589_, _02606_);
  or _46379_ (_37277_, _02607_, _02605_);
  and _46380_ (_02608_, _02589_, _35842_);
  not _46381_ (_02609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  nor _46382_ (_02610_, _02589_, _02609_);
  or _46383_ (_37278_, _02610_, _02608_);
  and _46384_ (_02611_, _02589_, _35846_);
  not _46385_ (_02612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  nor _46386_ (_02613_, _02589_, _02612_);
  or _46387_ (_37279_, _02613_, _02611_);
  and _46388_ (_02614_, _02313_, _36115_);
  and _46389_ (_02615_, _02614_, _35815_);
  not _46390_ (_02616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  nor _46391_ (_02617_, _02614_, _02616_);
  or _46392_ (_37288_, _02617_, _02615_);
  and _46393_ (_02618_, _02614_, _35822_);
  not _46394_ (_02619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  nor _46395_ (_02620_, _02614_, _02619_);
  or _46396_ (_37289_, _02620_, _02618_);
  and _46397_ (_02621_, _02614_, _35826_);
  not _46398_ (_02622_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  nor _46399_ (_02623_, _02614_, _02622_);
  or _46400_ (_37290_, _02623_, _02621_);
  and _46401_ (_02624_, _02614_, _35830_);
  not _46402_ (_02625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  nor _46403_ (_02626_, _02614_, _02625_);
  or _46404_ (_37291_, _02626_, _02624_);
  and _46405_ (_02627_, _02614_, _35834_);
  not _46406_ (_02628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  nor _46407_ (_02629_, _02614_, _02628_);
  or _46408_ (_37292_, _02629_, _02627_);
  and _46409_ (_02630_, _02614_, _35838_);
  not _46410_ (_02631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  nor _46411_ (_02632_, _02614_, _02631_);
  or _46412_ (_37293_, _02632_, _02630_);
  and _46413_ (_02633_, _02614_, _35842_);
  not _46414_ (_02634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  nor _46415_ (_02635_, _02614_, _02634_);
  or _46416_ (_37294_, _02635_, _02633_);
  and _46417_ (_02636_, _02614_, _35846_);
  not _46418_ (_02637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  nor _46419_ (_02638_, _02614_, _02637_);
  or _46420_ (_37295_, _02638_, _02636_);
  and _46421_ (_02639_, _02313_, _36141_);
  and _46422_ (_02640_, _02639_, _35815_);
  not _46423_ (_02641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  nor _46424_ (_02642_, _02639_, _02641_);
  or _46425_ (_37296_, _02642_, _02640_);
  and _46426_ (_02643_, _02639_, _35822_);
  not _46427_ (_02644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  nor _46428_ (_02645_, _02639_, _02644_);
  or _46429_ (_37297_, _02645_, _02643_);
  and _46430_ (_02646_, _02639_, _35826_);
  not _46431_ (_02647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  nor _46432_ (_02648_, _02639_, _02647_);
  or _46433_ (_37298_, _02648_, _02646_);
  and _46434_ (_02649_, _02639_, _35830_);
  not _46435_ (_02650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  nor _46436_ (_02651_, _02639_, _02650_);
  or _46437_ (_37299_, _02651_, _02649_);
  and _46438_ (_02652_, _02639_, _35834_);
  not _46439_ (_02653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  nor _46440_ (_02654_, _02639_, _02653_);
  or _46441_ (_37300_, _02654_, _02652_);
  and _46442_ (_02655_, _02639_, _35838_);
  not _46443_ (_02656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  nor _46444_ (_02657_, _02639_, _02656_);
  or _46445_ (_37301_, _02657_, _02655_);
  and _46446_ (_02658_, _02639_, _35842_);
  not _46447_ (_02659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  nor _46448_ (_02660_, _02639_, _02659_);
  or _46449_ (_37302_, _02660_, _02658_);
  and _46450_ (_02661_, _02639_, _35846_);
  not _46451_ (_02662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  nor _46452_ (_02663_, _02639_, _02662_);
  or _46453_ (_37303_, _02663_, _02661_);
  and _46454_ (_02664_, _02313_, _36167_);
  and _46455_ (_02665_, _02664_, _35815_);
  not _46456_ (_02666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  nor _46457_ (_02667_, _02664_, _02666_);
  or _46458_ (_37304_, _02667_, _02665_);
  and _46459_ (_02668_, _02664_, _35822_);
  not _46460_ (_02669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  nor _46461_ (_02670_, _02664_, _02669_);
  or _46462_ (_37305_, _02670_, _02668_);
  and _46463_ (_02671_, _02664_, _35826_);
  not _46464_ (_02672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  nor _46465_ (_02673_, _02664_, _02672_);
  or _46466_ (_37306_, _02673_, _02671_);
  and _46467_ (_02674_, _02664_, _35830_);
  not _46468_ (_02675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  nor _46469_ (_02676_, _02664_, _02675_);
  or _46470_ (_37307_, _02676_, _02674_);
  and _46471_ (_02677_, _02664_, _35834_);
  not _46472_ (_02678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  nor _46473_ (_02679_, _02664_, _02678_);
  or _46474_ (_37308_, _02679_, _02677_);
  and _46475_ (_02680_, _02664_, _35838_);
  not _46476_ (_02681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  nor _46477_ (_02682_, _02664_, _02681_);
  or _46478_ (_37309_, _02682_, _02680_);
  and _46479_ (_02683_, _02664_, _35842_);
  not _46480_ (_02684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  nor _46481_ (_02685_, _02664_, _02684_);
  or _46482_ (_37310_, _02685_, _02683_);
  and _46483_ (_02686_, _02664_, _35846_);
  not _46484_ (_02687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  nor _46485_ (_02688_, _02664_, _02687_);
  or _46486_ (_37311_, _02688_, _02686_);
  and _46487_ (_02689_, _02313_, _36193_);
  and _46488_ (_02690_, _02689_, _35815_);
  not _46489_ (_02691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  nor _46490_ (_02692_, _02689_, _02691_);
  or _46491_ (_37312_, _02692_, _02690_);
  and _46492_ (_02693_, _02689_, _35822_);
  not _46493_ (_02694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  nor _46494_ (_02695_, _02689_, _02694_);
  or _46495_ (_37313_, _02695_, _02693_);
  and _46496_ (_02696_, _02689_, _35826_);
  not _46497_ (_02697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  nor _46498_ (_02698_, _02689_, _02697_);
  or _46499_ (_37314_, _02698_, _02696_);
  and _46500_ (_02699_, _02689_, _35830_);
  not _46501_ (_02700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  nor _46502_ (_02701_, _02689_, _02700_);
  or _46503_ (_37315_, _02701_, _02699_);
  and _46504_ (_02702_, _02689_, _35834_);
  not _46505_ (_02703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  nor _46506_ (_02704_, _02689_, _02703_);
  or _46507_ (_37316_, _02704_, _02702_);
  and _46508_ (_02705_, _02689_, _35838_);
  not _46509_ (_02706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  nor _46510_ (_02707_, _02689_, _02706_);
  or _46511_ (_37317_, _02707_, _02705_);
  and _46512_ (_02708_, _02689_, _35842_);
  not _46513_ (_02709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  nor _46514_ (_02710_, _02689_, _02709_);
  or _46515_ (_37318_, _02710_, _02708_);
  and _46516_ (_02711_, _02689_, _35846_);
  not _46517_ (_02712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  nor _46518_ (_02713_, _02689_, _02712_);
  or _46519_ (_37319_, _02713_, _02711_);
  and _46520_ (_02714_, _36220_, _33632_);
  and _46521_ (_02715_, _02714_, _35572_);
  and _46522_ (_02716_, _02715_, _35815_);
  not _46523_ (_02717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  nor _46524_ (_02718_, _02715_, _02717_);
  or _46525_ (_37320_, _02718_, _02716_);
  and _46526_ (_02719_, _02715_, _35822_);
  not _46527_ (_02720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  nor _46528_ (_02721_, _02715_, _02720_);
  or _46529_ (_37321_, _02721_, _02719_);
  and _46530_ (_02722_, _02715_, _35826_);
  not _46531_ (_02723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  nor _46532_ (_02724_, _02715_, _02723_);
  or _46533_ (_37322_, _02724_, _02722_);
  and _46534_ (_02725_, _02715_, _35830_);
  not _46535_ (_02726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  nor _46536_ (_02727_, _02715_, _02726_);
  or _46537_ (_37323_, _02727_, _02725_);
  and _46538_ (_02728_, _02715_, _35834_);
  not _46539_ (_02729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  nor _46540_ (_02730_, _02715_, _02729_);
  or _46541_ (_37324_, _02730_, _02728_);
  and _46542_ (_02731_, _02715_, _35838_);
  not _46543_ (_02732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  nor _46544_ (_02733_, _02715_, _02732_);
  or _46545_ (_37325_, _02733_, _02731_);
  and _46546_ (_02734_, _02715_, _35842_);
  not _46547_ (_02735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  nor _46548_ (_02736_, _02715_, _02735_);
  or _46549_ (_37326_, _02736_, _02734_);
  and _46550_ (_02737_, _02715_, _35846_);
  not _46551_ (_02738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  nor _46552_ (_02739_, _02715_, _02738_);
  or _46553_ (_37327_, _02739_, _02737_);
  and _46554_ (_02740_, _02714_, _35817_);
  and _46555_ (_02741_, _02740_, _35815_);
  not _46556_ (_02742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  nor _46557_ (_02743_, _02740_, _02742_);
  or _46558_ (_37328_, _02743_, _02741_);
  and _46559_ (_02744_, _02740_, _35822_);
  not _46560_ (_02745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  nor _46561_ (_02746_, _02740_, _02745_);
  or _46562_ (_37329_, _02746_, _02744_);
  and _46563_ (_02747_, _02740_, _35826_);
  not _46564_ (_02748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  nor _46565_ (_02749_, _02740_, _02748_);
  or _46566_ (_37330_, _02749_, _02747_);
  and _46567_ (_02750_, _02740_, _35830_);
  not _46568_ (_02751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  nor _46569_ (_02752_, _02740_, _02751_);
  or _46570_ (_37331_, _02752_, _02750_);
  and _46571_ (_02753_, _02740_, _35834_);
  not _46572_ (_02754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  nor _46573_ (_02755_, _02740_, _02754_);
  or _46574_ (_37332_, _02755_, _02753_);
  and _46575_ (_02756_, _02740_, _35838_);
  not _46576_ (_02757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  nor _46577_ (_02758_, _02740_, _02757_);
  or _46578_ (_37333_, _02758_, _02756_);
  and _46579_ (_02759_, _02740_, _35842_);
  not _46580_ (_02760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  nor _46581_ (_02761_, _02740_, _02760_);
  or _46582_ (_37334_, _02761_, _02759_);
  and _46583_ (_02762_, _02740_, _35846_);
  not _46584_ (_02763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  nor _46585_ (_02764_, _02740_, _02763_);
  or _46586_ (_37335_, _02764_, _02762_);
  and _46587_ (_02765_, _02714_, _35851_);
  and _46588_ (_02766_, _02765_, _35815_);
  not _46589_ (_02767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  nor _46590_ (_02768_, _02765_, _02767_);
  or _46591_ (_37336_, _02768_, _02766_);
  and _46592_ (_02769_, _02765_, _35822_);
  not _46593_ (_02770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  nor _46594_ (_02771_, _02765_, _02770_);
  or _46595_ (_37337_, _02771_, _02769_);
  and _46596_ (_02772_, _02765_, _35826_);
  not _46597_ (_02773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  nor _46598_ (_02774_, _02765_, _02773_);
  or _46599_ (_37338_, _02774_, _02772_);
  and _46600_ (_02775_, _02765_, _35830_);
  not _46601_ (_02776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  nor _46602_ (_02777_, _02765_, _02776_);
  or _46603_ (_37339_, _02777_, _02775_);
  and _46604_ (_02778_, _02765_, _35834_);
  not _46605_ (_02779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  nor _46606_ (_02780_, _02765_, _02779_);
  or _46607_ (_37340_, _02780_, _02778_);
  and _46608_ (_02781_, _02765_, _35838_);
  not _46609_ (_02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  nor _46610_ (_02783_, _02765_, _02782_);
  or _46611_ (_37341_, _02783_, _02781_);
  and _46612_ (_02784_, _02765_, _35842_);
  not _46613_ (_02785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  nor _46614_ (_02786_, _02765_, _02785_);
  or _46615_ (_37342_, _02786_, _02784_);
  and _46616_ (_02787_, _02765_, _35846_);
  not _46617_ (_02788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  nor _46618_ (_02789_, _02765_, _02788_);
  or _46619_ (_37343_, _02789_, _02787_);
  and _46620_ (_02790_, _02714_, _35878_);
  and _46621_ (_02791_, _02790_, _35815_);
  not _46622_ (_02792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  nor _46623_ (_02793_, _02790_, _02792_);
  or _46624_ (_37344_, _02793_, _02791_);
  and _46625_ (_02794_, _02790_, _35822_);
  not _46626_ (_02795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  nor _46627_ (_02796_, _02790_, _02795_);
  or _46628_ (_37345_, _02796_, _02794_);
  and _46629_ (_02797_, _02790_, _35826_);
  not _46630_ (_02798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  nor _46631_ (_02799_, _02790_, _02798_);
  or _46632_ (_37346_, _02799_, _02797_);
  and _46633_ (_02800_, _02790_, _35830_);
  not _46634_ (_02801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  nor _46635_ (_02802_, _02790_, _02801_);
  or _46636_ (_37347_, _02802_, _02800_);
  and _46637_ (_02803_, _02790_, _35834_);
  not _46638_ (_02804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  nor _46639_ (_02805_, _02790_, _02804_);
  or _46640_ (_37348_, _02805_, _02803_);
  and _46641_ (_02806_, _02790_, _35838_);
  not _46642_ (_02807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  nor _46643_ (_02808_, _02790_, _02807_);
  or _46644_ (_37349_, _02808_, _02806_);
  and _46645_ (_02809_, _02790_, _35842_);
  not _46646_ (_02810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  nor _46647_ (_02811_, _02790_, _02810_);
  or _46648_ (_37350_, _02811_, _02809_);
  and _46649_ (_02812_, _02790_, _35846_);
  not _46650_ (_02813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  nor _46651_ (_02814_, _02790_, _02813_);
  or _46652_ (_37351_, _02814_, _02812_);
  and _46653_ (_02815_, _02714_, _35905_);
  and _46654_ (_02816_, _02815_, _35815_);
  not _46655_ (_02817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  nor _46656_ (_02818_, _02815_, _02817_);
  or _46657_ (_37352_, _02818_, _02816_);
  and _46658_ (_02819_, _02815_, _35822_);
  not _46659_ (_02820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  nor _46660_ (_02821_, _02815_, _02820_);
  or _46661_ (_37353_, _02821_, _02819_);
  and _46662_ (_02822_, _02815_, _35826_);
  not _46663_ (_02823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  nor _46664_ (_02824_, _02815_, _02823_);
  or _46665_ (_37354_, _02824_, _02822_);
  and _46666_ (_02825_, _02815_, _35830_);
  not _46667_ (_02826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  nor _46668_ (_02827_, _02815_, _02826_);
  or _46669_ (_37355_, _02827_, _02825_);
  and _46670_ (_02828_, _02815_, _35834_);
  not _46671_ (_02829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  nor _46672_ (_02830_, _02815_, _02829_);
  or _46673_ (_37356_, _02830_, _02828_);
  and _46674_ (_02831_, _02815_, _35838_);
  not _46675_ (_02832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  nor _46676_ (_02833_, _02815_, _02832_);
  or _46677_ (_37357_, _02833_, _02831_);
  and _46678_ (_02834_, _02815_, _35842_);
  not _46679_ (_02835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  nor _46680_ (_02836_, _02815_, _02835_);
  or _46681_ (_37358_, _02836_, _02834_);
  and _46682_ (_02837_, _02815_, _35846_);
  not _46683_ (_02838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  nor _46684_ (_02839_, _02815_, _02838_);
  or _46685_ (_37359_, _02839_, _02837_);
  and _46686_ (_02840_, _02714_, _35931_);
  and _46687_ (_02841_, _02840_, _35815_);
  not _46688_ (_02842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  nor _46689_ (_02843_, _02840_, _02842_);
  or _46690_ (_37360_, _02843_, _02841_);
  and _46691_ (_02844_, _02840_, _35822_);
  not _46692_ (_02845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  nor _46693_ (_02846_, _02840_, _02845_);
  or _46694_ (_37361_, _02846_, _02844_);
  and _46695_ (_02847_, _02840_, _35826_);
  not _46696_ (_02848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  nor _46697_ (_02849_, _02840_, _02848_);
  or _46698_ (_37362_, _02849_, _02847_);
  and _46699_ (_02850_, _02840_, _35830_);
  not _46700_ (_02851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  nor _46701_ (_02852_, _02840_, _02851_);
  or _46702_ (_37363_, _02852_, _02850_);
  and _46703_ (_02853_, _02840_, _35834_);
  not _46704_ (_02854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  nor _46705_ (_02855_, _02840_, _02854_);
  or _46706_ (_37364_, _02855_, _02853_);
  and _46707_ (_02856_, _02840_, _35838_);
  not _46708_ (_02857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  nor _46709_ (_02858_, _02840_, _02857_);
  or _46710_ (_37365_, _02858_, _02856_);
  and _46711_ (_02859_, _02840_, _35842_);
  not _46712_ (_02860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  nor _46713_ (_02861_, _02840_, _02860_);
  or _46714_ (_37366_, _02861_, _02859_);
  and _46715_ (_02862_, _02840_, _35846_);
  not _46716_ (_02863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  nor _46717_ (_02864_, _02840_, _02863_);
  or _46718_ (_37367_, _02864_, _02862_);
  and _46719_ (_02865_, _02714_, _35957_);
  and _46720_ (_02866_, _02865_, _35815_);
  not _46721_ (_02867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  nor _46722_ (_02868_, _02865_, _02867_);
  or _46723_ (_37376_, _02868_, _02866_);
  and _46724_ (_02869_, _02865_, _35822_);
  not _46725_ (_02870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  nor _46726_ (_02871_, _02865_, _02870_);
  or _46727_ (_37377_, _02871_, _02869_);
  and _46728_ (_02872_, _02865_, _35826_);
  not _46729_ (_02873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  nor _46730_ (_02874_, _02865_, _02873_);
  or _46731_ (_37378_, _02874_, _02872_);
  and _46732_ (_02875_, _02865_, _35830_);
  not _46733_ (_02876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  nor _46734_ (_02877_, _02865_, _02876_);
  or _46735_ (_37379_, _02877_, _02875_);
  and _46736_ (_02878_, _02865_, _35834_);
  not _46737_ (_02879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  nor _46738_ (_02880_, _02865_, _02879_);
  or _46739_ (_37380_, _02880_, _02878_);
  and _46740_ (_02881_, _02865_, _35838_);
  not _46741_ (_02882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  nor _46742_ (_02883_, _02865_, _02882_);
  or _46743_ (_37381_, _02883_, _02881_);
  and _46744_ (_02884_, _02865_, _35842_);
  not _46745_ (_02885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  nor _46746_ (_02886_, _02865_, _02885_);
  or _46747_ (_37382_, _02886_, _02884_);
  and _46748_ (_02887_, _02865_, _35846_);
  not _46749_ (_02888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  nor _46750_ (_02889_, _02865_, _02888_);
  or _46751_ (_37383_, _02889_, _02887_);
  and _46752_ (_02890_, _02714_, _35983_);
  and _46753_ (_02891_, _02890_, _35815_);
  not _46754_ (_02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  nor _46755_ (_02893_, _02890_, _02892_);
  or _46756_ (_37384_, _02893_, _02891_);
  and _46757_ (_02894_, _02890_, _35822_);
  not _46758_ (_02895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  nor _46759_ (_02896_, _02890_, _02895_);
  or _46760_ (_37385_, _02896_, _02894_);
  and _46761_ (_02897_, _02890_, _35826_);
  not _46762_ (_02898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  nor _46763_ (_02899_, _02890_, _02898_);
  or _46764_ (_37386_, _02899_, _02897_);
  and _46765_ (_02900_, _02890_, _35830_);
  not _46766_ (_02901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  nor _46767_ (_02902_, _02890_, _02901_);
  or _46768_ (_37387_, _02902_, _02900_);
  and _46769_ (_02903_, _02890_, _35834_);
  not _46770_ (_02904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  nor _46771_ (_02905_, _02890_, _02904_);
  or _46772_ (_37388_, _02905_, _02903_);
  and _46773_ (_02906_, _02890_, _35838_);
  not _46774_ (_02907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  nor _46775_ (_02908_, _02890_, _02907_);
  or _46776_ (_37389_, _02908_, _02906_);
  and _46777_ (_02909_, _02890_, _35842_);
  not _46778_ (_02910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  nor _46779_ (_02911_, _02890_, _02910_);
  or _46780_ (_37390_, _02911_, _02909_);
  and _46781_ (_02912_, _02890_, _35846_);
  not _46782_ (_02913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  nor _46783_ (_02914_, _02890_, _02913_);
  or _46784_ (_37391_, _02914_, _02912_);
  and _46785_ (_02915_, _02714_, _36010_);
  and _46786_ (_02916_, _02915_, _35815_);
  not _46787_ (_02917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  nor _46788_ (_02918_, _02915_, _02917_);
  or _46789_ (_37392_, _02918_, _02916_);
  and _46790_ (_02919_, _02915_, _35822_);
  not _46791_ (_02920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  nor _46792_ (_02921_, _02915_, _02920_);
  or _46793_ (_37393_, _02921_, _02919_);
  and _46794_ (_02922_, _02915_, _35826_);
  not _46795_ (_02923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  nor _46796_ (_02924_, _02915_, _02923_);
  or _46797_ (_37394_, _02924_, _02922_);
  and _46798_ (_02925_, _02915_, _35830_);
  not _46799_ (_02926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  nor _46800_ (_02927_, _02915_, _02926_);
  or _46801_ (_37395_, _02927_, _02925_);
  and _46802_ (_02928_, _02915_, _35834_);
  not _46803_ (_02929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  nor _46804_ (_02930_, _02915_, _02929_);
  or _46805_ (_37396_, _02930_, _02928_);
  and _46806_ (_02931_, _02915_, _35838_);
  not _46807_ (_02932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  nor _46808_ (_02933_, _02915_, _02932_);
  or _46809_ (_37397_, _02933_, _02931_);
  and _46810_ (_02934_, _02915_, _35842_);
  not _46811_ (_02935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  nor _46812_ (_02936_, _02915_, _02935_);
  or _46813_ (_37398_, _02936_, _02934_);
  and _46814_ (_02937_, _02915_, _35846_);
  not _46815_ (_02938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  nor _46816_ (_02939_, _02915_, _02938_);
  or _46817_ (_37399_, _02939_, _02937_);
  and _46818_ (_02940_, _02714_, _36036_);
  and _46819_ (_02941_, _02940_, _35815_);
  not _46820_ (_02942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  nor _46821_ (_02943_, _02940_, _02942_);
  or _46822_ (_37400_, _02943_, _02941_);
  and _46823_ (_02944_, _02940_, _35822_);
  not _46824_ (_02945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  nor _46825_ (_02946_, _02940_, _02945_);
  or _46826_ (_37401_, _02946_, _02944_);
  and _46827_ (_02947_, _02940_, _35826_);
  not _46828_ (_02948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  nor _46829_ (_02949_, _02940_, _02948_);
  or _46830_ (_37402_, _02949_, _02947_);
  and _46831_ (_02950_, _02940_, _35830_);
  not _46832_ (_02951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  nor _46833_ (_02952_, _02940_, _02951_);
  or _46834_ (_37403_, _02952_, _02950_);
  and _46835_ (_02953_, _02940_, _35834_);
  not _46836_ (_02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  nor _46837_ (_02955_, _02940_, _02954_);
  or _46838_ (_37404_, _02955_, _02953_);
  and _46839_ (_02956_, _02940_, _35838_);
  not _46840_ (_02957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  nor _46841_ (_02958_, _02940_, _02957_);
  or _46842_ (_37405_, _02958_, _02956_);
  and _46843_ (_02959_, _02940_, _35842_);
  not _46844_ (_02960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  nor _46845_ (_02961_, _02940_, _02960_);
  or _46846_ (_37406_, _02961_, _02959_);
  and _46847_ (_02962_, _02940_, _35846_);
  not _46848_ (_02963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  nor _46849_ (_02964_, _02940_, _02963_);
  or _46850_ (_37407_, _02964_, _02962_);
  and _46851_ (_02965_, _02714_, _36062_);
  and _46852_ (_02966_, _02965_, _35815_);
  not _46853_ (_02967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  nor _46854_ (_02968_, _02965_, _02967_);
  or _46855_ (_37408_, _02968_, _02966_);
  and _46856_ (_02969_, _02965_, _35822_);
  not _46857_ (_02970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  nor _46858_ (_02971_, _02965_, _02970_);
  or _46859_ (_37409_, _02971_, _02969_);
  and _46860_ (_02972_, _02965_, _35826_);
  not _46861_ (_02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  nor _46862_ (_02974_, _02965_, _02973_);
  or _46863_ (_37410_, _02974_, _02972_);
  and _46864_ (_02975_, _02965_, _35830_);
  not _46865_ (_02976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  nor _46866_ (_02977_, _02965_, _02976_);
  or _46867_ (_37411_, _02977_, _02975_);
  and _46868_ (_02978_, _02965_, _35834_);
  not _46869_ (_02979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  nor _46870_ (_02980_, _02965_, _02979_);
  or _46871_ (_37412_, _02980_, _02978_);
  and _46872_ (_02981_, _02965_, _35838_);
  not _46873_ (_02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  nor _46874_ (_02983_, _02965_, _02982_);
  or _46875_ (_37413_, _02983_, _02981_);
  and _46876_ (_02984_, _02965_, _35842_);
  not _46877_ (_02985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  nor _46878_ (_02986_, _02965_, _02985_);
  or _46879_ (_37414_, _02986_, _02984_);
  and _46880_ (_02987_, _02965_, _35846_);
  not _46881_ (_02988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  nor _46882_ (_02989_, _02965_, _02988_);
  or _46883_ (_37415_, _02989_, _02987_);
  and _46884_ (_02990_, _02714_, _36088_);
  and _46885_ (_02991_, _02990_, _35815_);
  not _46886_ (_02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  nor _46887_ (_02993_, _02990_, _02992_);
  or _46888_ (_37416_, _02993_, _02991_);
  and _46889_ (_02994_, _02990_, _35822_);
  not _46890_ (_02995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  nor _46891_ (_02996_, _02990_, _02995_);
  or _46892_ (_37417_, _02996_, _02994_);
  and _46893_ (_02997_, _02990_, _35826_);
  not _46894_ (_02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  nor _46895_ (_02999_, _02990_, _02998_);
  or _46896_ (_37418_, _02999_, _02997_);
  and _46897_ (_03000_, _02990_, _35830_);
  not _46898_ (_03001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  nor _46899_ (_03002_, _02990_, _03001_);
  or _46900_ (_37419_, _03002_, _03000_);
  and _46901_ (_03003_, _02990_, _35834_);
  not _46902_ (_03004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  nor _46903_ (_03005_, _02990_, _03004_);
  or _46904_ (_37420_, _03005_, _03003_);
  and _46905_ (_03006_, _02990_, _35838_);
  not _46906_ (_03007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  nor _46907_ (_03008_, _02990_, _03007_);
  or _46908_ (_37421_, _03008_, _03006_);
  and _46909_ (_03009_, _02990_, _35842_);
  not _46910_ (_03010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  nor _46911_ (_03011_, _02990_, _03010_);
  or _46912_ (_37422_, _03011_, _03009_);
  and _46913_ (_03012_, _02990_, _35846_);
  not _46914_ (_03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  nor _46915_ (_03014_, _02990_, _03013_);
  or _46916_ (_37423_, _03014_, _03012_);
  and _46917_ (_03015_, _02714_, _36115_);
  and _46918_ (_03016_, _03015_, _35815_);
  not _46919_ (_03017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  nor _46920_ (_03018_, _03015_, _03017_);
  or _46921_ (_37424_, _03018_, _03016_);
  and _46922_ (_03019_, _03015_, _35822_);
  not _46923_ (_03020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  nor _46924_ (_03021_, _03015_, _03020_);
  or _46925_ (_37425_, _03021_, _03019_);
  and _46926_ (_03022_, _03015_, _35826_);
  not _46927_ (_03023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  nor _46928_ (_03024_, _03015_, _03023_);
  or _46929_ (_37426_, _03024_, _03022_);
  and _46930_ (_03025_, _03015_, _35830_);
  not _46931_ (_03026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  nor _46932_ (_03027_, _03015_, _03026_);
  or _46933_ (_37427_, _03027_, _03025_);
  and _46934_ (_03028_, _03015_, _35834_);
  not _46935_ (_03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  nor _46936_ (_03030_, _03015_, _03029_);
  or _46937_ (_37428_, _03030_, _03028_);
  and _46938_ (_03031_, _03015_, _35838_);
  not _46939_ (_03032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  nor _46940_ (_03033_, _03015_, _03032_);
  or _46941_ (_37429_, _03033_, _03031_);
  and _46942_ (_03034_, _03015_, _35842_);
  not _46943_ (_03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  nor _46944_ (_03036_, _03015_, _03035_);
  or _46945_ (_37430_, _03036_, _03034_);
  and _46946_ (_03037_, _03015_, _35846_);
  not _46947_ (_03038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  nor _46948_ (_03039_, _03015_, _03038_);
  or _46949_ (_37431_, _03039_, _03037_);
  and _46950_ (_03040_, _02714_, _36141_);
  and _46951_ (_03041_, _03040_, _35815_);
  not _46952_ (_03042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  nor _46953_ (_03043_, _03040_, _03042_);
  or _46954_ (_37432_, _03043_, _03041_);
  and _46955_ (_03044_, _03040_, _35822_);
  not _46956_ (_03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  nor _46957_ (_03046_, _03040_, _03045_);
  or _46958_ (_37433_, _03046_, _03044_);
  and _46959_ (_03047_, _03040_, _35826_);
  not _46960_ (_03048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  nor _46961_ (_03049_, _03040_, _03048_);
  or _46962_ (_37434_, _03049_, _03047_);
  and _46963_ (_03050_, _03040_, _35830_);
  not _46964_ (_03051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  nor _46965_ (_03052_, _03040_, _03051_);
  or _46966_ (_37435_, _03052_, _03050_);
  and _46967_ (_03053_, _03040_, _35834_);
  not _46968_ (_03054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  nor _46969_ (_03055_, _03040_, _03054_);
  or _46970_ (_37436_, _03055_, _03053_);
  and _46971_ (_03056_, _03040_, _35838_);
  not _46972_ (_03057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  nor _46973_ (_03058_, _03040_, _03057_);
  or _46974_ (_37437_, _03058_, _03056_);
  and _46975_ (_03059_, _03040_, _35842_);
  not _46976_ (_03060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  nor _46977_ (_03061_, _03040_, _03060_);
  or _46978_ (_37438_, _03061_, _03059_);
  and _46979_ (_03062_, _03040_, _35846_);
  not _46980_ (_03063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  nor _46981_ (_03064_, _03040_, _03063_);
  or _46982_ (_37439_, _03064_, _03062_);
  and _46983_ (_03065_, _02714_, _36167_);
  and _46984_ (_03066_, _03065_, _35815_);
  not _46985_ (_03067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  nor _46986_ (_03068_, _03065_, _03067_);
  or _46987_ (_37440_, _03068_, _03066_);
  and _46988_ (_03069_, _03065_, _35822_);
  not _46989_ (_03070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  nor _46990_ (_03071_, _03065_, _03070_);
  or _46991_ (_37441_, _03071_, _03069_);
  and _46992_ (_03072_, _03065_, _35826_);
  not _46993_ (_03073_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  nor _46994_ (_03074_, _03065_, _03073_);
  or _46995_ (_37442_, _03074_, _03072_);
  and _46996_ (_03075_, _03065_, _35830_);
  not _46997_ (_03076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  nor _46998_ (_03077_, _03065_, _03076_);
  or _46999_ (_37443_, _03077_, _03075_);
  and _47000_ (_03078_, _03065_, _35834_);
  not _47001_ (_03079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  nor _47002_ (_03080_, _03065_, _03079_);
  or _47003_ (_37444_, _03080_, _03078_);
  and _47004_ (_03081_, _03065_, _35838_);
  not _47005_ (_03082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  nor _47006_ (_03083_, _03065_, _03082_);
  or _47007_ (_37445_, _03083_, _03081_);
  and _47008_ (_03084_, _03065_, _35842_);
  not _47009_ (_03085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  nor _47010_ (_03086_, _03065_, _03085_);
  or _47011_ (_37446_, _03086_, _03084_);
  and _47012_ (_03087_, _03065_, _35846_);
  not _47013_ (_03088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  nor _47014_ (_03089_, _03065_, _03088_);
  or _47015_ (_37447_, _03089_, _03087_);
  and _47016_ (_03090_, _02714_, _36193_);
  and _47017_ (_03091_, _03090_, _35815_);
  not _47018_ (_03092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  nor _47019_ (_03093_, _03090_, _03092_);
  or _47020_ (_37448_, _03093_, _03091_);
  and _47021_ (_03094_, _03090_, _35822_);
  not _47022_ (_03095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  nor _47023_ (_03096_, _03090_, _03095_);
  or _47024_ (_37449_, _03096_, _03094_);
  and _47025_ (_03097_, _03090_, _35826_);
  not _47026_ (_03098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  nor _47027_ (_03099_, _03090_, _03098_);
  or _47028_ (_37450_, _03099_, _03097_);
  and _47029_ (_03100_, _03090_, _35830_);
  not _47030_ (_03101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  nor _47031_ (_03102_, _03090_, _03101_);
  or _47032_ (_37451_, _03102_, _03100_);
  and _47033_ (_03103_, _03090_, _35834_);
  not _47034_ (_03104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  nor _47035_ (_03105_, _03090_, _03104_);
  or _47036_ (_37452_, _03105_, _03103_);
  and _47037_ (_03106_, _03090_, _35838_);
  not _47038_ (_03107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  nor _47039_ (_03108_, _03090_, _03107_);
  or _47040_ (_37453_, _03108_, _03106_);
  and _47041_ (_03109_, _03090_, _35842_);
  not _47042_ (_03110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  nor _47043_ (_03111_, _03090_, _03110_);
  or _47044_ (_37454_, _03111_, _03109_);
  and _47045_ (_03112_, _03090_, _35846_);
  not _47046_ (_03113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  nor _47047_ (_03114_, _03090_, _03113_);
  or _47048_ (_37455_, _03114_, _03112_);
  not _47049_ (_03115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  and _47050_ (_03116_, _02312_, _36622_);
  and _47051_ (_03117_, _03116_, _35572_);
  nor _47052_ (_03118_, _03117_, _03115_);
  and _47053_ (_03119_, _03117_, _35815_);
  or _47054_ (_37464_, _03119_, _03118_);
  not _47055_ (_03120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  nor _47056_ (_03121_, _03117_, _03120_);
  and _47057_ (_03122_, _03117_, _35822_);
  or _47058_ (_37465_, _03122_, _03121_);
  not _47059_ (_03123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  nor _47060_ (_03124_, _03117_, _03123_);
  and _47061_ (_03125_, _03117_, _35826_);
  or _47062_ (_37466_, _03125_, _03124_);
  not _47063_ (_03126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  nor _47064_ (_03127_, _03117_, _03126_);
  and _47065_ (_03128_, _03117_, _35830_);
  or _47066_ (_37467_, _03128_, _03127_);
  not _47067_ (_03129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  nor _47068_ (_03130_, _03117_, _03129_);
  and _47069_ (_03131_, _03117_, _35834_);
  or _47070_ (_37468_, _03131_, _03130_);
  not _47071_ (_03132_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  nor _47072_ (_03133_, _03117_, _03132_);
  and _47073_ (_03134_, _03117_, _35838_);
  or _47074_ (_37469_, _03134_, _03133_);
  not _47075_ (_03135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  nor _47076_ (_03136_, _03117_, _03135_);
  and _47077_ (_03137_, _03117_, _35842_);
  or _47078_ (_37470_, _03137_, _03136_);
  not _47079_ (_03138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  nor _47080_ (_03139_, _03117_, _03138_);
  and _47081_ (_03140_, _03117_, _35846_);
  or _47082_ (_37471_, _03140_, _03139_);
  not _47083_ (_03141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and _47084_ (_03142_, _03116_, _35817_);
  nor _47085_ (_03143_, _03142_, _03141_);
  and _47086_ (_03144_, _03142_, _35815_);
  or _47087_ (_37472_, _03144_, _03143_);
  not _47088_ (_03145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  nor _47089_ (_03146_, _03142_, _03145_);
  and _47090_ (_03147_, _03142_, _35822_);
  or _47091_ (_37473_, _03147_, _03146_);
  not _47092_ (_03148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  nor _47093_ (_03149_, _03142_, _03148_);
  and _47094_ (_03150_, _03142_, _35826_);
  or _47095_ (_37474_, _03150_, _03149_);
  not _47096_ (_03151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  nor _47097_ (_03152_, _03142_, _03151_);
  and _47098_ (_03153_, _03142_, _35830_);
  or _47099_ (_37475_, _03153_, _03152_);
  not _47100_ (_03154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  nor _47101_ (_03155_, _03142_, _03154_);
  and _47102_ (_03156_, _03142_, _35834_);
  or _47103_ (_37476_, _03156_, _03155_);
  not _47104_ (_03157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  nor _47105_ (_03158_, _03142_, _03157_);
  and _47106_ (_03159_, _03142_, _35838_);
  or _47107_ (_37477_, _03159_, _03158_);
  not _47108_ (_03160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  nor _47109_ (_03161_, _03142_, _03160_);
  and _47110_ (_03162_, _03142_, _35842_);
  or _47111_ (_37478_, _03162_, _03161_);
  not _47112_ (_03163_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  nor _47113_ (_03164_, _03142_, _03163_);
  and _47114_ (_03165_, _03142_, _35846_);
  or _47115_ (_37479_, _03165_, _03164_);
  not _47116_ (_03166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and _47117_ (_03167_, _03116_, _35851_);
  nor _47118_ (_03168_, _03167_, _03166_);
  and _47119_ (_03169_, _03167_, _35815_);
  or _47120_ (_37480_, _03169_, _03168_);
  not _47121_ (_03170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  nor _47122_ (_03171_, _03167_, _03170_);
  and _47123_ (_03172_, _03167_, _35822_);
  or _47124_ (_37481_, _03172_, _03171_);
  not _47125_ (_03173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  nor _47126_ (_03174_, _03167_, _03173_);
  and _47127_ (_03175_, _03167_, _35826_);
  or _47128_ (_37482_, _03175_, _03174_);
  not _47129_ (_03176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  nor _47130_ (_03177_, _03167_, _03176_);
  and _47131_ (_03178_, _03167_, _35830_);
  or _47132_ (_37483_, _03178_, _03177_);
  not _47133_ (_03179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  nor _47134_ (_03180_, _03167_, _03179_);
  and _47135_ (_03181_, _03167_, _35834_);
  or _47136_ (_37484_, _03181_, _03180_);
  not _47137_ (_03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  nor _47138_ (_03183_, _03167_, _03182_);
  and _47139_ (_03184_, _03167_, _35838_);
  or _47140_ (_37485_, _03184_, _03183_);
  not _47141_ (_03185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  nor _47142_ (_03186_, _03167_, _03185_);
  and _47143_ (_03187_, _03167_, _35842_);
  or _47144_ (_37486_, _03187_, _03186_);
  not _47145_ (_03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  nor _47146_ (_03189_, _03167_, _03188_);
  and _47147_ (_03190_, _03167_, _35846_);
  or _47148_ (_37487_, _03190_, _03189_);
  not _47149_ (_03191_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  and _47150_ (_03192_, _03116_, _35878_);
  nor _47151_ (_03193_, _03192_, _03191_);
  and _47152_ (_03194_, _03192_, _35815_);
  or _47153_ (_37488_, _03194_, _03193_);
  not _47154_ (_03195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  nor _47155_ (_03196_, _03192_, _03195_);
  and _47156_ (_03197_, _03192_, _35822_);
  or _47157_ (_37489_, _03197_, _03196_);
  not _47158_ (_03198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  nor _47159_ (_03199_, _03192_, _03198_);
  and _47160_ (_03200_, _03192_, _35826_);
  or _47161_ (_37490_, _03200_, _03199_);
  not _47162_ (_03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  nor _47163_ (_03202_, _03192_, _03201_);
  and _47164_ (_03203_, _03192_, _35830_);
  or _47165_ (_37491_, _03203_, _03202_);
  not _47166_ (_03204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  nor _47167_ (_03205_, _03192_, _03204_);
  and _47168_ (_03206_, _03192_, _35834_);
  or _47169_ (_37492_, _03206_, _03205_);
  not _47170_ (_03207_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  nor _47171_ (_03208_, _03192_, _03207_);
  and _47172_ (_03209_, _03192_, _35838_);
  or _47173_ (_37493_, _03209_, _03208_);
  not _47174_ (_03210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  nor _47175_ (_03211_, _03192_, _03210_);
  and _47176_ (_03212_, _03192_, _35842_);
  or _47177_ (_37494_, _03212_, _03211_);
  not _47178_ (_03213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  nor _47179_ (_03214_, _03192_, _03213_);
  and _47180_ (_03215_, _03192_, _35846_);
  or _47181_ (_37495_, _03215_, _03214_);
  not _47182_ (_03216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and _47183_ (_03217_, _03116_, _35905_);
  nor _47184_ (_03218_, _03217_, _03216_);
  and _47185_ (_03219_, _03217_, _35815_);
  or _47186_ (_37496_, _03219_, _03218_);
  not _47187_ (_03220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  nor _47188_ (_03221_, _03217_, _03220_);
  and _47189_ (_03222_, _03217_, _35822_);
  or _47190_ (_37497_, _03222_, _03221_);
  not _47191_ (_03223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  nor _47192_ (_03224_, _03217_, _03223_);
  and _47193_ (_03225_, _03217_, _35826_);
  or _47194_ (_37498_, _03225_, _03224_);
  not _47195_ (_03226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  nor _47196_ (_03227_, _03217_, _03226_);
  and _47197_ (_03228_, _03217_, _35830_);
  or _47198_ (_37499_, _03228_, _03227_);
  not _47199_ (_03229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  nor _47200_ (_03230_, _03217_, _03229_);
  and _47201_ (_03231_, _03217_, _35834_);
  or _47202_ (_37500_, _03231_, _03230_);
  not _47203_ (_03232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  nor _47204_ (_03233_, _03217_, _03232_);
  and _47205_ (_03234_, _03217_, _35838_);
  or _47206_ (_37501_, _03234_, _03233_);
  not _47207_ (_03235_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  nor _47208_ (_03236_, _03217_, _03235_);
  and _47209_ (_03237_, _03217_, _35842_);
  or _47210_ (_37502_, _03237_, _03236_);
  not _47211_ (_03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  nor _47212_ (_03239_, _03217_, _03238_);
  and _47213_ (_03240_, _03217_, _35846_);
  or _47214_ (_37503_, _03240_, _03239_);
  not _47215_ (_03241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and _47216_ (_03242_, _03116_, _35931_);
  nor _47217_ (_03243_, _03242_, _03241_);
  and _47218_ (_03244_, _03242_, _35815_);
  or _47219_ (_37504_, _03244_, _03243_);
  not _47220_ (_03245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  nor _47221_ (_03246_, _03242_, _03245_);
  and _47222_ (_03247_, _03242_, _35822_);
  or _47223_ (_37505_, _03247_, _03246_);
  not _47224_ (_03248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  nor _47225_ (_03249_, _03242_, _03248_);
  and _47226_ (_03250_, _03242_, _35826_);
  or _47227_ (_37506_, _03250_, _03249_);
  not _47228_ (_03251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  nor _47229_ (_03252_, _03242_, _03251_);
  and _47230_ (_03253_, _03242_, _35830_);
  or _47231_ (_37507_, _03253_, _03252_);
  not _47232_ (_03254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  nor _47233_ (_03255_, _03242_, _03254_);
  and _47234_ (_03256_, _03242_, _35834_);
  or _47235_ (_37508_, _03256_, _03255_);
  not _47236_ (_03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  nor _47237_ (_03258_, _03242_, _03257_);
  and _47238_ (_03259_, _03242_, _35838_);
  or _47239_ (_37509_, _03259_, _03258_);
  not _47240_ (_03260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  nor _47241_ (_03261_, _03242_, _03260_);
  and _47242_ (_03262_, _03242_, _35842_);
  or _47243_ (_37510_, _03262_, _03261_);
  not _47244_ (_03263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  nor _47245_ (_03264_, _03242_, _03263_);
  and _47246_ (_03265_, _03242_, _35846_);
  or _47247_ (_37511_, _03265_, _03264_);
  not _47248_ (_03266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and _47249_ (_03267_, _03116_, _35957_);
  nor _47250_ (_03268_, _03267_, _03266_);
  and _47251_ (_03269_, _03267_, _35815_);
  or _47252_ (_37512_, _03269_, _03268_);
  not _47253_ (_03270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  nor _47254_ (_03271_, _03267_, _03270_);
  and _47255_ (_03272_, _03267_, _35822_);
  or _47256_ (_37513_, _03272_, _03271_);
  not _47257_ (_03273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  nor _47258_ (_03274_, _03267_, _03273_);
  and _47259_ (_03275_, _03267_, _35826_);
  or _47260_ (_37514_, _03275_, _03274_);
  not _47261_ (_03276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  nor _47262_ (_03277_, _03267_, _03276_);
  and _47263_ (_03278_, _03267_, _35830_);
  or _47264_ (_37515_, _03278_, _03277_);
  not _47265_ (_03279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  nor _47266_ (_03280_, _03267_, _03279_);
  and _47267_ (_03281_, _03267_, _35834_);
  or _47268_ (_37516_, _03281_, _03280_);
  not _47269_ (_03282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  nor _47270_ (_03283_, _03267_, _03282_);
  and _47271_ (_03284_, _03267_, _35838_);
  or _47272_ (_37517_, _03284_, _03283_);
  not _47273_ (_03285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  nor _47274_ (_03286_, _03267_, _03285_);
  and _47275_ (_03287_, _03267_, _35842_);
  or _47276_ (_37518_, _03287_, _03286_);
  not _47277_ (_03288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  nor _47278_ (_03289_, _03267_, _03288_);
  and _47279_ (_03290_, _03267_, _35846_);
  or _47280_ (_37519_, _03290_, _03289_);
  not _47281_ (_03291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  and _47282_ (_03292_, _03116_, _35983_);
  nor _47283_ (_03293_, _03292_, _03291_);
  and _47284_ (_03294_, _03292_, _35815_);
  or _47285_ (_37520_, _03294_, _03293_);
  not _47286_ (_03295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  nor _47287_ (_03296_, _03292_, _03295_);
  and _47288_ (_03297_, _03292_, _35822_);
  or _47289_ (_37521_, _03297_, _03296_);
  not _47290_ (_03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  nor _47291_ (_03299_, _03292_, _03298_);
  and _47292_ (_03300_, _03292_, _35826_);
  or _47293_ (_37522_, _03300_, _03299_);
  not _47294_ (_03301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  nor _47295_ (_03302_, _03292_, _03301_);
  and _47296_ (_03303_, _03292_, _35830_);
  or _47297_ (_37523_, _03303_, _03302_);
  not _47298_ (_03304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  nor _47299_ (_03305_, _03292_, _03304_);
  and _47300_ (_03306_, _03292_, _35834_);
  or _47301_ (_37524_, _03306_, _03305_);
  not _47302_ (_03307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  nor _47303_ (_03308_, _03292_, _03307_);
  and _47304_ (_03309_, _03292_, _35838_);
  or _47305_ (_37525_, _03309_, _03308_);
  not _47306_ (_03310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  nor _47307_ (_03311_, _03292_, _03310_);
  and _47308_ (_03312_, _03292_, _35842_);
  or _47309_ (_37526_, _03312_, _03311_);
  not _47310_ (_03313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  nor _47311_ (_03314_, _03292_, _03313_);
  and _47312_ (_03315_, _03292_, _35846_);
  or _47313_ (_37527_, _03315_, _03314_);
  not _47314_ (_03316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and _47315_ (_03317_, _03116_, _36010_);
  nor _47316_ (_03318_, _03317_, _03316_);
  and _47317_ (_03319_, _03317_, _35815_);
  or _47318_ (_37528_, _03319_, _03318_);
  not _47319_ (_03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  nor _47320_ (_03321_, _03317_, _03320_);
  and _47321_ (_03322_, _03317_, _35822_);
  or _47322_ (_37529_, _03322_, _03321_);
  not _47323_ (_03323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  nor _47324_ (_03324_, _03317_, _03323_);
  and _47325_ (_03325_, _03317_, _35826_);
  or _47326_ (_37530_, _03325_, _03324_);
  not _47327_ (_03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  nor _47328_ (_03327_, _03317_, _03326_);
  and _47329_ (_03328_, _03317_, _35830_);
  or _47330_ (_37531_, _03328_, _03327_);
  not _47331_ (_03329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  nor _47332_ (_03330_, _03317_, _03329_);
  and _47333_ (_03331_, _03317_, _35834_);
  or _47334_ (_37532_, _03331_, _03330_);
  not _47335_ (_03332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  nor _47336_ (_03333_, _03317_, _03332_);
  and _47337_ (_03334_, _03317_, _35838_);
  or _47338_ (_37533_, _03334_, _03333_);
  not _47339_ (_03335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  nor _47340_ (_03336_, _03317_, _03335_);
  and _47341_ (_03337_, _03317_, _35842_);
  or _47342_ (_37534_, _03337_, _03336_);
  not _47343_ (_03338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  nor _47344_ (_03339_, _03317_, _03338_);
  and _47345_ (_03340_, _03317_, _35846_);
  or _47346_ (_37535_, _03340_, _03339_);
  not _47347_ (_03341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  and _47348_ (_03342_, _03116_, _36036_);
  nor _47349_ (_03343_, _03342_, _03341_);
  and _47350_ (_03344_, _03342_, _35815_);
  or _47351_ (_37536_, _03344_, _03343_);
  not _47352_ (_03345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  nor _47353_ (_03346_, _03342_, _03345_);
  and _47354_ (_03347_, _03342_, _35822_);
  or _47355_ (_37537_, _03347_, _03346_);
  not _47356_ (_03348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  nor _47357_ (_03349_, _03342_, _03348_);
  and _47358_ (_03350_, _03342_, _35826_);
  or _47359_ (_37538_, _03350_, _03349_);
  not _47360_ (_03351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  nor _47361_ (_03352_, _03342_, _03351_);
  and _47362_ (_03353_, _03342_, _35830_);
  or _47363_ (_37539_, _03353_, _03352_);
  not _47364_ (_03354_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  nor _47365_ (_03355_, _03342_, _03354_);
  and _47366_ (_03356_, _03342_, _35834_);
  or _47367_ (_37540_, _03356_, _03355_);
  not _47368_ (_03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  nor _47369_ (_03358_, _03342_, _03357_);
  and _47370_ (_03359_, _03342_, _35838_);
  or _47371_ (_37541_, _03359_, _03358_);
  not _47372_ (_03360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  nor _47373_ (_03361_, _03342_, _03360_);
  and _47374_ (_03362_, _03342_, _35842_);
  or _47375_ (_37542_, _03362_, _03361_);
  not _47376_ (_03363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  nor _47377_ (_03364_, _03342_, _03363_);
  and _47378_ (_03365_, _03342_, _35846_);
  or _47379_ (_37543_, _03365_, _03364_);
  not _47380_ (_03366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and _47381_ (_03367_, _03116_, _36062_);
  nor _47382_ (_03368_, _03367_, _03366_);
  and _47383_ (_03369_, _03367_, _35815_);
  or _47384_ (_37552_, _03369_, _03368_);
  not _47385_ (_03370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  nor _47386_ (_03371_, _03367_, _03370_);
  and _47387_ (_03372_, _03367_, _35822_);
  or _47388_ (_37553_, _03372_, _03371_);
  not _47389_ (_03373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  nor _47390_ (_03374_, _03367_, _03373_);
  and _47391_ (_03375_, _03367_, _35826_);
  or _47392_ (_37554_, _03375_, _03374_);
  not _47393_ (_03376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  nor _47394_ (_03377_, _03367_, _03376_);
  and _47395_ (_03378_, _03367_, _35830_);
  or _47396_ (_37555_, _03378_, _03377_);
  not _47397_ (_03379_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  nor _47398_ (_03380_, _03367_, _03379_);
  and _47399_ (_03381_, _03367_, _35834_);
  or _47400_ (_37556_, _03381_, _03380_);
  not _47401_ (_03382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  nor _47402_ (_03383_, _03367_, _03382_);
  and _47403_ (_03384_, _03367_, _35838_);
  or _47404_ (_37557_, _03384_, _03383_);
  not _47405_ (_03385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  nor _47406_ (_03386_, _03367_, _03385_);
  and _47407_ (_03387_, _03367_, _35842_);
  or _47408_ (_37558_, _03387_, _03386_);
  not _47409_ (_03388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  nor _47410_ (_03389_, _03367_, _03388_);
  and _47411_ (_03390_, _03367_, _35846_);
  or _47412_ (_37559_, _03390_, _03389_);
  not _47413_ (_03391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and _47414_ (_03392_, _03116_, _36088_);
  nor _47415_ (_03393_, _03392_, _03391_);
  and _47416_ (_03394_, _03392_, _35815_);
  or _47417_ (_37560_, _03394_, _03393_);
  not _47418_ (_03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  nor _47419_ (_03396_, _03392_, _03395_);
  and _47420_ (_03397_, _03392_, _35822_);
  or _47421_ (_37561_, _03397_, _03396_);
  not _47422_ (_03398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  nor _47423_ (_03399_, _03392_, _03398_);
  and _47424_ (_03400_, _03392_, _35826_);
  or _47425_ (_37562_, _03400_, _03399_);
  not _47426_ (_03401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  nor _47427_ (_03402_, _03392_, _03401_);
  and _47428_ (_03403_, _03392_, _35830_);
  or _47429_ (_37563_, _03403_, _03402_);
  not _47430_ (_03404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  nor _47431_ (_03405_, _03392_, _03404_);
  and _47432_ (_03406_, _03392_, _35834_);
  or _47433_ (_37564_, _03406_, _03405_);
  not _47434_ (_03407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  nor _47435_ (_03408_, _03392_, _03407_);
  and _47436_ (_03409_, _03392_, _35838_);
  or _47437_ (_37565_, _03409_, _03408_);
  not _47438_ (_03410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  nor _47439_ (_03411_, _03392_, _03410_);
  and _47440_ (_03412_, _03392_, _35842_);
  or _47441_ (_37566_, _03412_, _03411_);
  not _47442_ (_03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  nor _47443_ (_03414_, _03392_, _03413_);
  and _47444_ (_03415_, _03392_, _35846_);
  or _47445_ (_37567_, _03415_, _03414_);
  not _47446_ (_03416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and _47447_ (_03417_, _03116_, _36115_);
  nor _47448_ (_03418_, _03417_, _03416_);
  and _47449_ (_03419_, _03417_, _35815_);
  or _47450_ (_37568_, _03419_, _03418_);
  not _47451_ (_03420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  nor _47452_ (_03421_, _03417_, _03420_);
  and _47453_ (_03422_, _03417_, _35822_);
  or _47454_ (_37569_, _03422_, _03421_);
  not _47455_ (_03423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  nor _47456_ (_03424_, _03417_, _03423_);
  and _47457_ (_03425_, _03417_, _35826_);
  or _47458_ (_37570_, _03425_, _03424_);
  not _47459_ (_03426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  nor _47460_ (_03427_, _03417_, _03426_);
  and _47461_ (_03428_, _03417_, _35830_);
  or _47462_ (_37571_, _03428_, _03427_);
  not _47463_ (_03429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  nor _47464_ (_03430_, _03417_, _03429_);
  and _47465_ (_03431_, _03417_, _35834_);
  or _47466_ (_37572_, _03431_, _03430_);
  not _47467_ (_03432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  nor _47468_ (_03433_, _03417_, _03432_);
  and _47469_ (_03434_, _03417_, _35838_);
  or _47470_ (_37573_, _03434_, _03433_);
  not _47471_ (_03435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  nor _47472_ (_03436_, _03417_, _03435_);
  and _47473_ (_03437_, _03417_, _35842_);
  or _47474_ (_37574_, _03437_, _03436_);
  not _47475_ (_03438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  nor _47476_ (_03439_, _03417_, _03438_);
  and _47477_ (_03440_, _03417_, _35846_);
  or _47478_ (_37575_, _03440_, _03439_);
  not _47479_ (_03441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  and _47480_ (_03442_, _03116_, _36141_);
  nor _47481_ (_03443_, _03442_, _03441_);
  and _47482_ (_03444_, _03442_, _35815_);
  or _47483_ (_37576_, _03444_, _03443_);
  not _47484_ (_03445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  nor _47485_ (_03446_, _03442_, _03445_);
  and _47486_ (_03447_, _03442_, _35822_);
  or _47487_ (_37577_, _03447_, _03446_);
  not _47488_ (_03448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  nor _47489_ (_03449_, _03442_, _03448_);
  and _47490_ (_03450_, _03442_, _35826_);
  or _47491_ (_37578_, _03450_, _03449_);
  not _47492_ (_03451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  nor _47493_ (_03452_, _03442_, _03451_);
  and _47494_ (_03453_, _03442_, _35830_);
  or _47495_ (_37579_, _03453_, _03452_);
  not _47496_ (_03454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  nor _47497_ (_03455_, _03442_, _03454_);
  and _47498_ (_03456_, _03442_, _35834_);
  or _47499_ (_37580_, _03456_, _03455_);
  not _47500_ (_03457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  nor _47501_ (_03458_, _03442_, _03457_);
  and _47502_ (_03459_, _03442_, _35838_);
  or _47503_ (_37581_, _03459_, _03458_);
  not _47504_ (_03460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  nor _47505_ (_03461_, _03442_, _03460_);
  and _47506_ (_03462_, _03442_, _35842_);
  or _47507_ (_37582_, _03462_, _03461_);
  not _47508_ (_03463_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  nor _47509_ (_03464_, _03442_, _03463_);
  and _47510_ (_03465_, _03442_, _35846_);
  or _47511_ (_37583_, _03465_, _03464_);
  not _47512_ (_03466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  and _47513_ (_03467_, _03116_, _36167_);
  nor _47514_ (_03468_, _03467_, _03466_);
  and _47515_ (_03469_, _03467_, _35815_);
  or _47516_ (_37584_, _03469_, _03468_);
  not _47517_ (_03470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  nor _47518_ (_03471_, _03467_, _03470_);
  and _47519_ (_03472_, _03467_, _35822_);
  or _47520_ (_37585_, _03472_, _03471_);
  not _47521_ (_03473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  nor _47522_ (_03474_, _03467_, _03473_);
  and _47523_ (_03475_, _03467_, _35826_);
  or _47524_ (_37586_, _03475_, _03474_);
  not _47525_ (_03476_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  nor _47526_ (_03477_, _03467_, _03476_);
  and _47527_ (_03478_, _03467_, _35830_);
  or _47528_ (_37587_, _03478_, _03477_);
  not _47529_ (_03479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  nor _47530_ (_03480_, _03467_, _03479_);
  and _47531_ (_03481_, _03467_, _35834_);
  or _47532_ (_37588_, _03481_, _03480_);
  not _47533_ (_03482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  nor _47534_ (_03483_, _03467_, _03482_);
  and _47535_ (_03484_, _03467_, _35838_);
  or _47536_ (_37589_, _03484_, _03483_);
  not _47537_ (_03485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  nor _47538_ (_03486_, _03467_, _03485_);
  and _47539_ (_03487_, _03467_, _35842_);
  or _47540_ (_37590_, _03487_, _03486_);
  not _47541_ (_03488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  nor _47542_ (_03489_, _03467_, _03488_);
  and _47543_ (_03490_, _03467_, _35846_);
  or _47544_ (_37591_, _03490_, _03489_);
  not _47545_ (_03491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and _47546_ (_03492_, _03116_, _36193_);
  nor _47547_ (_03493_, _03492_, _03491_);
  and _47548_ (_03494_, _03492_, _35815_);
  or _47549_ (_37592_, _03494_, _03493_);
  not _47550_ (_03495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  nor _47551_ (_03496_, _03492_, _03495_);
  and _47552_ (_03497_, _03492_, _35822_);
  or _47553_ (_37593_, _03497_, _03496_);
  not _47554_ (_03498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  nor _47555_ (_03499_, _03492_, _03498_);
  and _47556_ (_03500_, _03492_, _35826_);
  or _47557_ (_37594_, _03500_, _03499_);
  not _47558_ (_03501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  nor _47559_ (_03502_, _03492_, _03501_);
  and _47560_ (_03503_, _03492_, _35830_);
  or _47561_ (_37595_, _03503_, _03502_);
  not _47562_ (_03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  nor _47563_ (_03505_, _03492_, _03504_);
  and _47564_ (_03506_, _03492_, _35834_);
  or _47565_ (_37596_, _03506_, _03505_);
  not _47566_ (_03507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  nor _47567_ (_03508_, _03492_, _03507_);
  and _47568_ (_03509_, _03492_, _35838_);
  or _47569_ (_37597_, _03509_, _03508_);
  not _47570_ (_03510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  nor _47571_ (_03511_, _03492_, _03510_);
  and _47572_ (_03512_, _03492_, _35842_);
  or _47573_ (_37598_, _03512_, _03511_);
  not _47574_ (_03513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  nor _47575_ (_03514_, _03492_, _03513_);
  and _47576_ (_03515_, _03492_, _35846_);
  or _47577_ (_37599_, _03515_, _03514_);
  and _47578_ (_03516_, _00304_, _33632_);
  and _47579_ (_03517_, _03516_, _35572_);
  and _47580_ (_03518_, _03517_, _35815_);
  not _47581_ (_03519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  nor _47582_ (_03520_, _03517_, _03519_);
  or _47583_ (_37600_, _03520_, _03518_);
  and _47584_ (_03521_, _03517_, _35822_);
  not _47585_ (_03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  nor _47586_ (_03523_, _03517_, _03522_);
  or _47587_ (_37601_, _03523_, _03521_);
  and _47588_ (_03524_, _03517_, _35826_);
  not _47589_ (_03525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  nor _47590_ (_03526_, _03517_, _03525_);
  or _47591_ (_37602_, _03526_, _03524_);
  and _47592_ (_03527_, _03517_, _35830_);
  not _47593_ (_03528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  nor _47594_ (_03529_, _03517_, _03528_);
  or _47595_ (_37603_, _03529_, _03527_);
  and _47596_ (_03530_, _03517_, _35834_);
  not _47597_ (_03531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  nor _47598_ (_03532_, _03517_, _03531_);
  or _47599_ (_37604_, _03532_, _03530_);
  and _47600_ (_03533_, _03517_, _35838_);
  not _47601_ (_03534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  nor _47602_ (_03535_, _03517_, _03534_);
  or _47603_ (_37605_, _03535_, _03533_);
  and _47604_ (_03536_, _03517_, _35842_);
  not _47605_ (_03537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  nor _47606_ (_03538_, _03517_, _03537_);
  or _47607_ (_37606_, _03538_, _03536_);
  and _47608_ (_03539_, _03517_, _35846_);
  not _47609_ (_03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  nor _47610_ (_03541_, _03517_, _03540_);
  or _47611_ (_37607_, _03541_, _03539_);
  and _47612_ (_03542_, _03516_, _35817_);
  and _47613_ (_03543_, _03542_, _35815_);
  not _47614_ (_03544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  nor _47615_ (_03545_, _03542_, _03544_);
  or _47616_ (_37608_, _03545_, _03543_);
  and _47617_ (_03546_, _03542_, _35822_);
  not _47618_ (_03547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  nor _47619_ (_03548_, _03542_, _03547_);
  or _47620_ (_37609_, _03548_, _03546_);
  and _47621_ (_03549_, _03542_, _35826_);
  not _47622_ (_03550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  nor _47623_ (_03551_, _03542_, _03550_);
  or _47624_ (_37610_, _03551_, _03549_);
  and _47625_ (_03552_, _03542_, _35830_);
  not _47626_ (_03553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  nor _47627_ (_03554_, _03542_, _03553_);
  or _47628_ (_37611_, _03554_, _03552_);
  and _47629_ (_03555_, _03542_, _35834_);
  not _47630_ (_03556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  nor _47631_ (_03557_, _03542_, _03556_);
  or _47632_ (_37612_, _03557_, _03555_);
  and _47633_ (_03558_, _03542_, _35838_);
  not _47634_ (_03559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  nor _47635_ (_03560_, _03542_, _03559_);
  or _47636_ (_37613_, _03560_, _03558_);
  and _47637_ (_03561_, _03542_, _35842_);
  not _47638_ (_03562_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  nor _47639_ (_03563_, _03542_, _03562_);
  or _47640_ (_37614_, _03563_, _03561_);
  and _47641_ (_03564_, _03542_, _35846_);
  not _47642_ (_03565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  nor _47643_ (_03566_, _03542_, _03565_);
  or _47644_ (_37615_, _03566_, _03564_);
  and _47645_ (_03567_, _03516_, _35851_);
  and _47646_ (_03568_, _03567_, _35815_);
  not _47647_ (_03569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  nor _47648_ (_03570_, _03567_, _03569_);
  or _47649_ (_37616_, _03570_, _03568_);
  and _47650_ (_03571_, _03567_, _35822_);
  not _47651_ (_03572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  nor _47652_ (_03573_, _03567_, _03572_);
  or _47653_ (_37617_, _03573_, _03571_);
  and _47654_ (_03574_, _03567_, _35826_);
  not _47655_ (_03575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  nor _47656_ (_03576_, _03567_, _03575_);
  or _47657_ (_37618_, _03576_, _03574_);
  and _47658_ (_03577_, _03567_, _35830_);
  not _47659_ (_03578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  nor _47660_ (_03579_, _03567_, _03578_);
  or _47661_ (_37619_, _03579_, _03577_);
  and _47662_ (_03580_, _03567_, _35834_);
  not _47663_ (_03581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  nor _47664_ (_03582_, _03567_, _03581_);
  or _47665_ (_37620_, _03582_, _03580_);
  and _47666_ (_03583_, _03567_, _35838_);
  not _47667_ (_03584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  nor _47668_ (_03585_, _03567_, _03584_);
  or _47669_ (_37621_, _03585_, _03583_);
  and _47670_ (_03586_, _03567_, _35842_);
  not _47671_ (_03587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  nor _47672_ (_03588_, _03567_, _03587_);
  or _47673_ (_37622_, _03588_, _03586_);
  and _47674_ (_03589_, _03567_, _35846_);
  not _47675_ (_03590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  nor _47676_ (_03591_, _03567_, _03590_);
  or _47677_ (_37623_, _03591_, _03589_);
  and _47678_ (_03592_, _03516_, _35878_);
  and _47679_ (_03593_, _03592_, _35815_);
  not _47680_ (_03594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  nor _47681_ (_03595_, _03592_, _03594_);
  or _47682_ (_37624_, _03595_, _03593_);
  and _47683_ (_03596_, _03592_, _35822_);
  not _47684_ (_03597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  nor _47685_ (_03598_, _03592_, _03597_);
  or _47686_ (_37625_, _03598_, _03596_);
  and _47687_ (_03599_, _03592_, _35826_);
  not _47688_ (_03600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  nor _47689_ (_03601_, _03592_, _03600_);
  or _47690_ (_37626_, _03601_, _03599_);
  and _47691_ (_03602_, _03592_, _35830_);
  not _47692_ (_03603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  nor _47693_ (_03604_, _03592_, _03603_);
  or _47694_ (_37627_, _03604_, _03602_);
  and _47695_ (_03605_, _03592_, _35834_);
  not _47696_ (_03606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  nor _47697_ (_03607_, _03592_, _03606_);
  or _47698_ (_37628_, _03607_, _03605_);
  and _47699_ (_03608_, _03592_, _35838_);
  not _47700_ (_03609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  nor _47701_ (_03610_, _03592_, _03609_);
  or _47702_ (_37629_, _03610_, _03608_);
  and _47703_ (_03611_, _03592_, _35842_);
  not _47704_ (_03612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  nor _47705_ (_03613_, _03592_, _03612_);
  or _47706_ (_37630_, _03613_, _03611_);
  and _47707_ (_03614_, _03592_, _35846_);
  not _47708_ (_03615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  nor _47709_ (_03616_, _03592_, _03615_);
  or _47710_ (_37631_, _03616_, _03614_);
  and _47711_ (_03617_, _03516_, _35905_);
  and _47712_ (_03618_, _03617_, _35815_);
  not _47713_ (_03619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  nor _47714_ (_03620_, _03617_, _03619_);
  or _47715_ (_37640_, _03620_, _03618_);
  and _47716_ (_03621_, _03617_, _35822_);
  not _47717_ (_03622_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  nor _47718_ (_03623_, _03617_, _03622_);
  or _47719_ (_37641_, _03623_, _03621_);
  and _47720_ (_03624_, _03617_, _35826_);
  not _47721_ (_03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  nor _47722_ (_03626_, _03617_, _03625_);
  or _47723_ (_37642_, _03626_, _03624_);
  and _47724_ (_03627_, _03617_, _35830_);
  not _47725_ (_03628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  nor _47726_ (_03629_, _03617_, _03628_);
  or _47727_ (_37643_, _03629_, _03627_);
  and _47728_ (_03630_, _03617_, _35834_);
  not _47729_ (_03631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  nor _47730_ (_03632_, _03617_, _03631_);
  or _47731_ (_37644_, _03632_, _03630_);
  and _47732_ (_03633_, _03617_, _35838_);
  not _47733_ (_03634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  nor _47734_ (_03635_, _03617_, _03634_);
  or _47735_ (_37645_, _03635_, _03633_);
  and _47736_ (_03636_, _03617_, _35842_);
  not _47737_ (_03637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  nor _47738_ (_03638_, _03617_, _03637_);
  or _47739_ (_37646_, _03638_, _03636_);
  and _47740_ (_03639_, _03617_, _35846_);
  not _47741_ (_03640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  nor _47742_ (_03641_, _03617_, _03640_);
  or _47743_ (_37647_, _03641_, _03639_);
  and _47744_ (_03642_, _03516_, _35931_);
  and _47745_ (_03643_, _03642_, _35815_);
  not _47746_ (_03644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  nor _47747_ (_03645_, _03642_, _03644_);
  or _47748_ (_37648_, _03645_, _03643_);
  and _47749_ (_03646_, _03642_, _35822_);
  not _47750_ (_03647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  nor _47751_ (_03648_, _03642_, _03647_);
  or _47752_ (_37649_, _03648_, _03646_);
  and _47753_ (_03649_, _03642_, _35826_);
  not _47754_ (_03650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  nor _47755_ (_03651_, _03642_, _03650_);
  or _47756_ (_37650_, _03651_, _03649_);
  and _47757_ (_03652_, _03642_, _35830_);
  not _47758_ (_03653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  nor _47759_ (_03654_, _03642_, _03653_);
  or _47760_ (_37651_, _03654_, _03652_);
  and _47761_ (_03655_, _03642_, _35834_);
  not _47762_ (_03656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  nor _47763_ (_03657_, _03642_, _03656_);
  or _47764_ (_37652_, _03657_, _03655_);
  and _47765_ (_03658_, _03642_, _35838_);
  not _47766_ (_03659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  nor _47767_ (_03660_, _03642_, _03659_);
  or _47768_ (_37653_, _03660_, _03658_);
  and _47769_ (_03661_, _03642_, _35842_);
  not _47770_ (_03662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  nor _47771_ (_03663_, _03642_, _03662_);
  or _47772_ (_37654_, _03663_, _03661_);
  and _47773_ (_03664_, _03642_, _35846_);
  not _47774_ (_03665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  nor _47775_ (_03666_, _03642_, _03665_);
  or _47776_ (_37655_, _03666_, _03664_);
  and _47777_ (_03667_, _03516_, _35957_);
  and _47778_ (_03668_, _03667_, _35815_);
  not _47779_ (_03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  nor _47780_ (_03670_, _03667_, _03669_);
  or _47781_ (_37656_, _03670_, _03668_);
  and _47782_ (_03671_, _03667_, _35822_);
  not _47783_ (_03672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  nor _47784_ (_03673_, _03667_, _03672_);
  or _47785_ (_37657_, _03673_, _03671_);
  and _47786_ (_03674_, _03667_, _35826_);
  not _47787_ (_03675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  nor _47788_ (_03676_, _03667_, _03675_);
  or _47789_ (_37658_, _03676_, _03674_);
  and _47790_ (_03677_, _03667_, _35830_);
  not _47791_ (_03678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  nor _47792_ (_03679_, _03667_, _03678_);
  or _47793_ (_37659_, _03679_, _03677_);
  and _47794_ (_03680_, _03667_, _35834_);
  not _47795_ (_03681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  nor _47796_ (_03682_, _03667_, _03681_);
  or _47797_ (_37660_, _03682_, _03680_);
  and _47798_ (_03683_, _03667_, _35838_);
  not _47799_ (_03684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  nor _47800_ (_03685_, _03667_, _03684_);
  or _47801_ (_37661_, _03685_, _03683_);
  and _47802_ (_03686_, _03667_, _35842_);
  not _47803_ (_03687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  nor _47804_ (_03688_, _03667_, _03687_);
  or _47805_ (_37662_, _03688_, _03686_);
  and _47806_ (_03689_, _03667_, _35846_);
  not _47807_ (_03690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  nor _47808_ (_03691_, _03667_, _03690_);
  or _47809_ (_37663_, _03691_, _03689_);
  and _47810_ (_03692_, _03516_, _35983_);
  and _47811_ (_03693_, _03692_, _35815_);
  not _47812_ (_03694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  nor _47813_ (_03695_, _03692_, _03694_);
  or _47814_ (_37664_, _03695_, _03693_);
  and _47815_ (_03696_, _03692_, _35822_);
  not _47816_ (_03697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  nor _47817_ (_03698_, _03692_, _03697_);
  or _47818_ (_37665_, _03698_, _03696_);
  and _47819_ (_03699_, _03692_, _35826_);
  not _47820_ (_03700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  nor _47821_ (_03701_, _03692_, _03700_);
  or _47822_ (_37666_, _03701_, _03699_);
  and _47823_ (_03702_, _03692_, _35830_);
  not _47824_ (_03703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  nor _47825_ (_03704_, _03692_, _03703_);
  or _47826_ (_37667_, _03704_, _03702_);
  and _47827_ (_03705_, _03692_, _35834_);
  not _47828_ (_03706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  nor _47829_ (_03707_, _03692_, _03706_);
  or _47830_ (_37668_, _03707_, _03705_);
  and _47831_ (_03708_, _03692_, _35838_);
  not _47832_ (_03709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  nor _47833_ (_03710_, _03692_, _03709_);
  or _47834_ (_37669_, _03710_, _03708_);
  and _47835_ (_03711_, _03692_, _35842_);
  not _47836_ (_03712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  nor _47837_ (_03713_, _03692_, _03712_);
  or _47838_ (_37670_, _03713_, _03711_);
  and _47839_ (_03714_, _03692_, _35846_);
  not _47840_ (_03715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  nor _47841_ (_03716_, _03692_, _03715_);
  or _47842_ (_37671_, _03716_, _03714_);
  and _47843_ (_03717_, _03516_, _36010_);
  and _47844_ (_03718_, _03717_, _35815_);
  not _47845_ (_03719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  nor _47846_ (_03720_, _03717_, _03719_);
  or _47847_ (_37672_, _03720_, _03718_);
  and _47848_ (_03721_, _03717_, _35822_);
  not _47849_ (_03722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  nor _47850_ (_03723_, _03717_, _03722_);
  or _47851_ (_37673_, _03723_, _03721_);
  and _47852_ (_03724_, _03717_, _35826_);
  not _47853_ (_03725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  nor _47854_ (_03726_, _03717_, _03725_);
  or _47855_ (_37674_, _03726_, _03724_);
  and _47856_ (_03727_, _03717_, _35830_);
  not _47857_ (_03728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  nor _47858_ (_03729_, _03717_, _03728_);
  or _47859_ (_37675_, _03729_, _03727_);
  and _47860_ (_03730_, _03717_, _35834_);
  not _47861_ (_03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  nor _47862_ (_03732_, _03717_, _03731_);
  or _47863_ (_37676_, _03732_, _03730_);
  and _47864_ (_03733_, _03717_, _35838_);
  not _47865_ (_03734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  nor _47866_ (_03735_, _03717_, _03734_);
  or _47867_ (_37677_, _03735_, _03733_);
  and _47868_ (_03736_, _03717_, _35842_);
  not _47869_ (_03737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  nor _47870_ (_03738_, _03717_, _03737_);
  or _47871_ (_37678_, _03738_, _03736_);
  and _47872_ (_03739_, _03717_, _35846_);
  not _47873_ (_03740_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  nor _47874_ (_03741_, _03717_, _03740_);
  or _47875_ (_37679_, _03741_, _03739_);
  and _47876_ (_03742_, _03516_, _36036_);
  and _47877_ (_03743_, _03742_, _35815_);
  not _47878_ (_03744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  nor _47879_ (_03745_, _03742_, _03744_);
  or _47880_ (_37680_, _03745_, _03743_);
  and _47881_ (_03746_, _03742_, _35822_);
  not _47882_ (_03747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  nor _47883_ (_03748_, _03742_, _03747_);
  or _47884_ (_37681_, _03748_, _03746_);
  and _47885_ (_03749_, _03742_, _35826_);
  not _47886_ (_03750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  nor _47887_ (_03751_, _03742_, _03750_);
  or _47888_ (_37682_, _03751_, _03749_);
  and _47889_ (_03752_, _03742_, _35830_);
  not _47890_ (_03753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  nor _47891_ (_03754_, _03742_, _03753_);
  or _47892_ (_37683_, _03754_, _03752_);
  and _47893_ (_03755_, _03742_, _35834_);
  not _47894_ (_03756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  nor _47895_ (_03757_, _03742_, _03756_);
  or _47896_ (_37684_, _03757_, _03755_);
  and _47897_ (_03758_, _03742_, _35838_);
  not _47898_ (_03759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  nor _47899_ (_03760_, _03742_, _03759_);
  or _47900_ (_37685_, _03760_, _03758_);
  and _47901_ (_03761_, _03742_, _35842_);
  not _47902_ (_03762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  nor _47903_ (_03763_, _03742_, _03762_);
  or _47904_ (_37686_, _03763_, _03761_);
  and _47905_ (_03764_, _03742_, _35846_);
  not _47906_ (_03765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  nor _47907_ (_03766_, _03742_, _03765_);
  or _47908_ (_37687_, _03766_, _03764_);
  and _47909_ (_03767_, _03516_, _36062_);
  and _47910_ (_03768_, _03767_, _35815_);
  not _47911_ (_03769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  nor _47912_ (_03770_, _03767_, _03769_);
  or _47913_ (_37688_, _03770_, _03768_);
  and _47914_ (_03771_, _03767_, _35822_);
  not _47915_ (_03772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  nor _47916_ (_03773_, _03767_, _03772_);
  or _47917_ (_37689_, _03773_, _03771_);
  and _47918_ (_03774_, _03767_, _35826_);
  not _47919_ (_03775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  nor _47920_ (_03776_, _03767_, _03775_);
  or _47921_ (_37690_, _03776_, _03774_);
  and _47922_ (_03777_, _03767_, _35830_);
  not _47923_ (_03778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  nor _47924_ (_03779_, _03767_, _03778_);
  or _47925_ (_37691_, _03779_, _03777_);
  and _47926_ (_03780_, _03767_, _35834_);
  not _47927_ (_03781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  nor _47928_ (_03782_, _03767_, _03781_);
  or _47929_ (_37692_, _03782_, _03780_);
  and _47930_ (_03783_, _03767_, _35838_);
  not _47931_ (_03784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  nor _47932_ (_03785_, _03767_, _03784_);
  or _47933_ (_37693_, _03785_, _03783_);
  and _47934_ (_03786_, _03767_, _35842_);
  not _47935_ (_03787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  nor _47936_ (_03788_, _03767_, _03787_);
  or _47937_ (_37694_, _03788_, _03786_);
  and _47938_ (_03789_, _03767_, _35846_);
  not _47939_ (_03790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  nor _47940_ (_03791_, _03767_, _03790_);
  or _47941_ (_37695_, _03791_, _03789_);
  and _47942_ (_03792_, _03516_, _36088_);
  and _47943_ (_03793_, _03792_, _35815_);
  not _47944_ (_03794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  nor _47945_ (_03795_, _03792_, _03794_);
  or _47946_ (_37696_, _03795_, _03793_);
  and _47947_ (_03796_, _03792_, _35822_);
  not _47948_ (_03797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  nor _47949_ (_03798_, _03792_, _03797_);
  or _47950_ (_37697_, _03798_, _03796_);
  and _47951_ (_03799_, _03792_, _35826_);
  not _47952_ (_03800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  nor _47953_ (_03801_, _03792_, _03800_);
  or _47954_ (_37698_, _03801_, _03799_);
  and _47955_ (_03802_, _03792_, _35830_);
  not _47956_ (_03803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  nor _47957_ (_03804_, _03792_, _03803_);
  or _47958_ (_37699_, _03804_, _03802_);
  and _47959_ (_03805_, _03792_, _35834_);
  not _47960_ (_03806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  nor _47961_ (_03807_, _03792_, _03806_);
  or _47962_ (_37700_, _03807_, _03805_);
  and _47963_ (_03808_, _03792_, _35838_);
  not _47964_ (_03809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  nor _47965_ (_03810_, _03792_, _03809_);
  or _47966_ (_37701_, _03810_, _03808_);
  and _47967_ (_03811_, _03792_, _35842_);
  not _47968_ (_03812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  nor _47969_ (_03813_, _03792_, _03812_);
  or _47970_ (_37702_, _03813_, _03811_);
  and _47971_ (_03814_, _03792_, _35846_);
  not _47972_ (_03815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  nor _47973_ (_03816_, _03792_, _03815_);
  or _47974_ (_37703_, _03816_, _03814_);
  and _47975_ (_03817_, _03516_, _36115_);
  and _47976_ (_03818_, _03817_, _35815_);
  not _47977_ (_03819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  nor _47978_ (_03820_, _03817_, _03819_);
  or _47979_ (_37704_, _03820_, _03818_);
  and _47980_ (_03821_, _03817_, _35822_);
  not _47981_ (_03822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  nor _47982_ (_03823_, _03817_, _03822_);
  or _47983_ (_37705_, _03823_, _03821_);
  and _47984_ (_03824_, _03817_, _35826_);
  not _47985_ (_03825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  nor _47986_ (_03826_, _03817_, _03825_);
  or _47987_ (_37706_, _03826_, _03824_);
  and _47988_ (_03827_, _03817_, _35830_);
  not _47989_ (_03828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  nor _47990_ (_03829_, _03817_, _03828_);
  or _47991_ (_37707_, _03829_, _03827_);
  and _47992_ (_03830_, _03817_, _35834_);
  not _47993_ (_03831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  nor _47994_ (_03832_, _03817_, _03831_);
  or _47995_ (_37708_, _03832_, _03830_);
  and _47996_ (_03833_, _03817_, _35838_);
  not _47997_ (_03834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  nor _47998_ (_03835_, _03817_, _03834_);
  or _47999_ (_37709_, _03835_, _03833_);
  and _48000_ (_03836_, _03817_, _35842_);
  not _48001_ (_03837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  nor _48002_ (_03838_, _03817_, _03837_);
  or _48003_ (_37710_, _03838_, _03836_);
  and _48004_ (_03839_, _03817_, _35846_);
  not _48005_ (_03840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  nor _48006_ (_03841_, _03817_, _03840_);
  or _48007_ (_37711_, _03841_, _03839_);
  and _48008_ (_03842_, _03516_, _36141_);
  and _48009_ (_03843_, _03842_, _35815_);
  not _48010_ (_03844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  nor _48011_ (_03845_, _03842_, _03844_);
  or _48012_ (_37712_, _03845_, _03843_);
  and _48013_ (_03846_, _03842_, _35822_);
  not _48014_ (_03847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  nor _48015_ (_03848_, _03842_, _03847_);
  or _48016_ (_37713_, _03848_, _03846_);
  and _48017_ (_03849_, _03842_, _35826_);
  not _48018_ (_03850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  nor _48019_ (_03851_, _03842_, _03850_);
  or _48020_ (_37714_, _03851_, _03849_);
  and _48021_ (_03852_, _03842_, _35830_);
  not _48022_ (_03853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  nor _48023_ (_03854_, _03842_, _03853_);
  or _48024_ (_37715_, _03854_, _03852_);
  and _48025_ (_03855_, _03842_, _35834_);
  not _48026_ (_03856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  nor _48027_ (_03857_, _03842_, _03856_);
  or _48028_ (_37716_, _03857_, _03855_);
  and _48029_ (_03858_, _03842_, _35838_);
  not _48030_ (_03859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  nor _48031_ (_03860_, _03842_, _03859_);
  or _48032_ (_37717_, _03860_, _03858_);
  and _48033_ (_03861_, _03842_, _35842_);
  not _48034_ (_03862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  nor _48035_ (_03863_, _03842_, _03862_);
  or _48036_ (_37718_, _03863_, _03861_);
  and _48037_ (_03864_, _03842_, _35846_);
  not _48038_ (_03865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  nor _48039_ (_03866_, _03842_, _03865_);
  or _48040_ (_37719_, _03866_, _03864_);
  and _48041_ (_03867_, _03516_, _36167_);
  and _48042_ (_03868_, _03867_, _35815_);
  not _48043_ (_03869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  nor _48044_ (_03870_, _03867_, _03869_);
  or _48045_ (_37728_, _03870_, _03868_);
  and _48046_ (_03871_, _03867_, _35822_);
  not _48047_ (_03872_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  nor _48048_ (_03873_, _03867_, _03872_);
  or _48049_ (_37729_, _03873_, _03871_);
  and _48050_ (_03874_, _03867_, _35826_);
  not _48051_ (_03875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  nor _48052_ (_03876_, _03867_, _03875_);
  or _48053_ (_37730_, _03876_, _03874_);
  and _48054_ (_03877_, _03867_, _35830_);
  not _48055_ (_03878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  nor _48056_ (_03879_, _03867_, _03878_);
  or _48057_ (_37731_, _03879_, _03877_);
  and _48058_ (_03880_, _03867_, _35834_);
  not _48059_ (_03881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  nor _48060_ (_03882_, _03867_, _03881_);
  or _48061_ (_37732_, _03882_, _03880_);
  and _48062_ (_03883_, _03867_, _35838_);
  not _48063_ (_03884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  nor _48064_ (_03885_, _03867_, _03884_);
  or _48065_ (_37733_, _03885_, _03883_);
  and _48066_ (_03886_, _03867_, _35842_);
  not _48067_ (_03887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  nor _48068_ (_03888_, _03867_, _03887_);
  or _48069_ (_37734_, _03888_, _03886_);
  and _48070_ (_03889_, _03867_, _35846_);
  not _48071_ (_03890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  nor _48072_ (_03891_, _03867_, _03890_);
  or _48073_ (_37735_, _03891_, _03889_);
  and _48074_ (_03892_, _03516_, _36193_);
  and _48075_ (_03893_, _03892_, _35815_);
  not _48076_ (_03894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  nor _48077_ (_03895_, _03892_, _03894_);
  or _48078_ (_37736_, _03895_, _03893_);
  and _48079_ (_03896_, _03892_, _35822_);
  not _48080_ (_03897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  nor _48081_ (_03898_, _03892_, _03897_);
  or _48082_ (_37737_, _03898_, _03896_);
  and _48083_ (_03899_, _03892_, _35826_);
  not _48084_ (_03900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  nor _48085_ (_03901_, _03892_, _03900_);
  or _48086_ (_37738_, _03901_, _03899_);
  and _48087_ (_03902_, _03892_, _35830_);
  not _48088_ (_03903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  nor _48089_ (_03904_, _03892_, _03903_);
  or _48090_ (_37739_, _03904_, _03902_);
  and _48091_ (_03905_, _03892_, _35834_);
  not _48092_ (_03906_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  nor _48093_ (_03907_, _03892_, _03906_);
  or _48094_ (_37740_, _03907_, _03905_);
  and _48095_ (_03908_, _03892_, _35838_);
  not _48096_ (_03909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  nor _48097_ (_03910_, _03892_, _03909_);
  or _48098_ (_37741_, _03910_, _03908_);
  and _48099_ (_03911_, _03892_, _35842_);
  not _48100_ (_03912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  nor _48101_ (_03913_, _03892_, _03912_);
  or _48102_ (_37742_, _03913_, _03911_);
  and _48103_ (_03914_, _03892_, _35846_);
  not _48104_ (_03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  nor _48105_ (_03916_, _03892_, _03915_);
  or _48106_ (_37743_, _03916_, _03914_);
  and _48107_ (_03917_, _34784_, _34231_);
  and _48108_ (_03918_, _03917_, _35575_);
  and _48109_ (_03919_, _03918_, _35572_);
  and _48110_ (_03920_, _03919_, _35815_);
  not _48111_ (_03921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  nor _48112_ (_03922_, _03919_, _03921_);
  or _48113_ (_37744_, _03922_, _03920_);
  and _48114_ (_03923_, _03919_, _35822_);
  not _48115_ (_03924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  nor _48116_ (_03925_, _03919_, _03924_);
  or _48117_ (_37745_, _03925_, _03923_);
  and _48118_ (_03926_, _03919_, _35826_);
  not _48119_ (_03927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  nor _48120_ (_03928_, _03919_, _03927_);
  or _48121_ (_37746_, _03928_, _03926_);
  and _48122_ (_03929_, _03919_, _35830_);
  not _48123_ (_03930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  nor _48124_ (_03931_, _03919_, _03930_);
  or _48125_ (_37747_, _03931_, _03929_);
  and _48126_ (_03932_, _03919_, _35834_);
  not _48127_ (_03933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  nor _48128_ (_03934_, _03919_, _03933_);
  or _48129_ (_37748_, _03934_, _03932_);
  and _48130_ (_03935_, _03919_, _35838_);
  not _48131_ (_03936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  nor _48132_ (_03937_, _03919_, _03936_);
  or _48133_ (_37749_, _03937_, _03935_);
  and _48134_ (_03938_, _03919_, _35842_);
  not _48135_ (_03939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  nor _48136_ (_03940_, _03919_, _03939_);
  or _48137_ (_37750_, _03940_, _03938_);
  and _48138_ (_03941_, _03919_, _35846_);
  not _48139_ (_03942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  nor _48140_ (_03943_, _03919_, _03942_);
  or _48141_ (_37751_, _03943_, _03941_);
  and _48142_ (_03944_, _03918_, _35817_);
  and _48143_ (_03945_, _03944_, _35815_);
  not _48144_ (_03946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  nor _48145_ (_03947_, _03944_, _03946_);
  or _48146_ (_37752_, _03947_, _03945_);
  and _48147_ (_03948_, _03944_, _35822_);
  not _48148_ (_03949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  nor _48149_ (_03950_, _03944_, _03949_);
  or _48150_ (_37753_, _03950_, _03948_);
  and _48151_ (_03951_, _03944_, _35826_);
  not _48152_ (_03952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  nor _48153_ (_03953_, _03944_, _03952_);
  or _48154_ (_37754_, _03953_, _03951_);
  and _48155_ (_03954_, _03944_, _35830_);
  not _48156_ (_03955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  nor _48157_ (_03956_, _03944_, _03955_);
  or _48158_ (_37755_, _03956_, _03954_);
  and _48159_ (_03957_, _03944_, _35834_);
  not _48160_ (_03958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  nor _48161_ (_03959_, _03944_, _03958_);
  or _48162_ (_37756_, _03959_, _03957_);
  and _48163_ (_03960_, _03944_, _35838_);
  not _48164_ (_03961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  nor _48165_ (_03962_, _03944_, _03961_);
  or _48166_ (_37757_, _03962_, _03960_);
  and _48167_ (_03963_, _03944_, _35842_);
  not _48168_ (_03964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  nor _48169_ (_03965_, _03944_, _03964_);
  or _48170_ (_37758_, _03965_, _03963_);
  and _48171_ (_03966_, _03944_, _35846_);
  not _48172_ (_03967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  nor _48173_ (_03968_, _03944_, _03967_);
  or _48174_ (_37759_, _03968_, _03966_);
  and _48175_ (_03969_, _03918_, _35851_);
  and _48176_ (_03970_, _03969_, _35815_);
  not _48177_ (_03971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  nor _48178_ (_03972_, _03969_, _03971_);
  or _48179_ (_37760_, _03972_, _03970_);
  and _48180_ (_03973_, _03969_, _35822_);
  not _48181_ (_03974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  nor _48182_ (_03975_, _03969_, _03974_);
  or _48183_ (_37761_, _03975_, _03973_);
  and _48184_ (_03976_, _03969_, _35826_);
  not _48185_ (_03977_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  nor _48186_ (_03978_, _03969_, _03977_);
  or _48187_ (_37762_, _03978_, _03976_);
  and _48188_ (_03979_, _03969_, _35830_);
  not _48189_ (_03980_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  nor _48190_ (_03981_, _03969_, _03980_);
  or _48191_ (_37763_, _03981_, _03979_);
  and _48192_ (_03982_, _03969_, _35834_);
  not _48193_ (_03983_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  nor _48194_ (_03984_, _03969_, _03983_);
  or _48195_ (_37764_, _03984_, _03982_);
  and _48196_ (_03985_, _03969_, _35838_);
  not _48197_ (_03986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  nor _48198_ (_03987_, _03969_, _03986_);
  or _48199_ (_37765_, _03987_, _03985_);
  and _48200_ (_03988_, _03969_, _35842_);
  not _48201_ (_03989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  nor _48202_ (_03990_, _03969_, _03989_);
  or _48203_ (_37766_, _03990_, _03988_);
  and _48204_ (_03991_, _03969_, _35846_);
  not _48205_ (_03992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  nor _48206_ (_03993_, _03969_, _03992_);
  or _48207_ (_37767_, _03993_, _03991_);
  and _48208_ (_03994_, _03918_, _35878_);
  and _48209_ (_03995_, _03994_, _35815_);
  not _48210_ (_03996_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  nor _48211_ (_03997_, _03994_, _03996_);
  or _48212_ (_37768_, _03997_, _03995_);
  and _48213_ (_03998_, _03994_, _35822_);
  not _48214_ (_03999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  nor _48215_ (_04000_, _03994_, _03999_);
  or _48216_ (_37769_, _04000_, _03998_);
  and _48217_ (_04001_, _03994_, _35826_);
  not _48218_ (_04002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  nor _48219_ (_04003_, _03994_, _04002_);
  or _48220_ (_37770_, _04003_, _04001_);
  and _48221_ (_04004_, _03994_, _35830_);
  not _48222_ (_04005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  nor _48223_ (_04006_, _03994_, _04005_);
  or _48224_ (_37771_, _04006_, _04004_);
  and _48225_ (_04007_, _03994_, _35834_);
  not _48226_ (_04008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  nor _48227_ (_04009_, _03994_, _04008_);
  or _48228_ (_37772_, _04009_, _04007_);
  and _48229_ (_04010_, _03994_, _35838_);
  not _48230_ (_04011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  nor _48231_ (_04012_, _03994_, _04011_);
  or _48232_ (_37773_, _04012_, _04010_);
  and _48233_ (_04013_, _03994_, _35842_);
  not _48234_ (_04014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  nor _48235_ (_04015_, _03994_, _04014_);
  or _48236_ (_37774_, _04015_, _04013_);
  and _48237_ (_04016_, _03994_, _35846_);
  not _48238_ (_04017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  nor _48239_ (_04018_, _03994_, _04017_);
  or _48240_ (_37775_, _04018_, _04016_);
  and _48241_ (_04019_, _03918_, _35905_);
  and _48242_ (_04020_, _04019_, _35815_);
  not _48243_ (_04021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  nor _48244_ (_04022_, _04019_, _04021_);
  or _48245_ (_37776_, _04022_, _04020_);
  and _48246_ (_04023_, _04019_, _35822_);
  not _48247_ (_04024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  nor _48248_ (_04025_, _04019_, _04024_);
  or _48249_ (_37777_, _04025_, _04023_);
  and _48250_ (_04026_, _04019_, _35826_);
  not _48251_ (_04027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  nor _48252_ (_04028_, _04019_, _04027_);
  or _48253_ (_37778_, _04028_, _04026_);
  and _48254_ (_04029_, _04019_, _35830_);
  not _48255_ (_04030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  nor _48256_ (_04031_, _04019_, _04030_);
  or _48257_ (_37779_, _04031_, _04029_);
  and _48258_ (_04032_, _04019_, _35834_);
  not _48259_ (_04033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  nor _48260_ (_04034_, _04019_, _04033_);
  or _48261_ (_37780_, _04034_, _04032_);
  and _48262_ (_04035_, _04019_, _35838_);
  not _48263_ (_04036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  nor _48264_ (_04037_, _04019_, _04036_);
  or _48265_ (_37781_, _04037_, _04035_);
  and _48266_ (_04038_, _04019_, _35842_);
  not _48267_ (_04039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  nor _48268_ (_04040_, _04019_, _04039_);
  or _48269_ (_37782_, _04040_, _04038_);
  and _48270_ (_04041_, _04019_, _35846_);
  not _48271_ (_04042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  nor _48272_ (_04043_, _04019_, _04042_);
  or _48273_ (_37783_, _04043_, _04041_);
  and _48274_ (_04044_, _03918_, _35931_);
  and _48275_ (_04045_, _04044_, _35815_);
  not _48276_ (_04046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  nor _48277_ (_04047_, _04044_, _04046_);
  or _48278_ (_37784_, _04047_, _04045_);
  and _48279_ (_04048_, _04044_, _35822_);
  not _48280_ (_04049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  nor _48281_ (_04050_, _04044_, _04049_);
  or _48282_ (_37785_, _04050_, _04048_);
  and _48283_ (_04051_, _04044_, _35826_);
  not _48284_ (_04052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  nor _48285_ (_04053_, _04044_, _04052_);
  or _48286_ (_37786_, _04053_, _04051_);
  and _48287_ (_04054_, _04044_, _35830_);
  not _48288_ (_04055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  nor _48289_ (_04056_, _04044_, _04055_);
  or _48290_ (_37787_, _04056_, _04054_);
  and _48291_ (_04057_, _04044_, _35834_);
  not _48292_ (_04058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  nor _48293_ (_04059_, _04044_, _04058_);
  or _48294_ (_37788_, _04059_, _04057_);
  and _48295_ (_04060_, _04044_, _35838_);
  not _48296_ (_04061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  nor _48297_ (_04062_, _04044_, _04061_);
  or _48298_ (_37789_, _04062_, _04060_);
  and _48299_ (_04063_, _04044_, _35842_);
  not _48300_ (_04064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  nor _48301_ (_04065_, _04044_, _04064_);
  or _48302_ (_37790_, _04065_, _04063_);
  and _48303_ (_04066_, _04044_, _35846_);
  not _48304_ (_04067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  nor _48305_ (_04068_, _04044_, _04067_);
  or _48306_ (_37791_, _04068_, _04066_);
  and _48307_ (_04069_, _03918_, _35957_);
  and _48308_ (_04070_, _04069_, _35815_);
  not _48309_ (_04071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  nor _48310_ (_04072_, _04069_, _04071_);
  or _48311_ (_37792_, _04072_, _04070_);
  and _48312_ (_04073_, _04069_, _35822_);
  not _48313_ (_04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  nor _48314_ (_04075_, _04069_, _04074_);
  or _48315_ (_37793_, _04075_, _04073_);
  and _48316_ (_04076_, _04069_, _35826_);
  not _48317_ (_04077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  nor _48318_ (_04078_, _04069_, _04077_);
  or _48319_ (_37794_, _04078_, _04076_);
  and _48320_ (_04079_, _04069_, _35830_);
  not _48321_ (_04080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  nor _48322_ (_04081_, _04069_, _04080_);
  or _48323_ (_37795_, _04081_, _04079_);
  and _48324_ (_04082_, _04069_, _35834_);
  not _48325_ (_04083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  nor _48326_ (_04084_, _04069_, _04083_);
  or _48327_ (_37796_, _04084_, _04082_);
  and _48328_ (_04085_, _04069_, _35838_);
  not _48329_ (_04086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  nor _48330_ (_04087_, _04069_, _04086_);
  or _48331_ (_37797_, _04087_, _04085_);
  and _48332_ (_04088_, _04069_, _35842_);
  not _48333_ (_04089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  nor _48334_ (_04090_, _04069_, _04089_);
  or _48335_ (_37798_, _04090_, _04088_);
  and _48336_ (_04091_, _04069_, _35846_);
  not _48337_ (_04092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  nor _48338_ (_04093_, _04069_, _04092_);
  or _48339_ (_37799_, _04093_, _04091_);
  and _48340_ (_04094_, _03918_, _35983_);
  and _48341_ (_04095_, _04094_, _35815_);
  not _48342_ (_04096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  nor _48343_ (_04097_, _04094_, _04096_);
  or _48344_ (_37800_, _04097_, _04095_);
  and _48345_ (_04098_, _04094_, _35822_);
  not _48346_ (_04099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  nor _48347_ (_04100_, _04094_, _04099_);
  or _48348_ (_37801_, _04100_, _04098_);
  and _48349_ (_04101_, _04094_, _35826_);
  not _48350_ (_04102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  nor _48351_ (_04103_, _04094_, _04102_);
  or _48352_ (_37802_, _04103_, _04101_);
  and _48353_ (_04104_, _04094_, _35830_);
  not _48354_ (_04105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  nor _48355_ (_04106_, _04094_, _04105_);
  or _48356_ (_37803_, _04106_, _04104_);
  and _48357_ (_04107_, _04094_, _35834_);
  not _48358_ (_04108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  nor _48359_ (_04109_, _04094_, _04108_);
  or _48360_ (_37804_, _04109_, _04107_);
  and _48361_ (_04110_, _04094_, _35838_);
  not _48362_ (_04111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  nor _48363_ (_04112_, _04094_, _04111_);
  or _48364_ (_37805_, _04112_, _04110_);
  and _48365_ (_04113_, _04094_, _35842_);
  not _48366_ (_04114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  nor _48367_ (_04115_, _04094_, _04114_);
  or _48368_ (_37806_, _04115_, _04113_);
  and _48369_ (_04116_, _04094_, _35846_);
  not _48370_ (_04117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  nor _48371_ (_04118_, _04094_, _04117_);
  or _48372_ (_37807_, _04118_, _04116_);
  and _48373_ (_04119_, _03918_, _36010_);
  and _48374_ (_04120_, _04119_, _35815_);
  not _48375_ (_04121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  nor _48376_ (_04122_, _04119_, _04121_);
  or _48377_ (_37824_, _04122_, _04120_);
  and _48378_ (_04123_, _04119_, _35822_);
  not _48379_ (_04124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  nor _48380_ (_04125_, _04119_, _04124_);
  or _48381_ (_37825_, _04125_, _04123_);
  and _48382_ (_04126_, _04119_, _35826_);
  not _48383_ (_04127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  nor _48384_ (_04128_, _04119_, _04127_);
  or _48385_ (_37826_, _04128_, _04126_);
  and _48386_ (_04129_, _04119_, _35830_);
  not _48387_ (_04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  nor _48388_ (_04131_, _04119_, _04130_);
  or _48389_ (_37827_, _04131_, _04129_);
  and _48390_ (_04132_, _04119_, _35834_);
  not _48391_ (_04133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  nor _48392_ (_04134_, _04119_, _04133_);
  or _48393_ (_37828_, _04134_, _04132_);
  and _48394_ (_04135_, _04119_, _35838_);
  not _48395_ (_04136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  nor _48396_ (_04137_, _04119_, _04136_);
  or _48397_ (_37829_, _04137_, _04135_);
  and _48398_ (_04138_, _04119_, _35842_);
  not _48399_ (_04139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  nor _48400_ (_04140_, _04119_, _04139_);
  or _48401_ (_37830_, _04140_, _04138_);
  and _48402_ (_04141_, _04119_, _35846_);
  not _48403_ (_04142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  nor _48404_ (_04143_, _04119_, _04142_);
  or _48405_ (_37831_, _04143_, _04141_);
  and _48406_ (_04144_, _03918_, _36036_);
  and _48407_ (_04145_, _04144_, _35815_);
  not _48408_ (_04146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  nor _48409_ (_04147_, _04144_, _04146_);
  or _48410_ (_37832_, _04147_, _04145_);
  and _48411_ (_04148_, _04144_, _35822_);
  not _48412_ (_04149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  nor _48413_ (_04150_, _04144_, _04149_);
  or _48414_ (_37833_, _04150_, _04148_);
  and _48415_ (_04151_, _04144_, _35826_);
  not _48416_ (_04152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  nor _48417_ (_04153_, _04144_, _04152_);
  or _48418_ (_37834_, _04153_, _04151_);
  and _48419_ (_04154_, _04144_, _35830_);
  not _48420_ (_04155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  nor _48421_ (_04156_, _04144_, _04155_);
  or _48422_ (_37835_, _04156_, _04154_);
  and _48423_ (_04157_, _04144_, _35834_);
  not _48424_ (_04158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  nor _48425_ (_04159_, _04144_, _04158_);
  or _48426_ (_37836_, _04159_, _04157_);
  and _48427_ (_04160_, _04144_, _35838_);
  not _48428_ (_04161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  nor _48429_ (_04162_, _04144_, _04161_);
  or _48430_ (_37837_, _04162_, _04160_);
  and _48431_ (_04163_, _04144_, _35842_);
  not _48432_ (_04164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  nor _48433_ (_04165_, _04144_, _04164_);
  or _48434_ (_37838_, _04165_, _04163_);
  and _48435_ (_04166_, _04144_, _35846_);
  not _48436_ (_04167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  nor _48437_ (_04168_, _04144_, _04167_);
  or _48438_ (_37839_, _04168_, _04166_);
  and _48439_ (_04169_, _03918_, _36062_);
  and _48440_ (_04170_, _04169_, _35815_);
  not _48441_ (_04171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  nor _48442_ (_04172_, _04169_, _04171_);
  or _48443_ (_37840_, _04172_, _04170_);
  and _48444_ (_04173_, _04169_, _35822_);
  not _48445_ (_04174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  nor _48446_ (_04175_, _04169_, _04174_);
  or _48447_ (_37841_, _04175_, _04173_);
  and _48448_ (_04176_, _04169_, _35826_);
  not _48449_ (_04177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  nor _48450_ (_04178_, _04169_, _04177_);
  or _48451_ (_37842_, _04178_, _04176_);
  and _48452_ (_04179_, _04169_, _35830_);
  not _48453_ (_04180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  nor _48454_ (_04181_, _04169_, _04180_);
  or _48455_ (_37843_, _04181_, _04179_);
  and _48456_ (_04182_, _04169_, _35834_);
  not _48457_ (_04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  nor _48458_ (_04184_, _04169_, _04183_);
  or _48459_ (_37844_, _04184_, _04182_);
  and _48460_ (_04185_, _04169_, _35838_);
  not _48461_ (_04186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  nor _48462_ (_04187_, _04169_, _04186_);
  or _48463_ (_37845_, _04187_, _04185_);
  and _48464_ (_04188_, _04169_, _35842_);
  not _48465_ (_04189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  nor _48466_ (_04190_, _04169_, _04189_);
  or _48467_ (_37846_, _04190_, _04188_);
  and _48468_ (_04191_, _04169_, _35846_);
  not _48469_ (_04192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  nor _48470_ (_04193_, _04169_, _04192_);
  or _48471_ (_37847_, _04193_, _04191_);
  and _48472_ (_04194_, _03918_, _36088_);
  and _48473_ (_04195_, _04194_, _35815_);
  not _48474_ (_04196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  nor _48475_ (_04197_, _04194_, _04196_);
  or _48476_ (_37848_, _04197_, _04195_);
  and _48477_ (_04198_, _04194_, _35822_);
  not _48478_ (_04199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  nor _48479_ (_04200_, _04194_, _04199_);
  or _48480_ (_37849_, _04200_, _04198_);
  and _48481_ (_04201_, _04194_, _35826_);
  not _48482_ (_04202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  nor _48483_ (_04203_, _04194_, _04202_);
  or _48484_ (_37850_, _04203_, _04201_);
  and _48485_ (_04204_, _04194_, _35830_);
  not _48486_ (_04205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  nor _48487_ (_04206_, _04194_, _04205_);
  or _48488_ (_37851_, _04206_, _04204_);
  and _48489_ (_04207_, _04194_, _35834_);
  not _48490_ (_04208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  nor _48491_ (_04209_, _04194_, _04208_);
  or _48492_ (_37852_, _04209_, _04207_);
  and _48493_ (_04210_, _04194_, _35838_);
  not _48494_ (_04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  nor _48495_ (_04212_, _04194_, _04211_);
  or _48496_ (_37853_, _04212_, _04210_);
  and _48497_ (_04213_, _04194_, _35842_);
  not _48498_ (_04214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  nor _48499_ (_04215_, _04194_, _04214_);
  or _48500_ (_37854_, _04215_, _04213_);
  and _48501_ (_04216_, _04194_, _35846_);
  not _48502_ (_04217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  nor _48503_ (_04218_, _04194_, _04217_);
  or _48504_ (_37855_, _04218_, _04216_);
  and _48505_ (_04219_, _03918_, _36115_);
  and _48506_ (_04220_, _04219_, _35815_);
  not _48507_ (_04221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  nor _48508_ (_04222_, _04219_, _04221_);
  or _48509_ (_37856_, _04222_, _04220_);
  and _48510_ (_04223_, _04219_, _35822_);
  not _48511_ (_04224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  nor _48512_ (_04225_, _04219_, _04224_);
  or _48513_ (_37857_, _04225_, _04223_);
  and _48514_ (_04226_, _04219_, _35826_);
  not _48515_ (_04227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  nor _48516_ (_04228_, _04219_, _04227_);
  or _48517_ (_37858_, _04228_, _04226_);
  and _48518_ (_04229_, _04219_, _35830_);
  not _48519_ (_04230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  nor _48520_ (_04231_, _04219_, _04230_);
  or _48521_ (_37859_, _04231_, _04229_);
  and _48522_ (_04232_, _04219_, _35834_);
  not _48523_ (_04233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  nor _48524_ (_04234_, _04219_, _04233_);
  or _48525_ (_37860_, _04234_, _04232_);
  and _48526_ (_04235_, _04219_, _35838_);
  not _48527_ (_04236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  nor _48528_ (_04237_, _04219_, _04236_);
  or _48529_ (_37861_, _04237_, _04235_);
  and _48530_ (_04238_, _04219_, _35842_);
  not _48531_ (_04239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  nor _48532_ (_04240_, _04219_, _04239_);
  or _48533_ (_37862_, _04240_, _04238_);
  and _48534_ (_04241_, _04219_, _35846_);
  not _48535_ (_04242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  nor _48536_ (_04243_, _04219_, _04242_);
  or _48537_ (_37863_, _04243_, _04241_);
  and _48538_ (_04244_, _03918_, _36141_);
  and _48539_ (_04245_, _04244_, _35815_);
  not _48540_ (_04246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  nor _48541_ (_04247_, _04244_, _04246_);
  or _48542_ (_37864_, _04247_, _04245_);
  and _48543_ (_04248_, _04244_, _35822_);
  not _48544_ (_04249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  nor _48545_ (_04250_, _04244_, _04249_);
  or _48546_ (_37865_, _04250_, _04248_);
  and _48547_ (_04251_, _04244_, _35826_);
  not _48548_ (_04252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  nor _48549_ (_04253_, _04244_, _04252_);
  or _48550_ (_37866_, _04253_, _04251_);
  and _48551_ (_04254_, _04244_, _35830_);
  not _48552_ (_04255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  nor _48553_ (_04256_, _04244_, _04255_);
  or _48554_ (_37867_, _04256_, _04254_);
  and _48555_ (_04257_, _04244_, _35834_);
  not _48556_ (_04258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  nor _48557_ (_04259_, _04244_, _04258_);
  or _48558_ (_37868_, _04259_, _04257_);
  and _48559_ (_04260_, _04244_, _35838_);
  not _48560_ (_04261_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  nor _48561_ (_04262_, _04244_, _04261_);
  or _48562_ (_37869_, _04262_, _04260_);
  and _48563_ (_04263_, _04244_, _35842_);
  not _48564_ (_04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  nor _48565_ (_04265_, _04244_, _04264_);
  or _48566_ (_37870_, _04265_, _04263_);
  and _48567_ (_04266_, _04244_, _35846_);
  not _48568_ (_04267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  nor _48569_ (_04268_, _04244_, _04267_);
  or _48570_ (_37871_, _04268_, _04266_);
  and _48571_ (_04269_, _03918_, _36167_);
  and _48572_ (_04270_, _04269_, _35815_);
  not _48573_ (_04271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  nor _48574_ (_04272_, _04269_, _04271_);
  or _48575_ (_37872_, _04272_, _04270_);
  and _48576_ (_04273_, _04269_, _35822_);
  not _48577_ (_04274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  nor _48578_ (_04275_, _04269_, _04274_);
  or _48579_ (_37873_, _04275_, _04273_);
  and _48580_ (_04276_, _04269_, _35826_);
  not _48581_ (_04277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  nor _48582_ (_04278_, _04269_, _04277_);
  or _48583_ (_37874_, _04278_, _04276_);
  and _48584_ (_04279_, _04269_, _35830_);
  not _48585_ (_04280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  nor _48586_ (_04281_, _04269_, _04280_);
  or _48587_ (_37875_, _04281_, _04279_);
  and _48588_ (_04282_, _04269_, _35834_);
  not _48589_ (_04283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  nor _48590_ (_04284_, _04269_, _04283_);
  or _48591_ (_37876_, _04284_, _04282_);
  and _48592_ (_04285_, _04269_, _35838_);
  not _48593_ (_04286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  nor _48594_ (_04287_, _04269_, _04286_);
  or _48595_ (_37877_, _04287_, _04285_);
  and _48596_ (_04288_, _04269_, _35842_);
  not _48597_ (_04289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  nor _48598_ (_04290_, _04269_, _04289_);
  or _48599_ (_37878_, _04290_, _04288_);
  and _48600_ (_04291_, _04269_, _35846_);
  not _48601_ (_04292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  nor _48602_ (_04293_, _04269_, _04292_);
  or _48603_ (_37879_, _04293_, _04291_);
  and _48604_ (_04294_, _03918_, _36193_);
  and _48605_ (_04295_, _04294_, _35815_);
  not _48606_ (_04296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  nor _48607_ (_04297_, _04294_, _04296_);
  or _48608_ (_37880_, _04297_, _04295_);
  and _48609_ (_04298_, _04294_, _35822_);
  not _48610_ (_04299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  nor _48611_ (_04300_, _04294_, _04299_);
  or _48612_ (_37881_, _04300_, _04298_);
  and _48613_ (_04301_, _04294_, _35826_);
  not _48614_ (_04302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  nor _48615_ (_04303_, _04294_, _04302_);
  or _48616_ (_37882_, _04303_, _04301_);
  and _48617_ (_04304_, _04294_, _35830_);
  not _48618_ (_04305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  nor _48619_ (_04306_, _04294_, _04305_);
  or _48620_ (_37883_, _04306_, _04304_);
  and _48621_ (_04307_, _04294_, _35834_);
  not _48622_ (_04308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  nor _48623_ (_04309_, _04294_, _04308_);
  or _48624_ (_37884_, _04309_, _04307_);
  and _48625_ (_04310_, _04294_, _35838_);
  not _48626_ (_04311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  nor _48627_ (_04312_, _04294_, _04311_);
  or _48628_ (_37885_, _04312_, _04310_);
  and _48629_ (_04313_, _04294_, _35842_);
  not _48630_ (_04314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  nor _48631_ (_04315_, _04294_, _04314_);
  or _48632_ (_37886_, _04315_, _04313_);
  and _48633_ (_04316_, _04294_, _35846_);
  not _48634_ (_04317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  nor _48635_ (_04318_, _04294_, _04317_);
  or _48636_ (_37887_, _04318_, _04316_);
  not _48637_ (_04319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and _48638_ (_04320_, _36220_, _34231_);
  and _48639_ (_04321_, _04320_, _35572_);
  nor _48640_ (_04322_, _04321_, _04319_);
  and _48641_ (_04323_, _04321_, _35815_);
  or _48642_ (_37888_, _04323_, _04322_);
  not _48643_ (_04324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  nor _48644_ (_04325_, _04321_, _04324_);
  and _48645_ (_04326_, _04321_, _35822_);
  or _48646_ (_37889_, _04326_, _04325_);
  not _48647_ (_04327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  nor _48648_ (_04328_, _04321_, _04327_);
  and _48649_ (_04329_, _04321_, _35826_);
  or _48650_ (_37890_, _04329_, _04328_);
  not _48651_ (_04330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  nor _48652_ (_04331_, _04321_, _04330_);
  and _48653_ (_04332_, _04321_, _35830_);
  or _48654_ (_37891_, _04332_, _04331_);
  not _48655_ (_04333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  nor _48656_ (_04334_, _04321_, _04333_);
  and _48657_ (_04335_, _04321_, _35834_);
  or _48658_ (_37892_, _04335_, _04334_);
  not _48659_ (_04336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  nor _48660_ (_04337_, _04321_, _04336_);
  and _48661_ (_04338_, _04321_, _35838_);
  or _48662_ (_37893_, _04338_, _04337_);
  not _48663_ (_04339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  nor _48664_ (_04340_, _04321_, _04339_);
  and _48665_ (_04341_, _04321_, _35842_);
  or _48666_ (_37894_, _04341_, _04340_);
  not _48667_ (_04342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  nor _48668_ (_04343_, _04321_, _04342_);
  and _48669_ (_04344_, _04321_, _35846_);
  or _48670_ (_37895_, _04344_, _04343_);
  not _48671_ (_04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  and _48672_ (_04346_, _04320_, _35817_);
  nor _48673_ (_04347_, _04346_, _04345_);
  and _48674_ (_04348_, _04346_, _35815_);
  or _48675_ (_37896_, _04348_, _04347_);
  not _48676_ (_04349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  nor _48677_ (_04350_, _04346_, _04349_);
  and _48678_ (_04351_, _04346_, _35822_);
  or _48679_ (_37897_, _04351_, _04350_);
  not _48680_ (_04352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  nor _48681_ (_04353_, _04346_, _04352_);
  and _48682_ (_04354_, _04346_, _35826_);
  or _48683_ (_37898_, _04354_, _04353_);
  not _48684_ (_04355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  nor _48685_ (_04356_, _04346_, _04355_);
  and _48686_ (_04357_, _04346_, _35830_);
  or _48687_ (_37899_, _04357_, _04356_);
  not _48688_ (_04358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  nor _48689_ (_04359_, _04346_, _04358_);
  and _48690_ (_04360_, _04346_, _35834_);
  or _48691_ (_37900_, _04360_, _04359_);
  not _48692_ (_04361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  nor _48693_ (_04362_, _04346_, _04361_);
  and _48694_ (_04363_, _04346_, _35838_);
  or _48695_ (_37901_, _04363_, _04362_);
  not _48696_ (_04364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  nor _48697_ (_04365_, _04346_, _04364_);
  and _48698_ (_04366_, _04346_, _35842_);
  or _48699_ (_37902_, _04366_, _04365_);
  not _48700_ (_04367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  nor _48701_ (_04368_, _04346_, _04367_);
  and _48702_ (_04369_, _04346_, _35846_);
  or _48703_ (_37903_, _04369_, _04368_);
  not _48704_ (_04370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  and _48705_ (_04371_, _04320_, _35851_);
  nor _48706_ (_04372_, _04371_, _04370_);
  and _48707_ (_04373_, _04371_, _35815_);
  or _48708_ (_37912_, _04373_, _04372_);
  not _48709_ (_04374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  nor _48710_ (_04375_, _04371_, _04374_);
  and _48711_ (_04376_, _04371_, _35822_);
  or _48712_ (_37913_, _04376_, _04375_);
  not _48713_ (_04377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  nor _48714_ (_04378_, _04371_, _04377_);
  and _48715_ (_04379_, _04371_, _35826_);
  or _48716_ (_37914_, _04379_, _04378_);
  not _48717_ (_04380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  nor _48718_ (_04381_, _04371_, _04380_);
  and _48719_ (_04382_, _04371_, _35830_);
  or _48720_ (_37915_, _04382_, _04381_);
  not _48721_ (_04383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  nor _48722_ (_04384_, _04371_, _04383_);
  and _48723_ (_04385_, _04371_, _35834_);
  or _48724_ (_37916_, _04385_, _04384_);
  not _48725_ (_04386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  nor _48726_ (_04387_, _04371_, _04386_);
  and _48727_ (_04388_, _04371_, _35838_);
  or _48728_ (_37917_, _04388_, _04387_);
  not _48729_ (_04389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  nor _48730_ (_04390_, _04371_, _04389_);
  and _48731_ (_04391_, _04371_, _35842_);
  or _48732_ (_37918_, _04391_, _04390_);
  not _48733_ (_04392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  nor _48734_ (_04393_, _04371_, _04392_);
  and _48735_ (_04394_, _04371_, _35846_);
  or _48736_ (_37919_, _04394_, _04393_);
  not _48737_ (_04395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and _48738_ (_04396_, _04320_, _35878_);
  nor _48739_ (_04397_, _04396_, _04395_);
  and _48740_ (_04398_, _04396_, _35815_);
  or _48741_ (_37920_, _04398_, _04397_);
  not _48742_ (_04399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  nor _48743_ (_04400_, _04396_, _04399_);
  and _48744_ (_04401_, _04396_, _35822_);
  or _48745_ (_37921_, _04401_, _04400_);
  not _48746_ (_04402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  nor _48747_ (_04403_, _04396_, _04402_);
  and _48748_ (_04404_, _04396_, _35826_);
  or _48749_ (_37922_, _04404_, _04403_);
  not _48750_ (_04405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  nor _48751_ (_04406_, _04396_, _04405_);
  and _48752_ (_04407_, _04396_, _35830_);
  or _48753_ (_37923_, _04407_, _04406_);
  not _48754_ (_04408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  nor _48755_ (_04409_, _04396_, _04408_);
  and _48756_ (_04410_, _04396_, _35834_);
  or _48757_ (_37924_, _04410_, _04409_);
  not _48758_ (_04411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  nor _48759_ (_04412_, _04396_, _04411_);
  and _48760_ (_04413_, _04396_, _35838_);
  or _48761_ (_37925_, _04413_, _04412_);
  not _48762_ (_04414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  nor _48763_ (_04415_, _04396_, _04414_);
  and _48764_ (_04416_, _04396_, _35842_);
  or _48765_ (_37926_, _04416_, _04415_);
  not _48766_ (_04417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  nor _48767_ (_04418_, _04396_, _04417_);
  and _48768_ (_04419_, _04396_, _35846_);
  or _48769_ (_37927_, _04419_, _04418_);
  not _48770_ (_04420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and _48771_ (_04421_, _04320_, _35905_);
  nor _48772_ (_04422_, _04421_, _04420_);
  and _48773_ (_04423_, _04421_, _35815_);
  or _48774_ (_37928_, _04423_, _04422_);
  not _48775_ (_04424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  nor _48776_ (_04425_, _04421_, _04424_);
  and _48777_ (_04426_, _04421_, _35822_);
  or _48778_ (_37929_, _04426_, _04425_);
  not _48779_ (_04427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  nor _48780_ (_04428_, _04421_, _04427_);
  and _48781_ (_04429_, _04421_, _35826_);
  or _48782_ (_37930_, _04429_, _04428_);
  not _48783_ (_04430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  nor _48784_ (_04431_, _04421_, _04430_);
  and _48785_ (_04432_, _04421_, _35830_);
  or _48786_ (_37931_, _04432_, _04431_);
  not _48787_ (_04433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  nor _48788_ (_04434_, _04421_, _04433_);
  and _48789_ (_04435_, _04421_, _35834_);
  or _48790_ (_37932_, _04435_, _04434_);
  not _48791_ (_04436_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  nor _48792_ (_04437_, _04421_, _04436_);
  and _48793_ (_04438_, _04421_, _35838_);
  or _48794_ (_37933_, _04438_, _04437_);
  not _48795_ (_04439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  nor _48796_ (_04440_, _04421_, _04439_);
  and _48797_ (_04441_, _04421_, _35842_);
  or _48798_ (_37934_, _04441_, _04440_);
  not _48799_ (_04442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  nor _48800_ (_04443_, _04421_, _04442_);
  and _48801_ (_04444_, _04421_, _35846_);
  or _48802_ (_37935_, _04444_, _04443_);
  not _48803_ (_04445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  and _48804_ (_04446_, _04320_, _35931_);
  nor _48805_ (_04447_, _04446_, _04445_);
  and _48806_ (_04448_, _04446_, _35815_);
  or _48807_ (_37936_, _04448_, _04447_);
  not _48808_ (_04449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  nor _48809_ (_04450_, _04446_, _04449_);
  and _48810_ (_04451_, _04446_, _35822_);
  or _48811_ (_37937_, _04451_, _04450_);
  not _48812_ (_04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  nor _48813_ (_04453_, _04446_, _04452_);
  and _48814_ (_04454_, _04446_, _35826_);
  or _48815_ (_37938_, _04454_, _04453_);
  not _48816_ (_04455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  nor _48817_ (_04456_, _04446_, _04455_);
  and _48818_ (_04457_, _04446_, _35830_);
  or _48819_ (_37939_, _04457_, _04456_);
  not _48820_ (_04458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  nor _48821_ (_04459_, _04446_, _04458_);
  and _48822_ (_04460_, _04446_, _35834_);
  or _48823_ (_37940_, _04460_, _04459_);
  not _48824_ (_04461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  nor _48825_ (_04462_, _04446_, _04461_);
  and _48826_ (_04463_, _04446_, _35838_);
  or _48827_ (_37941_, _04463_, _04462_);
  not _48828_ (_04464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  nor _48829_ (_04465_, _04446_, _04464_);
  and _48830_ (_04466_, _04446_, _35842_);
  or _48831_ (_37942_, _04466_, _04465_);
  not _48832_ (_04467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  nor _48833_ (_04468_, _04446_, _04467_);
  and _48834_ (_04469_, _04446_, _35846_);
  or _48835_ (_37943_, _04469_, _04468_);
  not _48836_ (_04470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  and _48837_ (_04471_, _04320_, _35957_);
  nor _48838_ (_04472_, _04471_, _04470_);
  and _48839_ (_04473_, _04471_, _35815_);
  or _48840_ (_37944_, _04473_, _04472_);
  not _48841_ (_04474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  nor _48842_ (_04475_, _04471_, _04474_);
  and _48843_ (_04476_, _04471_, _35822_);
  or _48844_ (_37945_, _04476_, _04475_);
  not _48845_ (_04477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  nor _48846_ (_04478_, _04471_, _04477_);
  and _48847_ (_04479_, _04471_, _35826_);
  or _48848_ (_37946_, _04479_, _04478_);
  not _48849_ (_04480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  nor _48850_ (_04481_, _04471_, _04480_);
  and _48851_ (_04482_, _04471_, _35830_);
  or _48852_ (_37947_, _04482_, _04481_);
  not _48853_ (_04483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  nor _48854_ (_04484_, _04471_, _04483_);
  and _48855_ (_04485_, _04471_, _35834_);
  or _48856_ (_37948_, _04485_, _04484_);
  not _48857_ (_04486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  nor _48858_ (_04487_, _04471_, _04486_);
  and _48859_ (_04488_, _04471_, _35838_);
  or _48860_ (_37949_, _04488_, _04487_);
  not _48861_ (_04489_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  nor _48862_ (_04490_, _04471_, _04489_);
  and _48863_ (_04491_, _04471_, _35842_);
  or _48864_ (_37950_, _04491_, _04490_);
  not _48865_ (_04492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  nor _48866_ (_04493_, _04471_, _04492_);
  and _48867_ (_04494_, _04471_, _35846_);
  or _48868_ (_37951_, _04494_, _04493_);
  not _48869_ (_04495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and _48870_ (_04496_, _04320_, _35983_);
  nor _48871_ (_04497_, _04496_, _04495_);
  and _48872_ (_04498_, _04496_, _35815_);
  or _48873_ (_37952_, _04498_, _04497_);
  not _48874_ (_04499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  nor _48875_ (_04500_, _04496_, _04499_);
  and _48876_ (_04501_, _04496_, _35822_);
  or _48877_ (_37953_, _04501_, _04500_);
  not _48878_ (_04502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  nor _48879_ (_04503_, _04496_, _04502_);
  and _48880_ (_04504_, _04496_, _35826_);
  or _48881_ (_37954_, _04504_, _04503_);
  not _48882_ (_04505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  nor _48883_ (_04506_, _04496_, _04505_);
  and _48884_ (_04507_, _04496_, _35830_);
  or _48885_ (_37955_, _04507_, _04506_);
  not _48886_ (_04508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  nor _48887_ (_04509_, _04496_, _04508_);
  and _48888_ (_04510_, _04496_, _35834_);
  or _48889_ (_37956_, _04510_, _04509_);
  not _48890_ (_04511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  nor _48891_ (_04512_, _04496_, _04511_);
  and _48892_ (_04513_, _04496_, _35838_);
  or _48893_ (_37957_, _04513_, _04512_);
  not _48894_ (_04514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  nor _48895_ (_04515_, _04496_, _04514_);
  and _48896_ (_04516_, _04496_, _35842_);
  or _48897_ (_37958_, _04516_, _04515_);
  not _48898_ (_04517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  nor _48899_ (_04518_, _04496_, _04517_);
  and _48900_ (_04519_, _04496_, _35846_);
  or _48901_ (_37959_, _04519_, _04518_);
  not _48902_ (_04520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  and _48903_ (_04521_, _04320_, _36010_);
  nor _48904_ (_04522_, _04521_, _04520_);
  and _48905_ (_04523_, _04521_, _35815_);
  or _48906_ (_37960_, _04523_, _04522_);
  not _48907_ (_04524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  nor _48908_ (_04525_, _04521_, _04524_);
  and _48909_ (_04526_, _04521_, _35822_);
  or _48910_ (_37961_, _04526_, _04525_);
  not _48911_ (_04527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  nor _48912_ (_04528_, _04521_, _04527_);
  and _48913_ (_04529_, _04521_, _35826_);
  or _48914_ (_37962_, _04529_, _04528_);
  not _48915_ (_04530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  nor _48916_ (_04531_, _04521_, _04530_);
  and _48917_ (_04532_, _04521_, _35830_);
  or _48918_ (_37963_, _04532_, _04531_);
  not _48919_ (_04533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  nor _48920_ (_04534_, _04521_, _04533_);
  and _48921_ (_04535_, _04521_, _35834_);
  or _48922_ (_37964_, _04535_, _04534_);
  not _48923_ (_04536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  nor _48924_ (_04537_, _04521_, _04536_);
  and _48925_ (_04538_, _04521_, _35838_);
  or _48926_ (_37965_, _04538_, _04537_);
  not _48927_ (_04539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  nor _48928_ (_04540_, _04521_, _04539_);
  and _48929_ (_04541_, _04521_, _35842_);
  or _48930_ (_37966_, _04541_, _04540_);
  not _48931_ (_04542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  nor _48932_ (_04543_, _04521_, _04542_);
  and _48933_ (_04544_, _04521_, _35846_);
  or _48934_ (_37967_, _04544_, _04543_);
  not _48935_ (_04545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and _48936_ (_04546_, _04320_, _36036_);
  nor _48937_ (_04547_, _04546_, _04545_);
  and _48938_ (_04548_, _04546_, _35815_);
  or _48939_ (_37968_, _04548_, _04547_);
  not _48940_ (_04549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  nor _48941_ (_04550_, _04546_, _04549_);
  and _48942_ (_04551_, _04546_, _35822_);
  or _48943_ (_37969_, _04551_, _04550_);
  not _48944_ (_04552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  nor _48945_ (_04553_, _04546_, _04552_);
  and _48946_ (_04554_, _04546_, _35826_);
  or _48947_ (_37970_, _04554_, _04553_);
  not _48948_ (_04555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  nor _48949_ (_04556_, _04546_, _04555_);
  and _48950_ (_04557_, _04546_, _35830_);
  or _48951_ (_37971_, _04557_, _04556_);
  not _48952_ (_04558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  nor _48953_ (_04559_, _04546_, _04558_);
  and _48954_ (_04560_, _04546_, _35834_);
  or _48955_ (_37972_, _04560_, _04559_);
  not _48956_ (_04561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  nor _48957_ (_04562_, _04546_, _04561_);
  and _48958_ (_04563_, _04546_, _35838_);
  or _48959_ (_37973_, _04563_, _04562_);
  not _48960_ (_04564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  nor _48961_ (_04565_, _04546_, _04564_);
  and _48962_ (_04566_, _04546_, _35842_);
  or _48963_ (_37974_, _04566_, _04565_);
  not _48964_ (_04567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  nor _48965_ (_04568_, _04546_, _04567_);
  and _48966_ (_04569_, _04546_, _35846_);
  or _48967_ (_37975_, _04569_, _04568_);
  not _48968_ (_04570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and _48969_ (_04571_, _04320_, _36062_);
  nor _48970_ (_04572_, _04571_, _04570_);
  and _48971_ (_04573_, _04571_, _35815_);
  or _48972_ (_37976_, _04573_, _04572_);
  not _48973_ (_04574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  nor _48974_ (_04575_, _04571_, _04574_);
  and _48975_ (_04576_, _04571_, _35822_);
  or _48976_ (_37977_, _04576_, _04575_);
  not _48977_ (_04577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  nor _48978_ (_04578_, _04571_, _04577_);
  and _48979_ (_04579_, _04571_, _35826_);
  or _48980_ (_37978_, _04579_, _04578_);
  not _48981_ (_04580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  nor _48982_ (_04581_, _04571_, _04580_);
  and _48983_ (_04582_, _04571_, _35830_);
  or _48984_ (_37979_, _04582_, _04581_);
  not _48985_ (_04583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  nor _48986_ (_04584_, _04571_, _04583_);
  and _48987_ (_04585_, _04571_, _35834_);
  or _48988_ (_37980_, _04585_, _04584_);
  not _48989_ (_04586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  nor _48990_ (_04587_, _04571_, _04586_);
  and _48991_ (_04588_, _04571_, _35838_);
  or _48992_ (_37981_, _04588_, _04587_);
  not _48993_ (_04589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  nor _48994_ (_04590_, _04571_, _04589_);
  and _48995_ (_04591_, _04571_, _35842_);
  or _48996_ (_37982_, _04591_, _04590_);
  not _48997_ (_04592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  nor _48998_ (_04593_, _04571_, _04592_);
  and _48999_ (_04594_, _04571_, _35846_);
  or _49000_ (_37983_, _04594_, _04593_);
  not _49001_ (_04595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  and _49002_ (_04596_, _04320_, _36088_);
  nor _49003_ (_04597_, _04596_, _04595_);
  and _49004_ (_04598_, _04596_, _35815_);
  or _49005_ (_37984_, _04598_, _04597_);
  not _49006_ (_04599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  nor _49007_ (_04600_, _04596_, _04599_);
  and _49008_ (_04601_, _04596_, _35822_);
  or _49009_ (_37985_, _04601_, _04600_);
  not _49010_ (_04602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  nor _49011_ (_04603_, _04596_, _04602_);
  and _49012_ (_04604_, _04596_, _35826_);
  or _49013_ (_37986_, _04604_, _04603_);
  not _49014_ (_04605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  nor _49015_ (_04606_, _04596_, _04605_);
  and _49016_ (_04607_, _04596_, _35830_);
  or _49017_ (_37987_, _04607_, _04606_);
  not _49018_ (_04608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  nor _49019_ (_04609_, _04596_, _04608_);
  and _49020_ (_04610_, _04596_, _35834_);
  or _49021_ (_37988_, _04610_, _04609_);
  not _49022_ (_04611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  nor _49023_ (_04612_, _04596_, _04611_);
  and _49024_ (_04613_, _04596_, _35838_);
  or _49025_ (_37989_, _04613_, _04612_);
  not _49026_ (_04614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  nor _49027_ (_04615_, _04596_, _04614_);
  and _49028_ (_04616_, _04596_, _35842_);
  or _49029_ (_37990_, _04616_, _04615_);
  not _49030_ (_04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  nor _49031_ (_04618_, _04596_, _04617_);
  and _49032_ (_04619_, _04596_, _35846_);
  or _49033_ (_37991_, _04619_, _04618_);
  not _49034_ (_04620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  and _49035_ (_04621_, _04320_, _36115_);
  nor _49036_ (_04622_, _04621_, _04620_);
  and _49037_ (_04623_, _04621_, _35815_);
  or _49038_ (_38000_, _04623_, _04622_);
  not _49039_ (_04624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  nor _49040_ (_04625_, _04621_, _04624_);
  and _49041_ (_04626_, _04621_, _35822_);
  or _49042_ (_38001_, _04626_, _04625_);
  not _49043_ (_04627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  nor _49044_ (_04628_, _04621_, _04627_);
  and _49045_ (_04629_, _04621_, _35826_);
  or _49046_ (_38002_, _04629_, _04628_);
  not _49047_ (_04630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  nor _49048_ (_04631_, _04621_, _04630_);
  and _49049_ (_04632_, _04621_, _35830_);
  or _49050_ (_38003_, _04632_, _04631_);
  not _49051_ (_04633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  nor _49052_ (_04634_, _04621_, _04633_);
  and _49053_ (_04635_, _04621_, _35834_);
  or _49054_ (_38004_, _04635_, _04634_);
  not _49055_ (_04636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  nor _49056_ (_04637_, _04621_, _04636_);
  and _49057_ (_04638_, _04621_, _35838_);
  or _49058_ (_38005_, _04638_, _04637_);
  not _49059_ (_04639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  nor _49060_ (_04640_, _04621_, _04639_);
  and _49061_ (_04641_, _04621_, _35842_);
  or _49062_ (_38006_, _04641_, _04640_);
  not _49063_ (_04642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  nor _49064_ (_04643_, _04621_, _04642_);
  and _49065_ (_04644_, _04621_, _35846_);
  or _49066_ (_38007_, _04644_, _04643_);
  not _49067_ (_04645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and _49068_ (_04646_, _04320_, _36141_);
  nor _49069_ (_04647_, _04646_, _04645_);
  and _49070_ (_04648_, _04646_, _35815_);
  or _49071_ (_38008_, _04648_, _04647_);
  not _49072_ (_04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  nor _49073_ (_04650_, _04646_, _04649_);
  and _49074_ (_04651_, _04646_, _35822_);
  or _49075_ (_38009_, _04651_, _04650_);
  not _49076_ (_04652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  nor _49077_ (_04653_, _04646_, _04652_);
  and _49078_ (_04654_, _04646_, _35826_);
  or _49079_ (_38010_, _04654_, _04653_);
  not _49080_ (_04655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  nor _49081_ (_04656_, _04646_, _04655_);
  and _49082_ (_04657_, _04646_, _35830_);
  or _49083_ (_38011_, _04657_, _04656_);
  not _49084_ (_04658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  nor _49085_ (_04659_, _04646_, _04658_);
  and _49086_ (_04660_, _04646_, _35834_);
  or _49087_ (_38012_, _04660_, _04659_);
  not _49088_ (_04661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  nor _49089_ (_04662_, _04646_, _04661_);
  and _49090_ (_04663_, _04646_, _35838_);
  or _49091_ (_38013_, _04663_, _04662_);
  not _49092_ (_04664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  nor _49093_ (_04665_, _04646_, _04664_);
  and _49094_ (_04666_, _04646_, _35842_);
  or _49095_ (_38014_, _04666_, _04665_);
  not _49096_ (_04667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  nor _49097_ (_04668_, _04646_, _04667_);
  and _49098_ (_04669_, _04646_, _35846_);
  or _49099_ (_38015_, _04669_, _04668_);
  not _49100_ (_04670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and _49101_ (_04671_, _04320_, _36167_);
  nor _49102_ (_04672_, _04671_, _04670_);
  and _49103_ (_04673_, _04671_, _35815_);
  or _49104_ (_38016_, _04673_, _04672_);
  not _49105_ (_04674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  nor _49106_ (_04675_, _04671_, _04674_);
  and _49107_ (_04676_, _04671_, _35822_);
  or _49108_ (_38017_, _04676_, _04675_);
  not _49109_ (_04677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  nor _49110_ (_04678_, _04671_, _04677_);
  and _49111_ (_04679_, _04671_, _35826_);
  or _49112_ (_38018_, _04679_, _04678_);
  not _49113_ (_04680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  nor _49114_ (_04681_, _04671_, _04680_);
  and _49115_ (_04682_, _04671_, _35830_);
  or _49116_ (_38019_, _04682_, _04681_);
  not _49117_ (_04683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  nor _49118_ (_04684_, _04671_, _04683_);
  and _49119_ (_04685_, _04671_, _35834_);
  or _49120_ (_38020_, _04685_, _04684_);
  not _49121_ (_04686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  nor _49122_ (_04687_, _04671_, _04686_);
  and _49123_ (_04688_, _04671_, _35838_);
  or _49124_ (_38021_, _04688_, _04687_);
  not _49125_ (_04689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  nor _49126_ (_04690_, _04671_, _04689_);
  and _49127_ (_04691_, _04671_, _35842_);
  or _49128_ (_38022_, _04691_, _04690_);
  not _49129_ (_04692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  nor _49130_ (_04693_, _04671_, _04692_);
  and _49131_ (_04694_, _04671_, _35846_);
  or _49132_ (_38023_, _04694_, _04693_);
  not _49133_ (_04695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  and _49134_ (_04696_, _04320_, _36193_);
  nor _49135_ (_04697_, _04696_, _04695_);
  and _49136_ (_04698_, _04696_, _35815_);
  or _49137_ (_38024_, _04698_, _04697_);
  not _49138_ (_04699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  nor _49139_ (_04700_, _04696_, _04699_);
  and _49140_ (_04701_, _04696_, _35822_);
  or _49141_ (_38025_, _04701_, _04700_);
  not _49142_ (_04702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  nor _49143_ (_04703_, _04696_, _04702_);
  and _49144_ (_04704_, _04696_, _35826_);
  or _49145_ (_38026_, _04704_, _04703_);
  not _49146_ (_04705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  nor _49147_ (_04706_, _04696_, _04705_);
  and _49148_ (_04707_, _04696_, _35830_);
  or _49149_ (_38027_, _04707_, _04706_);
  not _49150_ (_04708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  nor _49151_ (_04709_, _04696_, _04708_);
  and _49152_ (_04710_, _04696_, _35834_);
  or _49153_ (_38028_, _04710_, _04709_);
  not _49154_ (_04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  nor _49155_ (_04712_, _04696_, _04711_);
  and _49156_ (_04713_, _04696_, _35838_);
  or _49157_ (_38029_, _04713_, _04712_);
  not _49158_ (_04714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  nor _49159_ (_04715_, _04696_, _04714_);
  and _49160_ (_04716_, _04696_, _35842_);
  or _49161_ (_38030_, _04716_, _04715_);
  not _49162_ (_04717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  nor _49163_ (_04718_, _04696_, _04717_);
  and _49164_ (_04719_, _04696_, _35846_);
  or _49165_ (_38031_, _04719_, _04718_);
  and _49166_ (_04720_, _36622_, _34231_);
  and _49167_ (_04721_, _04720_, _35572_);
  and _49168_ (_04722_, _04721_, _35815_);
  not _49169_ (_04723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  nor _49170_ (_04724_, _04721_, _04723_);
  or _49171_ (_38032_, _04724_, _04722_);
  and _49172_ (_04725_, _04721_, _35822_);
  not _49173_ (_04726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  nor _49174_ (_04727_, _04721_, _04726_);
  or _49175_ (_38033_, _04727_, _04725_);
  and _49176_ (_04728_, _04721_, _35826_);
  not _49177_ (_04729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  nor _49178_ (_04730_, _04721_, _04729_);
  or _49179_ (_38034_, _04730_, _04728_);
  and _49180_ (_04731_, _04721_, _35830_);
  not _49181_ (_04732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  nor _49182_ (_04733_, _04721_, _04732_);
  or _49183_ (_38035_, _04733_, _04731_);
  and _49184_ (_04734_, _04721_, _35834_);
  not _49185_ (_04735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  nor _49186_ (_04736_, _04721_, _04735_);
  or _49187_ (_38036_, _04736_, _04734_);
  and _49188_ (_04737_, _04721_, _35838_);
  not _49189_ (_04738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  nor _49190_ (_04739_, _04721_, _04738_);
  or _49191_ (_38037_, _04739_, _04737_);
  and _49192_ (_04740_, _04721_, _35842_);
  not _49193_ (_04741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  nor _49194_ (_04742_, _04721_, _04741_);
  or _49195_ (_38038_, _04742_, _04740_);
  and _49196_ (_04743_, _04721_, _35846_);
  not _49197_ (_04744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  nor _49198_ (_04745_, _04721_, _04744_);
  or _49199_ (_38039_, _04745_, _04743_);
  and _49200_ (_04746_, _04720_, _35817_);
  and _49201_ (_04747_, _04746_, _35815_);
  not _49202_ (_04748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  nor _49203_ (_04749_, _04746_, _04748_);
  or _49204_ (_38040_, _04749_, _04747_);
  and _49205_ (_04750_, _04746_, _35822_);
  not _49206_ (_04751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  nor _49207_ (_04752_, _04746_, _04751_);
  or _49208_ (_38041_, _04752_, _04750_);
  and _49209_ (_04753_, _04746_, _35826_);
  not _49210_ (_04754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  nor _49211_ (_04755_, _04746_, _04754_);
  or _49212_ (_38042_, _04755_, _04753_);
  and _49213_ (_04756_, _04746_, _35830_);
  not _49214_ (_04757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  nor _49215_ (_04758_, _04746_, _04757_);
  or _49216_ (_38043_, _04758_, _04756_);
  and _49217_ (_04759_, _04746_, _35834_);
  not _49218_ (_04760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  nor _49219_ (_04761_, _04746_, _04760_);
  or _49220_ (_38044_, _04761_, _04759_);
  and _49221_ (_04762_, _04746_, _35838_);
  not _49222_ (_04763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  nor _49223_ (_04764_, _04746_, _04763_);
  or _49224_ (_38045_, _04764_, _04762_);
  and _49225_ (_04765_, _04746_, _35842_);
  not _49226_ (_04766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  nor _49227_ (_04767_, _04746_, _04766_);
  or _49228_ (_38046_, _04767_, _04765_);
  and _49229_ (_04768_, _04746_, _35846_);
  not _49230_ (_04769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  nor _49231_ (_04770_, _04746_, _04769_);
  or _49232_ (_38047_, _04770_, _04768_);
  and _49233_ (_04771_, _04720_, _35851_);
  and _49234_ (_04772_, _04771_, _35815_);
  not _49235_ (_04773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  nor _49236_ (_04774_, _04771_, _04773_);
  or _49237_ (_38048_, _04774_, _04772_);
  and _49238_ (_04775_, _04771_, _35822_);
  not _49239_ (_04776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  nor _49240_ (_04777_, _04771_, _04776_);
  or _49241_ (_38049_, _04777_, _04775_);
  and _49242_ (_04778_, _04771_, _35826_);
  not _49243_ (_04779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  nor _49244_ (_04780_, _04771_, _04779_);
  or _49245_ (_38050_, _04780_, _04778_);
  and _49246_ (_04781_, _04771_, _35830_);
  not _49247_ (_04782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  nor _49248_ (_04783_, _04771_, _04782_);
  or _49249_ (_38051_, _04783_, _04781_);
  and _49250_ (_04784_, _04771_, _35834_);
  not _49251_ (_04785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  nor _49252_ (_04786_, _04771_, _04785_);
  or _49253_ (_38052_, _04786_, _04784_);
  and _49254_ (_04787_, _04771_, _35838_);
  not _49255_ (_04788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  nor _49256_ (_04789_, _04771_, _04788_);
  or _49257_ (_38053_, _04789_, _04787_);
  and _49258_ (_04790_, _04771_, _35842_);
  not _49259_ (_04791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  nor _49260_ (_04792_, _04771_, _04791_);
  or _49261_ (_38054_, _04792_, _04790_);
  and _49262_ (_04793_, _04771_, _35846_);
  not _49263_ (_04794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  nor _49264_ (_04795_, _04771_, _04794_);
  or _49265_ (_38055_, _04795_, _04793_);
  and _49266_ (_04796_, _04720_, _35878_);
  and _49267_ (_04797_, _04796_, _35815_);
  not _49268_ (_04798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  nor _49269_ (_04799_, _04796_, _04798_);
  or _49270_ (_38056_, _04799_, _04797_);
  and _49271_ (_04800_, _04796_, _35822_);
  not _49272_ (_04801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  nor _49273_ (_04802_, _04796_, _04801_);
  or _49274_ (_38057_, _04802_, _04800_);
  and _49275_ (_04803_, _04796_, _35826_);
  not _49276_ (_04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  nor _49277_ (_04805_, _04796_, _04804_);
  or _49278_ (_38058_, _04805_, _04803_);
  and _49279_ (_04806_, _04796_, _35830_);
  not _49280_ (_04807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  nor _49281_ (_04808_, _04796_, _04807_);
  or _49282_ (_38059_, _04808_, _04806_);
  and _49283_ (_04809_, _04796_, _35834_);
  not _49284_ (_04810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  nor _49285_ (_04811_, _04796_, _04810_);
  or _49286_ (_38060_, _04811_, _04809_);
  and _49287_ (_04812_, _04796_, _35838_);
  not _49288_ (_04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  nor _49289_ (_04814_, _04796_, _04813_);
  or _49290_ (_38061_, _04814_, _04812_);
  and _49291_ (_04815_, _04796_, _35842_);
  not _49292_ (_04816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  nor _49293_ (_04817_, _04796_, _04816_);
  or _49294_ (_38062_, _04817_, _04815_);
  and _49295_ (_04818_, _04796_, _35846_);
  not _49296_ (_04819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  nor _49297_ (_04820_, _04796_, _04819_);
  or _49298_ (_38063_, _04820_, _04818_);
  and _49299_ (_04821_, _04720_, _35905_);
  and _49300_ (_04822_, _04821_, _35815_);
  not _49301_ (_04823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  nor _49302_ (_04824_, _04821_, _04823_);
  or _49303_ (_38064_, _04824_, _04822_);
  and _49304_ (_04825_, _04821_, _35822_);
  not _49305_ (_04826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  nor _49306_ (_04827_, _04821_, _04826_);
  or _49307_ (_38065_, _04827_, _04825_);
  and _49308_ (_04828_, _04821_, _35826_);
  not _49309_ (_04829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  nor _49310_ (_04830_, _04821_, _04829_);
  or _49311_ (_38066_, _04830_, _04828_);
  and _49312_ (_04831_, _04821_, _35830_);
  not _49313_ (_04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  nor _49314_ (_04833_, _04821_, _04832_);
  or _49315_ (_38067_, _04833_, _04831_);
  and _49316_ (_04834_, _04821_, _35834_);
  not _49317_ (_04835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  nor _49318_ (_04836_, _04821_, _04835_);
  or _49319_ (_38068_, _04836_, _04834_);
  and _49320_ (_04837_, _04821_, _35838_);
  not _49321_ (_04838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  nor _49322_ (_04839_, _04821_, _04838_);
  or _49323_ (_38069_, _04839_, _04837_);
  and _49324_ (_04840_, _04821_, _35842_);
  not _49325_ (_04841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  nor _49326_ (_04842_, _04821_, _04841_);
  or _49327_ (_38070_, _04842_, _04840_);
  and _49328_ (_04843_, _04821_, _35846_);
  not _49329_ (_04844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  nor _49330_ (_04845_, _04821_, _04844_);
  or _49331_ (_38071_, _04845_, _04843_);
  and _49332_ (_04846_, _04720_, _35931_);
  and _49333_ (_04847_, _04846_, _35815_);
  not _49334_ (_04848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  nor _49335_ (_04849_, _04846_, _04848_);
  or _49336_ (_38072_, _04849_, _04847_);
  and _49337_ (_04850_, _04846_, _35822_);
  not _49338_ (_04851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  nor _49339_ (_04852_, _04846_, _04851_);
  or _49340_ (_38073_, _04852_, _04850_);
  and _49341_ (_04853_, _04846_, _35826_);
  not _49342_ (_04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  nor _49343_ (_04855_, _04846_, _04854_);
  or _49344_ (_38074_, _04855_, _04853_);
  and _49345_ (_04856_, _04846_, _35830_);
  not _49346_ (_04857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  nor _49347_ (_04858_, _04846_, _04857_);
  or _49348_ (_38075_, _04858_, _04856_);
  and _49349_ (_04859_, _04846_, _35834_);
  not _49350_ (_04860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  nor _49351_ (_04861_, _04846_, _04860_);
  or _49352_ (_38076_, _04861_, _04859_);
  and _49353_ (_04862_, _04846_, _35838_);
  not _49354_ (_04863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  nor _49355_ (_04864_, _04846_, _04863_);
  or _49356_ (_38077_, _04864_, _04862_);
  and _49357_ (_04865_, _04846_, _35842_);
  not _49358_ (_04866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  nor _49359_ (_04867_, _04846_, _04866_);
  or _49360_ (_38078_, _04867_, _04865_);
  and _49361_ (_04868_, _04846_, _35846_);
  not _49362_ (_04869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  nor _49363_ (_04870_, _04846_, _04869_);
  or _49364_ (_38079_, _04870_, _04868_);
  and _49365_ (_04871_, _04720_, _35957_);
  and _49366_ (_04872_, _04871_, _35815_);
  not _49367_ (_04873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  nor _49368_ (_04874_, _04871_, _04873_);
  or _49369_ (_38088_, _04874_, _04872_);
  and _49370_ (_04875_, _04871_, _35822_);
  not _49371_ (_04876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  nor _49372_ (_04877_, _04871_, _04876_);
  or _49373_ (_38089_, _04877_, _04875_);
  and _49374_ (_04878_, _04871_, _35826_);
  not _49375_ (_04879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  nor _49376_ (_04880_, _04871_, _04879_);
  or _49377_ (_38090_, _04880_, _04878_);
  and _49378_ (_04881_, _04871_, _35830_);
  not _49379_ (_04882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  nor _49380_ (_04883_, _04871_, _04882_);
  or _49381_ (_38091_, _04883_, _04881_);
  and _49382_ (_04884_, _04871_, _35834_);
  not _49383_ (_04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  nor _49384_ (_04886_, _04871_, _04885_);
  or _49385_ (_38092_, _04886_, _04884_);
  and _49386_ (_04887_, _04871_, _35838_);
  not _49387_ (_04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  nor _49388_ (_04889_, _04871_, _04888_);
  or _49389_ (_38093_, _04889_, _04887_);
  and _49390_ (_04890_, _04871_, _35842_);
  not _49391_ (_04891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  nor _49392_ (_04892_, _04871_, _04891_);
  or _49393_ (_38094_, _04892_, _04890_);
  and _49394_ (_04893_, _04871_, _35846_);
  not _49395_ (_04894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  nor _49396_ (_04895_, _04871_, _04894_);
  or _49397_ (_38095_, _04895_, _04893_);
  and _49398_ (_04896_, _04720_, _35983_);
  and _49399_ (_04897_, _04896_, _35815_);
  not _49400_ (_04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  nor _49401_ (_04899_, _04896_, _04898_);
  or _49402_ (_38096_, _04899_, _04897_);
  and _49403_ (_04900_, _04896_, _35822_);
  not _49404_ (_04901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  nor _49405_ (_04902_, _04896_, _04901_);
  or _49406_ (_38097_, _04902_, _04900_);
  and _49407_ (_04903_, _04896_, _35826_);
  not _49408_ (_04904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  nor _49409_ (_04905_, _04896_, _04904_);
  or _49410_ (_38098_, _04905_, _04903_);
  and _49411_ (_04906_, _04896_, _35830_);
  not _49412_ (_04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  nor _49413_ (_04908_, _04896_, _04907_);
  or _49414_ (_38099_, _04908_, _04906_);
  and _49415_ (_04909_, _04896_, _35834_);
  not _49416_ (_04910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  nor _49417_ (_04911_, _04896_, _04910_);
  or _49418_ (_38100_, _04911_, _04909_);
  and _49419_ (_04912_, _04896_, _35838_);
  not _49420_ (_04913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  nor _49421_ (_04914_, _04896_, _04913_);
  or _49422_ (_38101_, _04914_, _04912_);
  and _49423_ (_04915_, _04896_, _35842_);
  not _49424_ (_04916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  nor _49425_ (_04917_, _04896_, _04916_);
  or _49426_ (_38102_, _04917_, _04915_);
  and _49427_ (_04918_, _04896_, _35846_);
  not _49428_ (_04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  nor _49429_ (_04920_, _04896_, _04919_);
  or _49430_ (_38103_, _04920_, _04918_);
  and _49431_ (_04921_, _04720_, _36010_);
  and _49432_ (_04922_, _04921_, _35815_);
  not _49433_ (_04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  nor _49434_ (_04924_, _04921_, _04923_);
  or _49435_ (_38104_, _04924_, _04922_);
  and _49436_ (_04925_, _04921_, _35822_);
  not _49437_ (_04926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  nor _49438_ (_04927_, _04921_, _04926_);
  or _49439_ (_38105_, _04927_, _04925_);
  and _49440_ (_04928_, _04921_, _35826_);
  not _49441_ (_04929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  nor _49442_ (_04930_, _04921_, _04929_);
  or _49443_ (_38106_, _04930_, _04928_);
  and _49444_ (_04931_, _04921_, _35830_);
  not _49445_ (_04932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  nor _49446_ (_04933_, _04921_, _04932_);
  or _49447_ (_38107_, _04933_, _04931_);
  and _49448_ (_04934_, _04921_, _35834_);
  not _49449_ (_04935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  nor _49450_ (_04936_, _04921_, _04935_);
  or _49451_ (_38108_, _04936_, _04934_);
  and _49452_ (_04937_, _04921_, _35838_);
  not _49453_ (_04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  nor _49454_ (_04939_, _04921_, _04938_);
  or _49455_ (_38109_, _04939_, _04937_);
  and _49456_ (_04940_, _04921_, _35842_);
  not _49457_ (_04941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  nor _49458_ (_04942_, _04921_, _04941_);
  or _49459_ (_38110_, _04942_, _04940_);
  and _49460_ (_04943_, _04921_, _35846_);
  not _49461_ (_04944_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  nor _49462_ (_04945_, _04921_, _04944_);
  or _49463_ (_38111_, _04945_, _04943_);
  and _49464_ (_04946_, _04720_, _36036_);
  and _49465_ (_04947_, _04946_, _35815_);
  not _49466_ (_04948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  nor _49467_ (_04949_, _04946_, _04948_);
  or _49468_ (_38112_, _04949_, _04947_);
  and _49469_ (_04950_, _04946_, _35822_);
  not _49470_ (_04951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  nor _49471_ (_04952_, _04946_, _04951_);
  or _49472_ (_38113_, _04952_, _04950_);
  and _49473_ (_04953_, _04946_, _35826_);
  not _49474_ (_04954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  nor _49475_ (_04955_, _04946_, _04954_);
  or _49476_ (_38114_, _04955_, _04953_);
  and _49477_ (_04956_, _04946_, _35830_);
  not _49478_ (_04957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  nor _49479_ (_04958_, _04946_, _04957_);
  or _49480_ (_38115_, _04958_, _04956_);
  and _49481_ (_04959_, _04946_, _35834_);
  not _49482_ (_04960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  nor _49483_ (_04961_, _04946_, _04960_);
  or _49484_ (_38116_, _04961_, _04959_);
  and _49485_ (_04962_, _04946_, _35838_);
  not _49486_ (_04963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  nor _49487_ (_04964_, _04946_, _04963_);
  or _49488_ (_38117_, _04964_, _04962_);
  and _49489_ (_04965_, _04946_, _35842_);
  not _49490_ (_04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  nor _49491_ (_04967_, _04946_, _04966_);
  or _49492_ (_38118_, _04967_, _04965_);
  and _49493_ (_04968_, _04946_, _35846_);
  not _49494_ (_04969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  nor _49495_ (_04970_, _04946_, _04969_);
  or _49496_ (_38119_, _04970_, _04968_);
  and _49497_ (_04971_, _04720_, _36062_);
  and _49498_ (_04972_, _04971_, _35815_);
  not _49499_ (_04973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  nor _49500_ (_04974_, _04971_, _04973_);
  or _49501_ (_38120_, _04974_, _04972_);
  and _49502_ (_04975_, _04971_, _35822_);
  not _49503_ (_04976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  nor _49504_ (_04977_, _04971_, _04976_);
  or _49505_ (_38121_, _04977_, _04975_);
  and _49506_ (_04978_, _04971_, _35826_);
  not _49507_ (_04979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  nor _49508_ (_04980_, _04971_, _04979_);
  or _49509_ (_38122_, _04980_, _04978_);
  and _49510_ (_04981_, _04971_, _35830_);
  not _49511_ (_04982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  nor _49512_ (_04983_, _04971_, _04982_);
  or _49513_ (_38123_, _04983_, _04981_);
  and _49514_ (_04984_, _04971_, _35834_);
  not _49515_ (_04985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  nor _49516_ (_04986_, _04971_, _04985_);
  or _49517_ (_38124_, _04986_, _04984_);
  and _49518_ (_04987_, _04971_, _35838_);
  not _49519_ (_04988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  nor _49520_ (_04989_, _04971_, _04988_);
  or _49521_ (_38125_, _04989_, _04987_);
  and _49522_ (_04990_, _04971_, _35842_);
  not _49523_ (_04991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  nor _49524_ (_04992_, _04971_, _04991_);
  or _49525_ (_38126_, _04992_, _04990_);
  and _49526_ (_04993_, _04971_, _35846_);
  not _49527_ (_04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  nor _49528_ (_04995_, _04971_, _04994_);
  or _49529_ (_38127_, _04995_, _04993_);
  and _49530_ (_04996_, _04720_, _36088_);
  and _49531_ (_04997_, _04996_, _35815_);
  not _49532_ (_04998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  nor _49533_ (_04999_, _04996_, _04998_);
  or _49534_ (_38128_, _04999_, _04997_);
  and _49535_ (_05000_, _04996_, _35822_);
  not _49536_ (_05001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  nor _49537_ (_05002_, _04996_, _05001_);
  or _49538_ (_38129_, _05002_, _05000_);
  and _49539_ (_05003_, _04996_, _35826_);
  not _49540_ (_05004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  nor _49541_ (_05005_, _04996_, _05004_);
  or _49542_ (_38130_, _05005_, _05003_);
  and _49543_ (_05006_, _04996_, _35830_);
  not _49544_ (_05007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  nor _49545_ (_05008_, _04996_, _05007_);
  or _49546_ (_38131_, _05008_, _05006_);
  and _49547_ (_05009_, _04996_, _35834_);
  not _49548_ (_05010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  nor _49549_ (_05011_, _04996_, _05010_);
  or _49550_ (_38132_, _05011_, _05009_);
  and _49551_ (_05012_, _04996_, _35838_);
  not _49552_ (_05013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  nor _49553_ (_05014_, _04996_, _05013_);
  or _49554_ (_38133_, _05014_, _05012_);
  and _49555_ (_05015_, _04996_, _35842_);
  not _49556_ (_05016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  nor _49557_ (_05017_, _04996_, _05016_);
  or _49558_ (_38134_, _05017_, _05015_);
  and _49559_ (_05018_, _04996_, _35846_);
  not _49560_ (_05019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  nor _49561_ (_05020_, _04996_, _05019_);
  or _49562_ (_38135_, _05020_, _05018_);
  and _49563_ (_05021_, _04720_, _36115_);
  and _49564_ (_05022_, _05021_, _35815_);
  not _49565_ (_05023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  nor _49566_ (_05024_, _05021_, _05023_);
  or _49567_ (_38136_, _05024_, _05022_);
  and _49568_ (_05025_, _05021_, _35822_);
  not _49569_ (_05026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  nor _49570_ (_05027_, _05021_, _05026_);
  or _49571_ (_38137_, _05027_, _05025_);
  and _49572_ (_05028_, _05021_, _35826_);
  not _49573_ (_05029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  nor _49574_ (_05030_, _05021_, _05029_);
  or _49575_ (_38138_, _05030_, _05028_);
  and _49576_ (_05031_, _05021_, _35830_);
  not _49577_ (_05032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  nor _49578_ (_05033_, _05021_, _05032_);
  or _49579_ (_38139_, _05033_, _05031_);
  and _49580_ (_05034_, _05021_, _35834_);
  not _49581_ (_05035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  nor _49582_ (_05036_, _05021_, _05035_);
  or _49583_ (_38140_, _05036_, _05034_);
  and _49584_ (_05037_, _05021_, _35838_);
  not _49585_ (_05038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  nor _49586_ (_05039_, _05021_, _05038_);
  or _49587_ (_38141_, _05039_, _05037_);
  and _49588_ (_05040_, _05021_, _35842_);
  not _49589_ (_05041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  nor _49590_ (_05042_, _05021_, _05041_);
  or _49591_ (_38142_, _05042_, _05040_);
  and _49592_ (_05043_, _05021_, _35846_);
  not _49593_ (_05044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  nor _49594_ (_05045_, _05021_, _05044_);
  or _49595_ (_38143_, _05045_, _05043_);
  and _49596_ (_05046_, _04720_, _36141_);
  and _49597_ (_05047_, _05046_, _35815_);
  not _49598_ (_05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  nor _49599_ (_05049_, _05046_, _05048_);
  or _49600_ (_38144_, _05049_, _05047_);
  and _49601_ (_05050_, _05046_, _35822_);
  not _49602_ (_05051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  nor _49603_ (_05052_, _05046_, _05051_);
  or _49604_ (_38145_, _05052_, _05050_);
  and _49605_ (_05053_, _05046_, _35826_);
  not _49606_ (_05054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  nor _49607_ (_05055_, _05046_, _05054_);
  or _49608_ (_38146_, _05055_, _05053_);
  and _49609_ (_05056_, _05046_, _35830_);
  not _49610_ (_05057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  nor _49611_ (_05058_, _05046_, _05057_);
  or _49612_ (_38147_, _05058_, _05056_);
  and _49613_ (_05059_, _05046_, _35834_);
  not _49614_ (_05060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  nor _49615_ (_05061_, _05046_, _05060_);
  or _49616_ (_38148_, _05061_, _05059_);
  and _49617_ (_05062_, _05046_, _35838_);
  not _49618_ (_05063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  nor _49619_ (_05064_, _05046_, _05063_);
  or _49620_ (_38149_, _05064_, _05062_);
  and _49621_ (_05065_, _05046_, _35842_);
  not _49622_ (_05066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  nor _49623_ (_05067_, _05046_, _05066_);
  or _49624_ (_38150_, _05067_, _05065_);
  and _49625_ (_05068_, _05046_, _35846_);
  not _49626_ (_05069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  nor _49627_ (_05070_, _05046_, _05069_);
  or _49628_ (_38151_, _05070_, _05068_);
  and _49629_ (_05071_, _04720_, _36167_);
  and _49630_ (_05072_, _05071_, _35815_);
  not _49631_ (_05073_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  nor _49632_ (_05074_, _05071_, _05073_);
  or _49633_ (_38152_, _05074_, _05072_);
  and _49634_ (_05075_, _05071_, _35822_);
  not _49635_ (_05076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  nor _49636_ (_05077_, _05071_, _05076_);
  or _49637_ (_38153_, _05077_, _05075_);
  and _49638_ (_05078_, _05071_, _35826_);
  not _49639_ (_05079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  nor _49640_ (_05080_, _05071_, _05079_);
  or _49641_ (_38154_, _05080_, _05078_);
  and _49642_ (_05081_, _05071_, _35830_);
  not _49643_ (_05082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  nor _49644_ (_05083_, _05071_, _05082_);
  or _49645_ (_38155_, _05083_, _05081_);
  and _49646_ (_05084_, _05071_, _35834_);
  not _49647_ (_05085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  nor _49648_ (_05086_, _05071_, _05085_);
  or _49649_ (_38156_, _05086_, _05084_);
  and _49650_ (_05087_, _05071_, _35838_);
  not _49651_ (_05088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  nor _49652_ (_05089_, _05071_, _05088_);
  or _49653_ (_38157_, _05089_, _05087_);
  and _49654_ (_05090_, _05071_, _35842_);
  not _49655_ (_05091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  nor _49656_ (_05092_, _05071_, _05091_);
  or _49657_ (_38158_, _05092_, _05090_);
  and _49658_ (_05093_, _05071_, _35846_);
  not _49659_ (_05094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  nor _49660_ (_05095_, _05071_, _05094_);
  or _49661_ (_38159_, _05095_, _05093_);
  and _49662_ (_05096_, _04720_, _36193_);
  and _49663_ (_05097_, _05096_, _35815_);
  not _49664_ (_05098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  nor _49665_ (_05099_, _05096_, _05098_);
  or _49666_ (_38160_, _05099_, _05097_);
  and _49667_ (_05100_, _05096_, _35822_);
  not _49668_ (_05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  nor _49669_ (_05102_, _05096_, _05101_);
  or _49670_ (_38161_, _05102_, _05100_);
  and _49671_ (_05103_, _05096_, _35826_);
  not _49672_ (_05104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  nor _49673_ (_05105_, _05096_, _05104_);
  or _49674_ (_38162_, _05105_, _05103_);
  and _49675_ (_05106_, _05096_, _35830_);
  not _49676_ (_05107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  nor _49677_ (_05108_, _05096_, _05107_);
  or _49678_ (_38163_, _05108_, _05106_);
  and _49679_ (_05109_, _05096_, _35834_);
  not _49680_ (_05110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  nor _49681_ (_05111_, _05096_, _05110_);
  or _49682_ (_38164_, _05111_, _05109_);
  and _49683_ (_05112_, _05096_, _35838_);
  not _49684_ (_05113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  nor _49685_ (_05114_, _05096_, _05113_);
  or _49686_ (_38165_, _05114_, _05112_);
  and _49687_ (_05115_, _05096_, _35842_);
  not _49688_ (_05116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  nor _49689_ (_05117_, _05096_, _05116_);
  or _49690_ (_38166_, _05117_, _05115_);
  and _49691_ (_05118_, _05096_, _35846_);
  not _49692_ (_05119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  nor _49693_ (_05120_, _05096_, _05119_);
  or _49694_ (_38167_, _05120_, _05118_);
  and _49695_ (_05121_, _00304_, _34231_);
  and _49696_ (_05122_, _05121_, _35572_);
  and _49697_ (_05123_, _05122_, _35815_);
  not _49698_ (_05124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  nor _49699_ (_05125_, _05122_, _05124_);
  or _49700_ (_38176_, _05125_, _05123_);
  and _49701_ (_05126_, _05122_, _35822_);
  not _49702_ (_05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  nor _49703_ (_05128_, _05122_, _05127_);
  or _49704_ (_38177_, _05128_, _05126_);
  and _49705_ (_05129_, _05122_, _35826_);
  not _49706_ (_05130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  nor _49707_ (_05131_, _05122_, _05130_);
  or _49708_ (_38178_, _05131_, _05129_);
  and _49709_ (_05132_, _05122_, _35830_);
  not _49710_ (_05133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  nor _49711_ (_05134_, _05122_, _05133_);
  or _49712_ (_38179_, _05134_, _05132_);
  and _49713_ (_05135_, _05122_, _35834_);
  not _49714_ (_05136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  nor _49715_ (_05137_, _05122_, _05136_);
  or _49716_ (_38180_, _05137_, _05135_);
  and _49717_ (_05138_, _05122_, _35838_);
  not _49718_ (_05139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  nor _49719_ (_05140_, _05122_, _05139_);
  or _49720_ (_38181_, _05140_, _05138_);
  and _49721_ (_05141_, _05122_, _35842_);
  not _49722_ (_05142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  nor _49723_ (_05143_, _05122_, _05142_);
  or _49724_ (_38182_, _05143_, _05141_);
  and _49725_ (_05144_, _05122_, _35846_);
  not _49726_ (_05145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  nor _49727_ (_05146_, _05122_, _05145_);
  or _49728_ (_38183_, _05146_, _05144_);
  and _49729_ (_05147_, _05121_, _35817_);
  and _49730_ (_05148_, _05147_, _35815_);
  not _49731_ (_05149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  nor _49732_ (_05150_, _05147_, _05149_);
  or _49733_ (_38184_, _05150_, _05148_);
  and _49734_ (_05151_, _05147_, _35822_);
  not _49735_ (_05152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  nor _49736_ (_05153_, _05147_, _05152_);
  or _49737_ (_38185_, _05153_, _05151_);
  and _49738_ (_05154_, _05147_, _35826_);
  not _49739_ (_05155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  nor _49740_ (_05156_, _05147_, _05155_);
  or _49741_ (_38186_, _05156_, _05154_);
  and _49742_ (_05157_, _05147_, _35830_);
  not _49743_ (_05158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  nor _49744_ (_05159_, _05147_, _05158_);
  or _49745_ (_38187_, _05159_, _05157_);
  and _49746_ (_05160_, _05147_, _35834_);
  not _49747_ (_05161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  nor _49748_ (_05162_, _05147_, _05161_);
  or _49749_ (_38188_, _05162_, _05160_);
  and _49750_ (_05163_, _05147_, _35838_);
  not _49751_ (_05164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  nor _49752_ (_05165_, _05147_, _05164_);
  or _49753_ (_38189_, _05165_, _05163_);
  and _49754_ (_05166_, _05147_, _35842_);
  not _49755_ (_05167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  nor _49756_ (_05168_, _05147_, _05167_);
  or _49757_ (_38190_, _05168_, _05166_);
  and _49758_ (_05169_, _05147_, _35846_);
  not _49759_ (_05170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  nor _49760_ (_05171_, _05147_, _05170_);
  or _49761_ (_38191_, _05171_, _05169_);
  and _49762_ (_05172_, _05121_, _35851_);
  and _49763_ (_05173_, _05172_, _35815_);
  not _49764_ (_05174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  nor _49765_ (_05175_, _05172_, _05174_);
  or _49766_ (_38192_, _05175_, _05173_);
  and _49767_ (_05176_, _05172_, _35822_);
  not _49768_ (_05177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  nor _49769_ (_05178_, _05172_, _05177_);
  or _49770_ (_38193_, _05178_, _05176_);
  and _49771_ (_05179_, _05172_, _35826_);
  not _49772_ (_05180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  nor _49773_ (_05181_, _05172_, _05180_);
  or _49774_ (_38194_, _05181_, _05179_);
  and _49775_ (_05182_, _05172_, _35830_);
  not _49776_ (_05183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  nor _49777_ (_05184_, _05172_, _05183_);
  or _49778_ (_38195_, _05184_, _05182_);
  and _49779_ (_05185_, _05172_, _35834_);
  not _49780_ (_05186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  nor _49781_ (_05187_, _05172_, _05186_);
  or _49782_ (_38196_, _05187_, _05185_);
  and _49783_ (_05188_, _05172_, _35838_);
  not _49784_ (_05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  nor _49785_ (_05190_, _05172_, _05189_);
  or _49786_ (_38197_, _05190_, _05188_);
  and _49787_ (_05191_, _05172_, _35842_);
  not _49788_ (_05192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  nor _49789_ (_05193_, _05172_, _05192_);
  or _49790_ (_38198_, _05193_, _05191_);
  and _49791_ (_05194_, _05172_, _35846_);
  not _49792_ (_05195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  nor _49793_ (_05196_, _05172_, _05195_);
  or _49794_ (_38199_, _05196_, _05194_);
  and _49795_ (_05197_, _05121_, _35878_);
  and _49796_ (_05198_, _05197_, _35815_);
  not _49797_ (_05199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  nor _49798_ (_05200_, _05197_, _05199_);
  or _49799_ (_38200_, _05200_, _05198_);
  and _49800_ (_05201_, _05197_, _35822_);
  not _49801_ (_05202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  nor _49802_ (_05203_, _05197_, _05202_);
  or _49803_ (_38201_, _05203_, _05201_);
  and _49804_ (_05204_, _05197_, _35826_);
  not _49805_ (_05205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  nor _49806_ (_05206_, _05197_, _05205_);
  or _49807_ (_38202_, _05206_, _05204_);
  and _49808_ (_05207_, _05197_, _35830_);
  not _49809_ (_05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  nor _49810_ (_05209_, _05197_, _05208_);
  or _49811_ (_38203_, _05209_, _05207_);
  and _49812_ (_05210_, _05197_, _35834_);
  not _49813_ (_05211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  nor _49814_ (_05212_, _05197_, _05211_);
  or _49815_ (_38204_, _05212_, _05210_);
  and _49816_ (_05213_, _05197_, _35838_);
  not _49817_ (_05214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  nor _49818_ (_05215_, _05197_, _05214_);
  or _49819_ (_38205_, _05215_, _05213_);
  and _49820_ (_05216_, _05197_, _35842_);
  not _49821_ (_05217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  nor _49822_ (_05218_, _05197_, _05217_);
  or _49823_ (_38206_, _05218_, _05216_);
  and _49824_ (_05219_, _05197_, _35846_);
  not _49825_ (_05220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  nor _49826_ (_05221_, _05197_, _05220_);
  or _49827_ (_38207_, _05221_, _05219_);
  and _49828_ (_05222_, _05121_, _35905_);
  and _49829_ (_05223_, _05222_, _35815_);
  not _49830_ (_05224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  nor _49831_ (_05225_, _05222_, _05224_);
  or _49832_ (_38208_, _05225_, _05223_);
  and _49833_ (_05226_, _05222_, _35822_);
  not _49834_ (_05227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  nor _49835_ (_05228_, _05222_, _05227_);
  or _49836_ (_38209_, _05228_, _05226_);
  and _49837_ (_05229_, _05222_, _35826_);
  not _49838_ (_05230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  nor _49839_ (_05231_, _05222_, _05230_);
  or _49840_ (_38210_, _05231_, _05229_);
  and _49841_ (_05232_, _05222_, _35830_);
  not _49842_ (_05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  nor _49843_ (_05234_, _05222_, _05233_);
  or _49844_ (_38211_, _05234_, _05232_);
  and _49845_ (_05235_, _05222_, _35834_);
  not _49846_ (_05236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  nor _49847_ (_05237_, _05222_, _05236_);
  or _49848_ (_38212_, _05237_, _05235_);
  and _49849_ (_05238_, _05222_, _35838_);
  not _49850_ (_05239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  nor _49851_ (_05240_, _05222_, _05239_);
  or _49852_ (_38213_, _05240_, _05238_);
  and _49853_ (_05241_, _05222_, _35842_);
  not _49854_ (_05242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  nor _49855_ (_05243_, _05222_, _05242_);
  or _49856_ (_38214_, _05243_, _05241_);
  and _49857_ (_05244_, _05222_, _35846_);
  not _49858_ (_05245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  nor _49859_ (_05246_, _05222_, _05245_);
  or _49860_ (_38215_, _05246_, _05244_);
  and _49861_ (_05247_, _05121_, _35931_);
  and _49862_ (_05248_, _05247_, _35815_);
  not _49863_ (_05249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  nor _49864_ (_05250_, _05247_, _05249_);
  or _49865_ (_38216_, _05250_, _05248_);
  and _49866_ (_05251_, _05247_, _35822_);
  not _49867_ (_05252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  nor _49868_ (_05253_, _05247_, _05252_);
  or _49869_ (_38217_, _05253_, _05251_);
  and _49870_ (_05254_, _05247_, _35826_);
  not _49871_ (_05255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  nor _49872_ (_05256_, _05247_, _05255_);
  or _49873_ (_38218_, _05256_, _05254_);
  and _49874_ (_05257_, _05247_, _35830_);
  not _49875_ (_05258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  nor _49876_ (_05259_, _05247_, _05258_);
  or _49877_ (_38219_, _05259_, _05257_);
  and _49878_ (_05260_, _05247_, _35834_);
  not _49879_ (_05261_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  nor _49880_ (_05262_, _05247_, _05261_);
  or _49881_ (_38220_, _05262_, _05260_);
  and _49882_ (_05263_, _05247_, _35838_);
  not _49883_ (_05264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  nor _49884_ (_05265_, _05247_, _05264_);
  or _49885_ (_38221_, _05265_, _05263_);
  and _49886_ (_05266_, _05247_, _35842_);
  not _49887_ (_05267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  nor _49888_ (_05268_, _05247_, _05267_);
  or _49889_ (_38222_, _05268_, _05266_);
  and _49890_ (_05269_, _05247_, _35846_);
  not _49891_ (_05270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  nor _49892_ (_05271_, _05247_, _05270_);
  or _49893_ (_38223_, _05271_, _05269_);
  and _49894_ (_05272_, _05121_, _35957_);
  and _49895_ (_05273_, _05272_, _35815_);
  not _49896_ (_05274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  nor _49897_ (_05275_, _05272_, _05274_);
  or _49898_ (_38224_, _05275_, _05273_);
  and _49899_ (_05276_, _05272_, _35822_);
  not _49900_ (_05277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  nor _49901_ (_05278_, _05272_, _05277_);
  or _49902_ (_38225_, _05278_, _05276_);
  and _49903_ (_05279_, _05272_, _35826_);
  not _49904_ (_05280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  nor _49905_ (_05281_, _05272_, _05280_);
  or _49906_ (_38226_, _05281_, _05279_);
  and _49907_ (_05282_, _05272_, _35830_);
  not _49908_ (_05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  nor _49909_ (_05284_, _05272_, _05283_);
  or _49910_ (_38227_, _05284_, _05282_);
  and _49911_ (_05285_, _05272_, _35834_);
  not _49912_ (_05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  nor _49913_ (_05287_, _05272_, _05286_);
  or _49914_ (_38228_, _05287_, _05285_);
  and _49915_ (_05288_, _05272_, _35838_);
  not _49916_ (_05289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  nor _49917_ (_05290_, _05272_, _05289_);
  or _49918_ (_38229_, _05290_, _05288_);
  and _49919_ (_05291_, _05272_, _35842_);
  not _49920_ (_05292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  nor _49921_ (_05293_, _05272_, _05292_);
  or _49922_ (_38230_, _05293_, _05291_);
  and _49923_ (_05294_, _05272_, _35846_);
  not _49924_ (_05295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  nor _49925_ (_05296_, _05272_, _05295_);
  or _49926_ (_38231_, _05296_, _05294_);
  and _49927_ (_05297_, _05121_, _35983_);
  and _49928_ (_05298_, _05297_, _35815_);
  not _49929_ (_05299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  nor _49930_ (_05300_, _05297_, _05299_);
  or _49931_ (_38232_, _05300_, _05298_);
  and _49932_ (_05301_, _05297_, _35822_);
  not _49933_ (_05302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  nor _49934_ (_05303_, _05297_, _05302_);
  or _49935_ (_38233_, _05303_, _05301_);
  and _49936_ (_05304_, _05297_, _35826_);
  not _49937_ (_05305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  nor _49938_ (_05306_, _05297_, _05305_);
  or _49939_ (_38234_, _05306_, _05304_);
  and _49940_ (_05307_, _05297_, _35830_);
  not _49941_ (_05308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  nor _49942_ (_05309_, _05297_, _05308_);
  or _49943_ (_38235_, _05309_, _05307_);
  and _49944_ (_05310_, _05297_, _35834_);
  not _49945_ (_05311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  nor _49946_ (_05312_, _05297_, _05311_);
  or _49947_ (_38236_, _05312_, _05310_);
  and _49948_ (_05313_, _05297_, _35838_);
  not _49949_ (_05314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  nor _49950_ (_05315_, _05297_, _05314_);
  or _49951_ (_38237_, _05315_, _05313_);
  and _49952_ (_05316_, _05297_, _35842_);
  not _49953_ (_05317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  nor _49954_ (_05318_, _05297_, _05317_);
  or _49955_ (_38238_, _05318_, _05316_);
  and _49956_ (_05319_, _05297_, _35846_);
  not _49957_ (_05320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  nor _49958_ (_05321_, _05297_, _05320_);
  or _49959_ (_38239_, _05321_, _05319_);
  and _49960_ (_05322_, _05121_, _36010_);
  and _49961_ (_05323_, _05322_, _35815_);
  not _49962_ (_05324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  nor _49963_ (_05325_, _05322_, _05324_);
  or _49964_ (_38240_, _05325_, _05323_);
  and _49965_ (_05326_, _05322_, _35822_);
  not _49966_ (_05327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  nor _49967_ (_05328_, _05322_, _05327_);
  or _49968_ (_38241_, _05328_, _05326_);
  and _49969_ (_05329_, _05322_, _35826_);
  not _49970_ (_05330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  nor _49971_ (_05331_, _05322_, _05330_);
  or _49972_ (_38242_, _05331_, _05329_);
  and _49973_ (_05332_, _05322_, _35830_);
  not _49974_ (_05333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  nor _49975_ (_05334_, _05322_, _05333_);
  or _49976_ (_38243_, _05334_, _05332_);
  and _49977_ (_05335_, _05322_, _35834_);
  not _49978_ (_05336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  nor _49979_ (_05337_, _05322_, _05336_);
  or _49980_ (_38244_, _05337_, _05335_);
  and _49981_ (_05338_, _05322_, _35838_);
  not _49982_ (_05339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  nor _49983_ (_05340_, _05322_, _05339_);
  or _49984_ (_38245_, _05340_, _05338_);
  and _49985_ (_05341_, _05322_, _35842_);
  not _49986_ (_05342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  nor _49987_ (_05343_, _05322_, _05342_);
  or _49988_ (_38246_, _05343_, _05341_);
  and _49989_ (_05344_, _05322_, _35846_);
  not _49990_ (_05345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  nor _49991_ (_05346_, _05322_, _05345_);
  or _49992_ (_38247_, _05346_, _05344_);
  and _49993_ (_05347_, _05121_, _36036_);
  and _49994_ (_05348_, _05347_, _35815_);
  not _49995_ (_05349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  nor _49996_ (_05350_, _05347_, _05349_);
  or _49997_ (_38248_, _05350_, _05348_);
  and _49998_ (_05351_, _05347_, _35822_);
  not _49999_ (_05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  nor _50000_ (_05353_, _05347_, _05352_);
  or _50001_ (_38249_, _05353_, _05351_);
  and _50002_ (_05354_, _05347_, _35826_);
  not _50003_ (_05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  nor _50004_ (_05356_, _05347_, _05355_);
  or _50005_ (_38250_, _05356_, _05354_);
  and _50006_ (_05357_, _05347_, _35830_);
  not _50007_ (_05358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  nor _50008_ (_05359_, _05347_, _05358_);
  or _50009_ (_38251_, _05359_, _05357_);
  and _50010_ (_05360_, _05347_, _35834_);
  not _50011_ (_05361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  nor _50012_ (_05362_, _05347_, _05361_);
  or _50013_ (_38252_, _05362_, _05360_);
  and _50014_ (_05363_, _05347_, _35838_);
  not _50015_ (_05364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  nor _50016_ (_05365_, _05347_, _05364_);
  or _50017_ (_38253_, _05365_, _05363_);
  and _50018_ (_05366_, _05347_, _35842_);
  not _50019_ (_05367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  nor _50020_ (_05368_, _05347_, _05367_);
  or _50021_ (_38254_, _05368_, _05366_);
  and _50022_ (_05369_, _05347_, _35846_);
  not _50023_ (_05370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  nor _50024_ (_05371_, _05347_, _05370_);
  or _50025_ (_38255_, _05371_, _05369_);
  and _50026_ (_05372_, _05121_, _36062_);
  and _50027_ (_05373_, _05372_, _35815_);
  not _50028_ (_05374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  nor _50029_ (_05375_, _05372_, _05374_);
  or _50030_ (_38264_, _05375_, _05373_);
  and _50031_ (_05376_, _05372_, _35822_);
  not _50032_ (_05377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  nor _50033_ (_05378_, _05372_, _05377_);
  or _50034_ (_38265_, _05378_, _05376_);
  and _50035_ (_05379_, _05372_, _35826_);
  not _50036_ (_05380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  nor _50037_ (_05381_, _05372_, _05380_);
  or _50038_ (_38266_, _05381_, _05379_);
  and _50039_ (_05382_, _05372_, _35830_);
  not _50040_ (_05383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  nor _50041_ (_05384_, _05372_, _05383_);
  or _50042_ (_38267_, _05384_, _05382_);
  and _50043_ (_05385_, _05372_, _35834_);
  not _50044_ (_05386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  nor _50045_ (_05387_, _05372_, _05386_);
  or _50046_ (_38268_, _05387_, _05385_);
  and _50047_ (_05388_, _05372_, _35838_);
  not _50048_ (_05389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  nor _50049_ (_05390_, _05372_, _05389_);
  or _50050_ (_38269_, _05390_, _05388_);
  and _50051_ (_05391_, _05372_, _35842_);
  not _50052_ (_05392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  nor _50053_ (_05393_, _05372_, _05392_);
  or _50054_ (_38270_, _05393_, _05391_);
  and _50055_ (_05394_, _05372_, _35846_);
  not _50056_ (_05395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  nor _50057_ (_05396_, _05372_, _05395_);
  or _50058_ (_38271_, _05396_, _05394_);
  and _50059_ (_05397_, _05121_, _36088_);
  and _50060_ (_05398_, _05397_, _35815_);
  not _50061_ (_05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  nor _50062_ (_05400_, _05397_, _05399_);
  or _50063_ (_38272_, _05400_, _05398_);
  and _50064_ (_05401_, _05397_, _35822_);
  not _50065_ (_05402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  nor _50066_ (_05403_, _05397_, _05402_);
  or _50067_ (_38273_, _05403_, _05401_);
  and _50068_ (_05404_, _05397_, _35826_);
  not _50069_ (_05405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  nor _50070_ (_05406_, _05397_, _05405_);
  or _50071_ (_38274_, _05406_, _05404_);
  and _50072_ (_05407_, _05397_, _35830_);
  not _50073_ (_05408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  nor _50074_ (_05409_, _05397_, _05408_);
  or _50075_ (_38275_, _05409_, _05407_);
  and _50076_ (_05410_, _05397_, _35834_);
  not _50077_ (_05411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  nor _50078_ (_05412_, _05397_, _05411_);
  or _50079_ (_38276_, _05412_, _05410_);
  and _50080_ (_05413_, _05397_, _35838_);
  not _50081_ (_05414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  nor _50082_ (_05415_, _05397_, _05414_);
  or _50083_ (_38277_, _05415_, _05413_);
  and _50084_ (_05416_, _05397_, _35842_);
  not _50085_ (_05417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  nor _50086_ (_05418_, _05397_, _05417_);
  or _50087_ (_38278_, _05418_, _05416_);
  and _50088_ (_05419_, _05397_, _35846_);
  not _50089_ (_05420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  nor _50090_ (_05421_, _05397_, _05420_);
  or _50091_ (_38279_, _05421_, _05419_);
  and _50092_ (_05422_, _05121_, _36115_);
  and _50093_ (_05423_, _05422_, _35815_);
  not _50094_ (_05424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  nor _50095_ (_05425_, _05422_, _05424_);
  or _50096_ (_38280_, _05425_, _05423_);
  and _50097_ (_05426_, _05422_, _35822_);
  not _50098_ (_05427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  nor _50099_ (_05428_, _05422_, _05427_);
  or _50100_ (_38281_, _05428_, _05426_);
  and _50101_ (_05429_, _05422_, _35826_);
  not _50102_ (_05430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  nor _50103_ (_05431_, _05422_, _05430_);
  or _50104_ (_38282_, _05431_, _05429_);
  and _50105_ (_05432_, _05422_, _35830_);
  not _50106_ (_05433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  nor _50107_ (_05434_, _05422_, _05433_);
  or _50108_ (_38283_, _05434_, _05432_);
  and _50109_ (_05435_, _05422_, _35834_);
  not _50110_ (_05436_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  nor _50111_ (_05437_, _05422_, _05436_);
  or _50112_ (_38284_, _05437_, _05435_);
  and _50113_ (_05438_, _05422_, _35838_);
  not _50114_ (_05439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  nor _50115_ (_05440_, _05422_, _05439_);
  or _50116_ (_38285_, _05440_, _05438_);
  and _50117_ (_05441_, _05422_, _35842_);
  not _50118_ (_05442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  nor _50119_ (_05443_, _05422_, _05442_);
  or _50120_ (_38286_, _05443_, _05441_);
  and _50121_ (_05444_, _05422_, _35846_);
  not _50122_ (_05445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  nor _50123_ (_05446_, _05422_, _05445_);
  or _50124_ (_38287_, _05446_, _05444_);
  and _50125_ (_05447_, _05121_, _36141_);
  and _50126_ (_05448_, _05447_, _35815_);
  not _50127_ (_05449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  nor _50128_ (_05450_, _05447_, _05449_);
  or _50129_ (_38288_, _05450_, _05448_);
  and _50130_ (_05451_, _05447_, _35822_);
  not _50131_ (_05452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  nor _50132_ (_05453_, _05447_, _05452_);
  or _50133_ (_38289_, _05453_, _05451_);
  and _50134_ (_05454_, _05447_, _35826_);
  not _50135_ (_05455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  nor _50136_ (_05456_, _05447_, _05455_);
  or _50137_ (_38290_, _05456_, _05454_);
  and _50138_ (_05457_, _05447_, _35830_);
  not _50139_ (_05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  nor _50140_ (_05459_, _05447_, _05458_);
  or _50141_ (_38291_, _05459_, _05457_);
  and _50142_ (_05460_, _05447_, _35834_);
  not _50143_ (_05461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  nor _50144_ (_05462_, _05447_, _05461_);
  or _50145_ (_38292_, _05462_, _05460_);
  and _50146_ (_05463_, _05447_, _35838_);
  not _50147_ (_05464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  nor _50148_ (_05465_, _05447_, _05464_);
  or _50149_ (_38293_, _05465_, _05463_);
  and _50150_ (_05466_, _05447_, _35842_);
  not _50151_ (_05467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  nor _50152_ (_05468_, _05447_, _05467_);
  or _50153_ (_38294_, _05468_, _05466_);
  and _50154_ (_05469_, _05447_, _35846_);
  not _50155_ (_05470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  nor _50156_ (_05471_, _05447_, _05470_);
  or _50157_ (_38295_, _05471_, _05469_);
  and _50158_ (_05472_, _05121_, _36167_);
  and _50159_ (_05473_, _05472_, _35815_);
  not _50160_ (_05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  nor _50161_ (_05475_, _05472_, _05474_);
  or _50162_ (_38296_, _05475_, _05473_);
  and _50163_ (_05476_, _05472_, _35822_);
  not _50164_ (_05477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  nor _50165_ (_05478_, _05472_, _05477_);
  or _50166_ (_38297_, _05478_, _05476_);
  and _50167_ (_05479_, _05472_, _35826_);
  not _50168_ (_05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  nor _50169_ (_05481_, _05472_, _05480_);
  or _50170_ (_38298_, _05481_, _05479_);
  and _50171_ (_05482_, _05472_, _35830_);
  not _50172_ (_05483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  nor _50173_ (_05484_, _05472_, _05483_);
  or _50174_ (_38299_, _05484_, _05482_);
  and _50175_ (_05485_, _05472_, _35834_);
  not _50176_ (_05486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  nor _50177_ (_05487_, _05472_, _05486_);
  or _50178_ (_38300_, _05487_, _05485_);
  and _50179_ (_05488_, _05472_, _35838_);
  not _50180_ (_05489_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  nor _50181_ (_05490_, _05472_, _05489_);
  or _50182_ (_38301_, _05490_, _05488_);
  and _50183_ (_05491_, _05472_, _35842_);
  not _50184_ (_05492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  nor _50185_ (_05493_, _05472_, _05492_);
  or _50186_ (_38302_, _05493_, _05491_);
  and _50187_ (_05494_, _05472_, _35846_);
  not _50188_ (_05495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  nor _50189_ (_05496_, _05472_, _05495_);
  or _50190_ (_38303_, _05496_, _05494_);
  and _50191_ (_05497_, _05121_, _36193_);
  and _50192_ (_05498_, _05497_, _35815_);
  not _50193_ (_05499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  nor _50194_ (_05500_, _05497_, _05499_);
  or _50195_ (_38304_, _05500_, _05498_);
  and _50196_ (_05501_, _05497_, _35822_);
  not _50197_ (_05502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  nor _50198_ (_05503_, _05497_, _05502_);
  or _50199_ (_38305_, _05503_, _05501_);
  and _50200_ (_05504_, _05497_, _35826_);
  not _50201_ (_05505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  nor _50202_ (_05506_, _05497_, _05505_);
  or _50203_ (_38306_, _05506_, _05504_);
  and _50204_ (_05507_, _05497_, _35830_);
  not _50205_ (_05508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  nor _50206_ (_05509_, _05497_, _05508_);
  or _50207_ (_38307_, _05509_, _05507_);
  and _50208_ (_05510_, _05497_, _35834_);
  not _50209_ (_05511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  nor _50210_ (_05512_, _05497_, _05511_);
  or _50211_ (_38308_, _05512_, _05510_);
  and _50212_ (_05513_, _05497_, _35838_);
  not _50213_ (_05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  nor _50214_ (_05515_, _05497_, _05514_);
  or _50215_ (_38309_, _05515_, _05513_);
  and _50216_ (_05516_, _05497_, _35842_);
  not _50217_ (_05517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  nor _50218_ (_05518_, _05497_, _05517_);
  or _50219_ (_38310_, _05518_, _05516_);
  and _50220_ (_05519_, _05497_, _35846_);
  not _50221_ (_05520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  nor _50222_ (_05521_, _05497_, _05520_);
  or _50223_ (_38311_, _05521_, _05519_);
  and _50224_ (_05522_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and _50225_ (_05523_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or _50226_ (_05524_, _05523_, _05522_);
  and _50227_ (_05525_, _05524_, _34581_);
  and _50228_ (_05526_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and _50229_ (_05527_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or _50230_ (_05528_, _05527_, _05526_);
  and _50231_ (_05529_, _05528_, _34796_);
  or _50232_ (_05530_, _05529_, _05525_);
  and _50233_ (_05531_, _05530_, _34772_);
  and _50234_ (_05532_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and _50235_ (_05533_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or _50236_ (_05534_, _05533_, _05532_);
  and _50237_ (_05535_, _05534_, _34581_);
  and _50238_ (_05536_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and _50239_ (_05537_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or _50240_ (_05538_, _05537_, _05536_);
  and _50241_ (_05539_, _05538_, _34796_);
  or _50242_ (_05540_, _05539_, _05535_);
  and _50243_ (_05541_, _05540_, _34790_);
  or _50244_ (_05542_, _05541_, _34719_);
  or _50245_ (_05543_, _05542_, _05531_);
  or _50246_ (_05544_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or _50247_ (_05545_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and _50248_ (_05546_, _05545_, _34796_);
  and _50249_ (_05547_, _05546_, _05544_);
  or _50250_ (_05548_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or _50251_ (_05549_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and _50252_ (_05550_, _05549_, _34581_);
  and _50253_ (_05551_, _05550_, _05548_);
  or _50254_ (_05552_, _05551_, _05547_);
  and _50255_ (_05553_, _05552_, _34772_);
  or _50256_ (_05554_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or _50257_ (_05555_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and _50258_ (_05556_, _05555_, _34796_);
  and _50259_ (_05557_, _05556_, _05554_);
  or _50260_ (_05558_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or _50261_ (_05559_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and _50262_ (_05560_, _05559_, _34581_);
  and _50263_ (_05561_, _05560_, _05558_);
  or _50264_ (_05562_, _05561_, _05557_);
  and _50265_ (_05563_, _05562_, _34790_);
  or _50266_ (_05564_, _05563_, _34803_);
  or _50267_ (_05565_, _05564_, _05553_);
  and _50268_ (_05566_, _05565_, _05543_);
  or _50269_ (_05567_, _05566_, _34700_);
  and _50270_ (_05568_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and _50271_ (_05569_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or _50272_ (_05570_, _05569_, _05568_);
  and _50273_ (_05571_, _05570_, _34581_);
  and _50274_ (_05572_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and _50275_ (_05573_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or _50276_ (_05574_, _05573_, _05572_);
  and _50277_ (_05575_, _05574_, _34796_);
  or _50278_ (_05576_, _05575_, _05571_);
  and _50279_ (_05577_, _05576_, _34772_);
  and _50280_ (_05578_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and _50281_ (_05579_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or _50282_ (_05580_, _05579_, _05578_);
  and _50283_ (_05581_, _05580_, _34581_);
  and _50284_ (_05582_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and _50285_ (_05583_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or _50286_ (_05584_, _05583_, _05582_);
  and _50287_ (_05585_, _05584_, _34796_);
  or _50288_ (_05586_, _05585_, _05581_);
  and _50289_ (_05587_, _05586_, _34790_);
  or _50290_ (_05588_, _05587_, _34719_);
  or _50291_ (_05589_, _05588_, _05577_);
  or _50292_ (_05590_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or _50293_ (_05591_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and _50294_ (_05592_, _05591_, _05590_);
  and _50295_ (_05593_, _05592_, _34581_);
  or _50296_ (_05594_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or _50297_ (_05595_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and _50298_ (_05596_, _05595_, _05594_);
  and _50299_ (_05597_, _05596_, _34796_);
  or _50300_ (_05598_, _05597_, _05593_);
  and _50301_ (_05599_, _05598_, _34772_);
  or _50302_ (_05600_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or _50303_ (_05601_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and _50304_ (_05602_, _05601_, _05600_);
  and _50305_ (_05603_, _05602_, _34581_);
  or _50306_ (_05604_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or _50307_ (_05605_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and _50308_ (_05606_, _05605_, _05604_);
  and _50309_ (_05607_, _05606_, _34796_);
  or _50310_ (_05608_, _05607_, _05603_);
  and _50311_ (_05609_, _05608_, _34790_);
  or _50312_ (_05610_, _05609_, _34803_);
  or _50313_ (_05611_, _05610_, _05599_);
  and _50314_ (_05612_, _05611_, _05589_);
  or _50315_ (_05613_, _05612_, _34789_);
  and _50316_ (_05614_, _05613_, _34638_);
  and _50317_ (_05615_, _05614_, _05567_);
  and _50318_ (_05616_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and _50319_ (_05617_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or _50320_ (_05618_, _05617_, _05616_);
  and _50321_ (_05619_, _05618_, _34581_);
  and _50322_ (_05620_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and _50323_ (_05621_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or _50324_ (_05622_, _05621_, _05620_);
  and _50325_ (_05623_, _05622_, _34796_);
  or _50326_ (_05624_, _05623_, _05619_);
  or _50327_ (_05625_, _05624_, _34790_);
  and _50328_ (_05626_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and _50329_ (_05627_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or _50330_ (_05628_, _05627_, _05626_);
  and _50331_ (_05629_, _05628_, _34581_);
  and _50332_ (_05630_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and _50333_ (_05631_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or _50334_ (_05632_, _05631_, _05630_);
  and _50335_ (_05633_, _05632_, _34796_);
  or _50336_ (_05634_, _05633_, _05629_);
  or _50337_ (_05635_, _05634_, _34772_);
  and _50338_ (_05636_, _05635_, _34803_);
  and _50339_ (_05637_, _05636_, _05625_);
  or _50340_ (_05638_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or _50341_ (_05639_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and _50342_ (_05640_, _05639_, _05638_);
  and _50343_ (_05641_, _05640_, _34581_);
  or _50344_ (_05642_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or _50345_ (_05643_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and _50346_ (_05644_, _05643_, _05642_);
  and _50347_ (_05645_, _05644_, _34796_);
  or _50348_ (_05646_, _05645_, _05641_);
  or _50349_ (_05647_, _05646_, _34790_);
  or _50350_ (_05648_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or _50351_ (_05649_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and _50352_ (_05650_, _05649_, _05648_);
  and _50353_ (_05651_, _05650_, _34581_);
  or _50354_ (_05652_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or _50355_ (_05653_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and _50356_ (_05654_, _05653_, _05652_);
  and _50357_ (_05655_, _05654_, _34796_);
  or _50358_ (_05656_, _05655_, _05651_);
  or _50359_ (_05657_, _05656_, _34772_);
  and _50360_ (_05658_, _05657_, _34719_);
  and _50361_ (_05659_, _05658_, _05647_);
  or _50362_ (_05660_, _05659_, _05637_);
  or _50363_ (_05661_, _05660_, _34789_);
  and _50364_ (_05662_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and _50365_ (_05663_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or _50366_ (_05664_, _05663_, _05662_);
  and _50367_ (_05665_, _05664_, _34581_);
  and _50368_ (_05666_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and _50369_ (_05667_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or _50370_ (_05668_, _05667_, _05666_);
  and _50371_ (_05669_, _05668_, _34796_);
  or _50372_ (_05670_, _05669_, _05665_);
  or _50373_ (_05671_, _05670_, _34790_);
  and _50374_ (_05672_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and _50375_ (_05673_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or _50376_ (_05674_, _05673_, _05672_);
  and _50377_ (_05675_, _05674_, _34581_);
  and _50378_ (_05676_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and _50379_ (_05677_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or _50380_ (_05678_, _05677_, _05676_);
  and _50381_ (_05679_, _05678_, _34796_);
  or _50382_ (_05680_, _05679_, _05675_);
  or _50383_ (_05681_, _05680_, _34772_);
  and _50384_ (_05682_, _05681_, _34803_);
  and _50385_ (_05683_, _05682_, _05671_);
  or _50386_ (_05684_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or _50387_ (_05685_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and _50388_ (_05686_, _05685_, _34796_);
  and _50389_ (_05687_, _05686_, _05684_);
  or _50390_ (_05688_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or _50391_ (_05689_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and _50392_ (_05690_, _05689_, _34581_);
  and _50393_ (_05691_, _05690_, _05688_);
  or _50394_ (_05692_, _05691_, _05687_);
  or _50395_ (_05693_, _05692_, _34790_);
  or _50396_ (_05694_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or _50397_ (_05695_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and _50398_ (_05696_, _05695_, _34796_);
  and _50399_ (_05697_, _05696_, _05694_);
  or _50400_ (_05698_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or _50401_ (_05699_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and _50402_ (_05700_, _05699_, _34581_);
  and _50403_ (_05701_, _05700_, _05698_);
  or _50404_ (_05702_, _05701_, _05697_);
  or _50405_ (_05703_, _05702_, _34772_);
  and _50406_ (_05704_, _05703_, _34719_);
  and _50407_ (_05705_, _05704_, _05693_);
  or _50408_ (_05706_, _05705_, _05683_);
  or _50409_ (_05707_, _05706_, _34700_);
  and _50410_ (_05708_, _05707_, _34840_);
  and _50411_ (_05709_, _05708_, _05661_);
  or _50412_ (_05710_, _05709_, _05615_);
  or _50413_ (_05711_, _05710_, _34692_);
  and _50414_ (_05712_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and _50415_ (_05713_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or _50416_ (_05714_, _05713_, _05712_);
  and _50417_ (_05715_, _05714_, _34581_);
  and _50418_ (_05716_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and _50419_ (_05717_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or _50420_ (_05718_, _05717_, _05716_);
  and _50421_ (_05719_, _05718_, _34796_);
  or _50422_ (_05720_, _05719_, _05715_);
  and _50423_ (_05721_, _05720_, _34790_);
  and _50424_ (_05722_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and _50425_ (_05723_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or _50426_ (_05724_, _05723_, _05722_);
  and _50427_ (_05725_, _05724_, _34581_);
  and _50428_ (_05726_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and _50429_ (_05727_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or _50430_ (_05728_, _05727_, _05726_);
  and _50431_ (_05729_, _05728_, _34796_);
  or _50432_ (_05730_, _05729_, _05725_);
  and _50433_ (_05731_, _05730_, _34772_);
  or _50434_ (_05732_, _05731_, _05721_);
  and _50435_ (_05733_, _05732_, _34803_);
  or _50436_ (_05734_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or _50437_ (_05735_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and _50438_ (_05736_, _05735_, _05734_);
  and _50439_ (_05737_, _05736_, _34581_);
  or _50440_ (_05738_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or _50441_ (_05739_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and _50442_ (_05740_, _05739_, _05738_);
  and _50443_ (_05741_, _05740_, _34796_);
  or _50444_ (_05742_, _05741_, _05737_);
  and _50445_ (_05743_, _05742_, _34790_);
  or _50446_ (_05744_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or _50447_ (_05745_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and _50448_ (_05746_, _05745_, _05744_);
  and _50449_ (_05747_, _05746_, _34581_);
  or _50450_ (_05748_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or _50451_ (_05749_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and _50452_ (_05750_, _05749_, _05748_);
  and _50453_ (_05751_, _05750_, _34796_);
  or _50454_ (_05752_, _05751_, _05747_);
  and _50455_ (_05753_, _05752_, _34772_);
  or _50456_ (_05754_, _05753_, _05743_);
  and _50457_ (_05755_, _05754_, _34719_);
  or _50458_ (_05756_, _05755_, _05733_);
  or _50459_ (_05757_, _05756_, _34789_);
  and _50460_ (_05758_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  and _50461_ (_05759_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or _50462_ (_05760_, _05759_, _05758_);
  and _50463_ (_05761_, _05760_, _34581_);
  and _50464_ (_05762_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  and _50465_ (_05763_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or _50466_ (_05764_, _05763_, _05762_);
  and _50467_ (_05765_, _05764_, _34796_);
  or _50468_ (_05766_, _05765_, _05761_);
  and _50469_ (_05767_, _05766_, _34790_);
  and _50470_ (_05768_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and _50471_ (_05769_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or _50472_ (_05770_, _05769_, _05768_);
  and _50473_ (_05771_, _05770_, _34581_);
  and _50474_ (_05772_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  and _50475_ (_05773_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or _50476_ (_05774_, _05773_, _05772_);
  and _50477_ (_05775_, _05774_, _34796_);
  or _50478_ (_05776_, _05775_, _05771_);
  and _50479_ (_05777_, _05776_, _34772_);
  or _50480_ (_05778_, _05777_, _05767_);
  and _50481_ (_05779_, _05778_, _34803_);
  or _50482_ (_05780_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or _50483_ (_05781_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  and _50484_ (_05782_, _05781_, _34796_);
  and _50485_ (_05783_, _05782_, _05780_);
  or _50486_ (_05784_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or _50487_ (_05785_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  and _50488_ (_05786_, _05785_, _34581_);
  and _50489_ (_05787_, _05786_, _05784_);
  or _50490_ (_05788_, _05787_, _05783_);
  and _50491_ (_05789_, _05788_, _34790_);
  or _50492_ (_05790_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or _50493_ (_05791_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and _50494_ (_05792_, _05791_, _34796_);
  and _50495_ (_05793_, _05792_, _05790_);
  or _50496_ (_05794_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or _50497_ (_05795_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  and _50498_ (_05796_, _05795_, _34581_);
  and _50499_ (_05797_, _05796_, _05794_);
  or _50500_ (_05798_, _05797_, _05793_);
  and _50501_ (_05799_, _05798_, _34772_);
  or _50502_ (_05800_, _05799_, _05789_);
  and _50503_ (_05801_, _05800_, _34719_);
  or _50504_ (_05802_, _05801_, _05779_);
  or _50505_ (_05803_, _05802_, _34700_);
  and _50506_ (_05804_, _05803_, _34638_);
  and _50507_ (_05805_, _05804_, _05757_);
  and _50508_ (_05806_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and _50509_ (_05807_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or _50510_ (_05808_, _05807_, _05806_);
  and _50511_ (_05809_, _05808_, _34581_);
  and _50512_ (_05810_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and _50513_ (_05811_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or _50514_ (_05812_, _05811_, _05810_);
  and _50515_ (_05813_, _05812_, _34796_);
  or _50516_ (_05814_, _05813_, _05809_);
  or _50517_ (_05815_, _05814_, _34790_);
  and _50518_ (_05816_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and _50519_ (_05817_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or _50520_ (_05818_, _05817_, _05816_);
  and _50521_ (_05819_, _05818_, _34581_);
  and _50522_ (_05820_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and _50523_ (_05821_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or _50524_ (_05822_, _05821_, _05820_);
  and _50525_ (_05823_, _05822_, _34796_);
  or _50526_ (_05824_, _05823_, _05819_);
  or _50527_ (_05825_, _05824_, _34772_);
  and _50528_ (_05826_, _05825_, _34803_);
  and _50529_ (_05827_, _05826_, _05815_);
  or _50530_ (_05828_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or _50531_ (_05829_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and _50532_ (_05830_, _05829_, _34796_);
  and _50533_ (_05831_, _05830_, _05828_);
  or _50534_ (_05832_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or _50535_ (_05833_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and _50536_ (_05834_, _05833_, _34581_);
  and _50537_ (_05835_, _05834_, _05832_);
  or _50538_ (_05836_, _05835_, _05831_);
  or _50539_ (_05837_, _05836_, _34790_);
  or _50540_ (_05838_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or _50541_ (_05839_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and _50542_ (_05840_, _05839_, _34796_);
  and _50543_ (_05841_, _05840_, _05838_);
  or _50544_ (_05842_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or _50545_ (_05843_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and _50546_ (_05844_, _05843_, _34581_);
  and _50547_ (_05845_, _05844_, _05842_);
  or _50548_ (_05846_, _05845_, _05841_);
  or _50549_ (_05847_, _05846_, _34772_);
  and _50550_ (_05848_, _05847_, _34719_);
  and _50551_ (_05849_, _05848_, _05837_);
  or _50552_ (_05850_, _05849_, _05827_);
  or _50553_ (_05851_, _05850_, _34700_);
  and _50554_ (_05852_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and _50555_ (_05853_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or _50556_ (_05854_, _05853_, _05852_);
  and _50557_ (_05855_, _05854_, _34581_);
  and _50558_ (_05856_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and _50559_ (_05857_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or _50560_ (_05858_, _05857_, _05856_);
  and _50561_ (_05859_, _05858_, _34796_);
  or _50562_ (_05860_, _05859_, _05855_);
  or _50563_ (_05861_, _05860_, _34790_);
  and _50564_ (_05862_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and _50565_ (_05863_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or _50566_ (_05864_, _05863_, _05862_);
  and _50567_ (_05865_, _05864_, _34581_);
  and _50568_ (_05866_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and _50569_ (_05867_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or _50570_ (_05868_, _05867_, _05866_);
  and _50571_ (_05869_, _05868_, _34796_);
  or _50572_ (_05870_, _05869_, _05865_);
  or _50573_ (_05871_, _05870_, _34772_);
  and _50574_ (_05872_, _05871_, _34803_);
  and _50575_ (_05873_, _05872_, _05861_);
  or _50576_ (_05874_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or _50577_ (_05875_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and _50578_ (_05876_, _05875_, _05874_);
  and _50579_ (_05877_, _05876_, _34581_);
  or _50580_ (_05878_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or _50581_ (_05879_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and _50582_ (_05880_, _05879_, _05878_);
  and _50583_ (_05881_, _05880_, _34796_);
  or _50584_ (_05882_, _05881_, _05877_);
  or _50585_ (_05883_, _05882_, _34790_);
  or _50586_ (_05884_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or _50587_ (_05885_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and _50588_ (_05886_, _05885_, _05884_);
  and _50589_ (_05887_, _05886_, _34581_);
  or _50590_ (_05888_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or _50591_ (_05889_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and _50592_ (_05890_, _05889_, _05888_);
  and _50593_ (_05891_, _05890_, _34796_);
  or _50594_ (_05892_, _05891_, _05887_);
  or _50595_ (_05893_, _05892_, _34772_);
  and _50596_ (_05894_, _05893_, _34719_);
  and _50597_ (_05895_, _05894_, _05883_);
  or _50598_ (_05896_, _05895_, _05873_);
  or _50599_ (_05897_, _05896_, _34789_);
  and _50600_ (_05898_, _05897_, _34840_);
  and _50601_ (_05899_, _05898_, _05851_);
  or _50602_ (_05900_, _05899_, _05805_);
  or _50603_ (_05901_, _05900_, _34985_);
  and _50604_ (_05902_, _05901_, _34346_);
  and _50605_ (_05903_, _05902_, _05711_);
  and _50606_ (_05904_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and _50607_ (_05905_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or _50608_ (_05906_, _05905_, _05904_);
  and _50609_ (_05907_, _05906_, _34581_);
  and _50610_ (_05908_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and _50611_ (_05909_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or _50612_ (_05910_, _05909_, _05908_);
  and _50613_ (_05911_, _05910_, _34796_);
  or _50614_ (_05912_, _05911_, _05907_);
  or _50615_ (_05913_, _05912_, _34790_);
  and _50616_ (_05914_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and _50617_ (_05915_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or _50618_ (_05916_, _05915_, _05914_);
  and _50619_ (_05917_, _05916_, _34581_);
  and _50620_ (_05918_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and _50621_ (_05919_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or _50622_ (_05920_, _05919_, _05918_);
  and _50623_ (_05921_, _05920_, _34796_);
  or _50624_ (_05922_, _05921_, _05917_);
  or _50625_ (_05923_, _05922_, _34772_);
  and _50626_ (_05924_, _05923_, _34803_);
  and _50627_ (_05925_, _05924_, _05913_);
  or _50628_ (_05926_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or _50629_ (_05927_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and _50630_ (_05928_, _05927_, _05926_);
  and _50631_ (_05929_, _05928_, _34581_);
  or _50632_ (_05930_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or _50633_ (_05931_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and _50634_ (_05932_, _05931_, _05930_);
  and _50635_ (_05933_, _05932_, _34796_);
  or _50636_ (_05934_, _05933_, _05929_);
  or _50637_ (_05935_, _05934_, _34790_);
  or _50638_ (_05936_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or _50639_ (_05937_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and _50640_ (_05938_, _05937_, _05936_);
  and _50641_ (_05939_, _05938_, _34581_);
  or _50642_ (_05940_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or _50643_ (_05941_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and _50644_ (_05942_, _05941_, _05940_);
  and _50645_ (_05943_, _05942_, _34796_);
  or _50646_ (_05944_, _05943_, _05939_);
  or _50647_ (_05945_, _05944_, _34772_);
  and _50648_ (_05946_, _05945_, _34719_);
  and _50649_ (_05947_, _05946_, _05935_);
  or _50650_ (_05948_, _05947_, _05925_);
  and _50651_ (_05949_, _05948_, _34700_);
  and _50652_ (_05950_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and _50653_ (_05951_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or _50654_ (_05952_, _05951_, _05950_);
  and _50655_ (_05953_, _05952_, _34581_);
  and _50656_ (_05954_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and _50657_ (_05955_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or _50658_ (_05956_, _05955_, _05954_);
  and _50659_ (_05957_, _05956_, _34796_);
  or _50660_ (_05958_, _05957_, _05953_);
  or _50661_ (_05959_, _05958_, _34790_);
  and _50662_ (_05960_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and _50663_ (_05961_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or _50664_ (_05962_, _05961_, _05960_);
  and _50665_ (_05963_, _05962_, _34581_);
  and _50666_ (_05964_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and _50667_ (_05965_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or _50668_ (_05966_, _05965_, _05964_);
  and _50669_ (_05967_, _05966_, _34796_);
  or _50670_ (_05968_, _05967_, _05963_);
  or _50671_ (_05969_, _05968_, _34772_);
  and _50672_ (_05970_, _05969_, _34803_);
  and _50673_ (_05971_, _05970_, _05959_);
  or _50674_ (_05972_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or _50675_ (_05973_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  and _50676_ (_05974_, _05973_, _34796_);
  and _50677_ (_05975_, _05974_, _05972_);
  or _50678_ (_05976_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or _50679_ (_05977_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and _50680_ (_05978_, _05977_, _34581_);
  and _50681_ (_05979_, _05978_, _05976_);
  or _50682_ (_05980_, _05979_, _05975_);
  or _50683_ (_05981_, _05980_, _34790_);
  or _50684_ (_05982_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or _50685_ (_05983_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and _50686_ (_05984_, _05983_, _34796_);
  and _50687_ (_05985_, _05984_, _05982_);
  or _50688_ (_05986_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or _50689_ (_05987_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and _50690_ (_05988_, _05987_, _34581_);
  and _50691_ (_05989_, _05988_, _05986_);
  or _50692_ (_05990_, _05989_, _05985_);
  or _50693_ (_05991_, _05990_, _34772_);
  and _50694_ (_05992_, _05991_, _34719_);
  and _50695_ (_05993_, _05992_, _05981_);
  or _50696_ (_05994_, _05993_, _05971_);
  and _50697_ (_05995_, _05994_, _34789_);
  or _50698_ (_05996_, _05995_, _05949_);
  and _50699_ (_05997_, _05996_, _34840_);
  and _50700_ (_05998_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  and _50701_ (_05999_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or _50702_ (_06000_, _05999_, _05998_);
  and _50703_ (_06001_, _06000_, _34581_);
  and _50704_ (_06002_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and _50705_ (_06003_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or _50706_ (_06004_, _06003_, _06002_);
  and _50707_ (_06005_, _06004_, _34796_);
  or _50708_ (_06006_, _06005_, _06001_);
  and _50709_ (_06007_, _06006_, _34772_);
  and _50710_ (_06008_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and _50711_ (_06009_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or _50712_ (_06010_, _06009_, _06008_);
  and _50713_ (_06011_, _06010_, _34581_);
  and _50714_ (_06012_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and _50715_ (_06013_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or _50716_ (_06014_, _06013_, _06012_);
  and _50717_ (_06015_, _06014_, _34796_);
  or _50718_ (_06016_, _06015_, _06011_);
  and _50719_ (_06017_, _06016_, _34790_);
  or _50720_ (_06018_, _06017_, _06007_);
  and _50721_ (_06019_, _06018_, _34803_);
  or _50722_ (_06020_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or _50723_ (_06021_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and _50724_ (_06022_, _06021_, _34796_);
  and _50725_ (_06023_, _06022_, _06020_);
  or _50726_ (_06024_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or _50727_ (_06025_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  and _50728_ (_06026_, _06025_, _34581_);
  and _50729_ (_06027_, _06026_, _06024_);
  or _50730_ (_06028_, _06027_, _06023_);
  and _50731_ (_06029_, _06028_, _34772_);
  or _50732_ (_06030_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or _50733_ (_06031_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and _50734_ (_06032_, _06031_, _34796_);
  and _50735_ (_06033_, _06032_, _06030_);
  or _50736_ (_06034_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or _50737_ (_06035_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and _50738_ (_06036_, _06035_, _34581_);
  and _50739_ (_06037_, _06036_, _06034_);
  or _50740_ (_06038_, _06037_, _06033_);
  and _50741_ (_06039_, _06038_, _34790_);
  or _50742_ (_06040_, _06039_, _06029_);
  and _50743_ (_06041_, _06040_, _34719_);
  or _50744_ (_06042_, _06041_, _06019_);
  and _50745_ (_06043_, _06042_, _34789_);
  and _50746_ (_06044_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and _50747_ (_06045_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or _50748_ (_06046_, _06045_, _06044_);
  and _50749_ (_06047_, _06046_, _34581_);
  and _50750_ (_06048_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and _50751_ (_06049_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or _50752_ (_06050_, _06049_, _06048_);
  and _50753_ (_06051_, _06050_, _34796_);
  or _50754_ (_06052_, _06051_, _06047_);
  and _50755_ (_06053_, _06052_, _34772_);
  and _50756_ (_06054_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and _50757_ (_06055_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or _50758_ (_06056_, _06055_, _06054_);
  and _50759_ (_06057_, _06056_, _34581_);
  and _50760_ (_06058_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and _50761_ (_06059_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or _50762_ (_06060_, _06059_, _06058_);
  and _50763_ (_06061_, _06060_, _34796_);
  or _50764_ (_06062_, _06061_, _06057_);
  and _50765_ (_06063_, _06062_, _34790_);
  or _50766_ (_06064_, _06063_, _06053_);
  and _50767_ (_06065_, _06064_, _34803_);
  or _50768_ (_06066_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or _50769_ (_06067_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and _50770_ (_06068_, _06067_, _06066_);
  and _50771_ (_06069_, _06068_, _34581_);
  or _50772_ (_06070_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or _50773_ (_06071_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and _50774_ (_06072_, _06071_, _06070_);
  and _50775_ (_06073_, _06072_, _34796_);
  or _50776_ (_06074_, _06073_, _06069_);
  and _50777_ (_06075_, _06074_, _34772_);
  or _50778_ (_06076_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or _50779_ (_06077_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and _50780_ (_06078_, _06077_, _06076_);
  and _50781_ (_06079_, _06078_, _34581_);
  or _50782_ (_06080_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or _50783_ (_06081_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and _50784_ (_06082_, _06081_, _06080_);
  and _50785_ (_06083_, _06082_, _34796_);
  or _50786_ (_06084_, _06083_, _06079_);
  and _50787_ (_06085_, _06084_, _34790_);
  or _50788_ (_06086_, _06085_, _06075_);
  and _50789_ (_06087_, _06086_, _34719_);
  or _50790_ (_06088_, _06087_, _06065_);
  and _50791_ (_06089_, _06088_, _34700_);
  or _50792_ (_06090_, _06089_, _06043_);
  and _50793_ (_06091_, _06090_, _34638_);
  or _50794_ (_06092_, _06091_, _05997_);
  or _50795_ (_06093_, _06092_, _34985_);
  or _50796_ (_06094_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or _50797_ (_06095_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and _50798_ (_06096_, _06095_, _06094_);
  and _50799_ (_06097_, _06096_, _34581_);
  or _50800_ (_06098_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or _50801_ (_06099_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and _50802_ (_06100_, _06099_, _06098_);
  and _50803_ (_06101_, _06100_, _34796_);
  or _50804_ (_06102_, _06101_, _06097_);
  and _50805_ (_06103_, _06102_, _34790_);
  or _50806_ (_06104_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or _50807_ (_06105_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and _50808_ (_06106_, _06105_, _06104_);
  and _50809_ (_06107_, _06106_, _34581_);
  or _50810_ (_06108_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or _50811_ (_06109_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and _50812_ (_06110_, _06109_, _06108_);
  and _50813_ (_06111_, _06110_, _34796_);
  or _50814_ (_06112_, _06111_, _06107_);
  and _50815_ (_06113_, _06112_, _34772_);
  or _50816_ (_06114_, _06113_, _06103_);
  and _50817_ (_06115_, _06114_, _34719_);
  and _50818_ (_06116_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and _50819_ (_06117_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or _50820_ (_06118_, _06117_, _06116_);
  and _50821_ (_06119_, _06118_, _34581_);
  and _50822_ (_06120_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and _50823_ (_06121_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or _50824_ (_06122_, _06121_, _06120_);
  and _50825_ (_06123_, _06122_, _34796_);
  or _50826_ (_06124_, _06123_, _06119_);
  and _50827_ (_06125_, _06124_, _34790_);
  and _50828_ (_06126_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and _50829_ (_06127_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or _50830_ (_06128_, _06127_, _06126_);
  and _50831_ (_06129_, _06128_, _34581_);
  and _50832_ (_06130_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  and _50833_ (_06131_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or _50834_ (_06132_, _06131_, _06130_);
  and _50835_ (_06133_, _06132_, _34796_);
  or _50836_ (_06134_, _06133_, _06129_);
  and _50837_ (_06135_, _06134_, _34772_);
  or _50838_ (_06136_, _06135_, _06125_);
  and _50839_ (_06137_, _06136_, _34803_);
  or _50840_ (_06138_, _06137_, _06115_);
  and _50841_ (_06139_, _06138_, _34700_);
  or _50842_ (_06140_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or _50843_ (_06141_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and _50844_ (_06142_, _06141_, _34796_);
  and _50845_ (_06143_, _06142_, _06140_);
  or _50846_ (_06144_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or _50847_ (_06145_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and _50848_ (_06146_, _06145_, _34581_);
  and _50849_ (_06147_, _06146_, _06144_);
  or _50850_ (_06148_, _06147_, _06143_);
  and _50851_ (_06149_, _06148_, _34790_);
  or _50852_ (_06150_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or _50853_ (_06151_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and _50854_ (_06152_, _06151_, _34796_);
  and _50855_ (_06153_, _06152_, _06150_);
  or _50856_ (_06154_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or _50857_ (_06155_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and _50858_ (_06156_, _06155_, _34581_);
  and _50859_ (_06157_, _06156_, _06154_);
  or _50860_ (_06158_, _06157_, _06153_);
  and _50861_ (_06159_, _06158_, _34772_);
  or _50862_ (_06160_, _06159_, _06149_);
  and _50863_ (_06161_, _06160_, _34719_);
  and _50864_ (_06162_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and _50865_ (_06163_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or _50866_ (_06164_, _06163_, _06162_);
  and _50867_ (_06165_, _06164_, _34581_);
  and _50868_ (_06166_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and _50869_ (_06167_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or _50870_ (_06168_, _06167_, _06166_);
  and _50871_ (_06169_, _06168_, _34796_);
  or _50872_ (_06170_, _06169_, _06165_);
  and _50873_ (_06171_, _06170_, _34790_);
  and _50874_ (_06172_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and _50875_ (_06173_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or _50876_ (_06174_, _06173_, _06172_);
  and _50877_ (_06175_, _06174_, _34581_);
  and _50878_ (_06176_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and _50879_ (_06177_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or _50880_ (_06178_, _06177_, _06176_);
  and _50881_ (_06179_, _06178_, _34796_);
  or _50882_ (_06180_, _06179_, _06175_);
  and _50883_ (_06181_, _06180_, _34772_);
  or _50884_ (_06182_, _06181_, _06171_);
  and _50885_ (_06183_, _06182_, _34803_);
  or _50886_ (_06184_, _06183_, _06161_);
  and _50887_ (_06185_, _06184_, _34789_);
  or _50888_ (_06186_, _06185_, _06139_);
  and _50889_ (_06187_, _06186_, _34638_);
  and _50890_ (_06188_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and _50891_ (_06189_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or _50892_ (_06190_, _06189_, _06188_);
  and _50893_ (_06191_, _06190_, _34581_);
  and _50894_ (_06192_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  and _50895_ (_06193_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or _50896_ (_06194_, _06193_, _06192_);
  and _50897_ (_06195_, _06194_, _34796_);
  or _50898_ (_06196_, _06195_, _06191_);
  or _50899_ (_06197_, _06196_, _34790_);
  and _50900_ (_06198_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and _50901_ (_06199_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or _50902_ (_06200_, _06199_, _06198_);
  and _50903_ (_06201_, _06200_, _34581_);
  and _50904_ (_06202_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  and _50905_ (_06203_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or _50906_ (_06204_, _06203_, _06202_);
  and _50907_ (_06205_, _06204_, _34796_);
  or _50908_ (_06206_, _06205_, _06201_);
  or _50909_ (_06207_, _06206_, _34772_);
  and _50910_ (_06208_, _06207_, _34803_);
  and _50911_ (_06209_, _06208_, _06197_);
  or _50912_ (_06210_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or _50913_ (_06211_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  and _50914_ (_06212_, _06211_, _34796_);
  and _50915_ (_06213_, _06212_, _06210_);
  or _50916_ (_06214_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or _50917_ (_06215_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and _50918_ (_06216_, _06215_, _34581_);
  and _50919_ (_06217_, _06216_, _06214_);
  or _50920_ (_06218_, _06217_, _06213_);
  or _50921_ (_06219_, _06218_, _34790_);
  or _50922_ (_06220_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or _50923_ (_06221_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and _50924_ (_06222_, _06221_, _34796_);
  and _50925_ (_06223_, _06222_, _06220_);
  or _50926_ (_06224_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or _50927_ (_06225_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and _50928_ (_06226_, _06225_, _34581_);
  and _50929_ (_06227_, _06226_, _06224_);
  or _50930_ (_06228_, _06227_, _06223_);
  or _50931_ (_06229_, _06228_, _34772_);
  and _50932_ (_06230_, _06229_, _34719_);
  and _50933_ (_06231_, _06230_, _06219_);
  or _50934_ (_06232_, _06231_, _06209_);
  and _50935_ (_06233_, _06232_, _34789_);
  and _50936_ (_06234_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and _50937_ (_06235_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or _50938_ (_06236_, _06235_, _06234_);
  and _50939_ (_06237_, _06236_, _34581_);
  and _50940_ (_06238_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  and _50941_ (_06239_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or _50942_ (_06240_, _06239_, _06238_);
  and _50943_ (_06241_, _06240_, _34796_);
  or _50944_ (_06242_, _06241_, _06237_);
  or _50945_ (_06243_, _06242_, _34790_);
  and _50946_ (_06244_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and _50947_ (_06245_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or _50948_ (_06246_, _06245_, _06244_);
  and _50949_ (_06247_, _06246_, _34581_);
  and _50950_ (_06248_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and _50951_ (_06249_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or _50952_ (_06250_, _06249_, _06248_);
  and _50953_ (_06251_, _06250_, _34796_);
  or _50954_ (_06252_, _06251_, _06247_);
  or _50955_ (_06253_, _06252_, _34772_);
  and _50956_ (_06254_, _06253_, _34803_);
  and _50957_ (_06255_, _06254_, _06243_);
  or _50958_ (_06256_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or _50959_ (_06257_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  and _50960_ (_06258_, _06257_, _06256_);
  and _50961_ (_06259_, _06258_, _34581_);
  or _50962_ (_06260_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or _50963_ (_06261_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and _50964_ (_06262_, _06261_, _06260_);
  and _50965_ (_06263_, _06262_, _34796_);
  or _50966_ (_06264_, _06263_, _06259_);
  or _50967_ (_06265_, _06264_, _34790_);
  or _50968_ (_06266_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or _50969_ (_06267_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and _50970_ (_06268_, _06267_, _06266_);
  and _50971_ (_06269_, _06268_, _34581_);
  or _50972_ (_06270_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or _50973_ (_06271_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  and _50974_ (_06272_, _06271_, _06270_);
  and _50975_ (_06273_, _06272_, _34796_);
  or _50976_ (_06274_, _06273_, _06269_);
  or _50977_ (_06275_, _06274_, _34772_);
  and _50978_ (_06276_, _06275_, _34719_);
  and _50979_ (_06277_, _06276_, _06265_);
  or _50980_ (_06278_, _06277_, _06255_);
  and _50981_ (_06279_, _06278_, _34700_);
  or _50982_ (_06280_, _06279_, _06233_);
  and _50983_ (_06281_, _06280_, _34840_);
  or _50984_ (_06282_, _06281_, _06187_);
  or _50985_ (_06283_, _06282_, _34692_);
  and _50986_ (_06284_, _06283_, _35178_);
  and _50987_ (_06285_, _06284_, _06093_);
  or _50988_ (_06286_, _06285_, _05903_);
  or _50989_ (_06287_, _06286_, _34788_);
  or _50990_ (_06288_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and _50991_ (_06289_, _06288_, _38997_);
  and _50992_ (_38984_[0], _06289_, _06287_);
  and _50993_ (_06290_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and _50994_ (_06291_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or _50995_ (_06292_, _06291_, _06290_);
  and _50996_ (_06293_, _06292_, _34796_);
  and _50997_ (_06294_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and _50998_ (_06295_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or _50999_ (_06296_, _06295_, _06294_);
  and _51000_ (_06297_, _06296_, _34581_);
  or _51001_ (_06298_, _06297_, _06293_);
  or _51002_ (_06299_, _06298_, _34790_);
  and _51003_ (_06300_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and _51004_ (_06301_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or _51005_ (_06302_, _06301_, _06300_);
  and _51006_ (_06303_, _06302_, _34796_);
  and _51007_ (_06304_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  and _51008_ (_06305_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or _51009_ (_06306_, _06305_, _06304_);
  and _51010_ (_06307_, _06306_, _34581_);
  or _51011_ (_06308_, _06307_, _06303_);
  or _51012_ (_06309_, _06308_, _34772_);
  and _51013_ (_06310_, _06309_, _34803_);
  and _51014_ (_06311_, _06310_, _06299_);
  or _51015_ (_06312_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or _51016_ (_06313_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and _51017_ (_06314_, _06313_, _34581_);
  and _51018_ (_06315_, _06314_, _06312_);
  or _51019_ (_06316_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or _51020_ (_06317_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  and _51021_ (_06318_, _06317_, _34796_);
  and _51022_ (_06319_, _06318_, _06316_);
  or _51023_ (_06320_, _06319_, _06315_);
  or _51024_ (_06321_, _06320_, _34790_);
  or _51025_ (_06322_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or _51026_ (_06323_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and _51027_ (_06324_, _06323_, _34581_);
  and _51028_ (_06325_, _06324_, _06322_);
  or _51029_ (_06326_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or _51030_ (_06327_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  and _51031_ (_06328_, _06327_, _34796_);
  and _51032_ (_06329_, _06328_, _06326_);
  or _51033_ (_06330_, _06329_, _06325_);
  or _51034_ (_06331_, _06330_, _34772_);
  and _51035_ (_06332_, _06331_, _34719_);
  and _51036_ (_06333_, _06332_, _06321_);
  or _51037_ (_06334_, _06333_, _06311_);
  or _51038_ (_06335_, _06334_, _34700_);
  and _51039_ (_06336_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and _51040_ (_06337_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or _51041_ (_06338_, _06337_, _34581_);
  or _51042_ (_06339_, _06338_, _06336_);
  and _51043_ (_06340_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and _51044_ (_06341_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or _51045_ (_06342_, _06341_, _34796_);
  or _51046_ (_06343_, _06342_, _06340_);
  and _51047_ (_06344_, _06343_, _06339_);
  or _51048_ (_06345_, _06344_, _34790_);
  and _51049_ (_06346_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  and _51050_ (_06347_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or _51051_ (_06348_, _06347_, _34581_);
  or _51052_ (_06349_, _06348_, _06346_);
  and _51053_ (_06350_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and _51054_ (_06351_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or _51055_ (_06352_, _06351_, _34796_);
  or _51056_ (_06353_, _06352_, _06350_);
  and _51057_ (_06354_, _06353_, _06349_);
  or _51058_ (_06355_, _06354_, _34772_);
  and _51059_ (_06356_, _06355_, _34803_);
  and _51060_ (_06357_, _06356_, _06345_);
  or _51061_ (_06358_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or _51062_ (_06359_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and _51063_ (_06360_, _06359_, _06358_);
  or _51064_ (_06361_, _06360_, _34796_);
  or _51065_ (_06362_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or _51066_ (_06363_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and _51067_ (_06364_, _06363_, _06362_);
  or _51068_ (_06365_, _06364_, _34581_);
  and _51069_ (_06366_, _06365_, _06361_);
  or _51070_ (_06367_, _06366_, _34790_);
  or _51071_ (_06368_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or _51072_ (_06369_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  and _51073_ (_06370_, _06369_, _06368_);
  or _51074_ (_06371_, _06370_, _34796_);
  or _51075_ (_06372_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or _51076_ (_06373_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and _51077_ (_06374_, _06373_, _06372_);
  or _51078_ (_06375_, _06374_, _34581_);
  and _51079_ (_06376_, _06375_, _06371_);
  or _51080_ (_06377_, _06376_, _34772_);
  and _51081_ (_06378_, _06377_, _34719_);
  and _51082_ (_06379_, _06378_, _06367_);
  or _51083_ (_06380_, _06379_, _06357_);
  or _51084_ (_06381_, _06380_, _34789_);
  and _51085_ (_06382_, _06381_, _34840_);
  and _51086_ (_06383_, _06382_, _06335_);
  and _51087_ (_06384_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and _51088_ (_06385_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or _51089_ (_06386_, _06385_, _06384_);
  and _51090_ (_06387_, _06386_, _34581_);
  and _51091_ (_06388_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and _51092_ (_06389_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _51093_ (_06390_, _06389_, _06388_);
  and _51094_ (_06391_, _06390_, _34796_);
  or _51095_ (_06392_, _06391_, _06387_);
  and _51096_ (_06393_, _06392_, _34772_);
  and _51097_ (_06394_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and _51098_ (_06395_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or _51099_ (_06396_, _06395_, _06394_);
  and _51100_ (_06397_, _06396_, _34581_);
  and _51101_ (_06398_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and _51102_ (_06399_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _51103_ (_06400_, _06399_, _06398_);
  and _51104_ (_06401_, _06400_, _34796_);
  or _51105_ (_06402_, _06401_, _06397_);
  and _51106_ (_06403_, _06402_, _34790_);
  or _51107_ (_06404_, _06403_, _06393_);
  and _51108_ (_06405_, _06404_, _34803_);
  or _51109_ (_06406_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or _51110_ (_06407_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _51111_ (_06408_, _06407_, _06406_);
  and _51112_ (_06409_, _06408_, _34581_);
  or _51113_ (_06410_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or _51114_ (_06411_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and _51115_ (_06412_, _06411_, _06410_);
  and _51116_ (_06413_, _06412_, _34796_);
  or _51117_ (_06414_, _06413_, _06409_);
  and _51118_ (_06415_, _06414_, _34772_);
  or _51119_ (_06416_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or _51120_ (_06417_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _51121_ (_06418_, _06417_, _06416_);
  and _51122_ (_06419_, _06418_, _34581_);
  or _51123_ (_06420_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or _51124_ (_06421_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and _51125_ (_06422_, _06421_, _06420_);
  and _51126_ (_06423_, _06422_, _34796_);
  or _51127_ (_06424_, _06423_, _06419_);
  and _51128_ (_06425_, _06424_, _34790_);
  or _51129_ (_06426_, _06425_, _06415_);
  and _51130_ (_06427_, _06426_, _34719_);
  or _51131_ (_06428_, _06427_, _06405_);
  and _51132_ (_06429_, _06428_, _34789_);
  and _51133_ (_06430_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  and _51134_ (_06431_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or _51135_ (_06432_, _06431_, _06430_);
  and _51136_ (_06433_, _06432_, _34581_);
  and _51137_ (_06434_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and _51138_ (_06435_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or _51139_ (_06436_, _06435_, _06434_);
  and _51140_ (_06437_, _06436_, _34796_);
  or _51141_ (_06438_, _06437_, _06433_);
  and _51142_ (_06439_, _06438_, _34772_);
  and _51143_ (_06440_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and _51144_ (_06441_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or _51145_ (_06442_, _06441_, _06440_);
  and _51146_ (_06443_, _06442_, _34581_);
  and _51147_ (_06444_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and _51148_ (_06445_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or _51149_ (_06446_, _06445_, _06444_);
  and _51150_ (_06447_, _06446_, _34796_);
  or _51151_ (_06448_, _06447_, _06443_);
  and _51152_ (_06449_, _06448_, _34790_);
  or _51153_ (_06450_, _06449_, _06439_);
  and _51154_ (_06451_, _06450_, _34803_);
  or _51155_ (_06452_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or _51156_ (_06453_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  and _51157_ (_06454_, _06453_, _06452_);
  and _51158_ (_06455_, _06454_, _34581_);
  or _51159_ (_06456_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or _51160_ (_06457_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and _51161_ (_06458_, _06457_, _06456_);
  and _51162_ (_06459_, _06458_, _34796_);
  or _51163_ (_06460_, _06459_, _06455_);
  and _51164_ (_06461_, _06460_, _34772_);
  or _51165_ (_06462_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or _51166_ (_06463_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and _51167_ (_06464_, _06463_, _06462_);
  and _51168_ (_06465_, _06464_, _34581_);
  or _51169_ (_06466_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or _51170_ (_06467_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and _51171_ (_06468_, _06467_, _06466_);
  and _51172_ (_06469_, _06468_, _34796_);
  or _51173_ (_06470_, _06469_, _06465_);
  and _51174_ (_06471_, _06470_, _34790_);
  or _51175_ (_06472_, _06471_, _06461_);
  and _51176_ (_06473_, _06472_, _34719_);
  or _51177_ (_06474_, _06473_, _06451_);
  and _51178_ (_06475_, _06474_, _34700_);
  or _51179_ (_06476_, _06475_, _06429_);
  and _51180_ (_06477_, _06476_, _34638_);
  or _51181_ (_06478_, _06477_, _06383_);
  or _51182_ (_06479_, _06478_, _34692_);
  and _51183_ (_06480_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  and _51184_ (_06481_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or _51185_ (_06482_, _06481_, _06480_);
  and _51186_ (_06483_, _06482_, _34581_);
  and _51187_ (_06484_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and _51188_ (_06485_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or _51189_ (_06486_, _06485_, _06484_);
  and _51190_ (_06487_, _06486_, _34796_);
  or _51191_ (_06488_, _06487_, _06483_);
  or _51192_ (_06489_, _06488_, _34790_);
  and _51193_ (_06490_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  and _51194_ (_06491_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or _51195_ (_06492_, _06491_, _06490_);
  and _51196_ (_06493_, _06492_, _34581_);
  and _51197_ (_06494_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and _51198_ (_06495_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or _51199_ (_06496_, _06495_, _06494_);
  and _51200_ (_06497_, _06496_, _34796_);
  or _51201_ (_06498_, _06497_, _06493_);
  or _51202_ (_06499_, _06498_, _34772_);
  and _51203_ (_06500_, _06499_, _34803_);
  and _51204_ (_06501_, _06500_, _06489_);
  or _51205_ (_06502_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or _51206_ (_06503_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and _51207_ (_06504_, _06503_, _34796_);
  and _51208_ (_06505_, _06504_, _06502_);
  or _51209_ (_06506_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or _51210_ (_06507_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and _51211_ (_06508_, _06507_, _34581_);
  and _51212_ (_06509_, _06508_, _06506_);
  or _51213_ (_06510_, _06509_, _06505_);
  or _51214_ (_06511_, _06510_, _34790_);
  or _51215_ (_06512_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or _51216_ (_06513_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and _51217_ (_06514_, _06513_, _34796_);
  and _51218_ (_06515_, _06514_, _06512_);
  or _51219_ (_06516_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or _51220_ (_06517_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  and _51221_ (_06518_, _06517_, _34581_);
  and _51222_ (_06519_, _06518_, _06516_);
  or _51223_ (_06520_, _06519_, _06515_);
  or _51224_ (_06521_, _06520_, _34772_);
  and _51225_ (_06522_, _06521_, _34719_);
  and _51226_ (_06523_, _06522_, _06511_);
  or _51227_ (_06524_, _06523_, _06501_);
  and _51228_ (_06525_, _06524_, _34789_);
  and _51229_ (_06526_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and _51230_ (_06527_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or _51231_ (_06528_, _06527_, _06526_);
  and _51232_ (_06529_, _06528_, _34581_);
  and _51233_ (_06530_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and _51234_ (_06531_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or _51235_ (_06532_, _06531_, _06530_);
  and _51236_ (_06533_, _06532_, _34796_);
  or _51237_ (_06534_, _06533_, _06529_);
  or _51238_ (_06535_, _06534_, _34790_);
  and _51239_ (_06536_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and _51240_ (_06537_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or _51241_ (_06538_, _06537_, _06536_);
  and _51242_ (_06539_, _06538_, _34581_);
  and _51243_ (_06540_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and _51244_ (_06541_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or _51245_ (_06542_, _06541_, _06540_);
  and _51246_ (_06543_, _06542_, _34796_);
  or _51247_ (_06544_, _06543_, _06539_);
  or _51248_ (_06545_, _06544_, _34772_);
  and _51249_ (_06546_, _06545_, _34803_);
  and _51250_ (_06547_, _06546_, _06535_);
  or _51251_ (_06548_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or _51252_ (_06549_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and _51253_ (_06550_, _06549_, _06548_);
  and _51254_ (_06551_, _06550_, _34581_);
  or _51255_ (_06552_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or _51256_ (_06553_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and _51257_ (_06554_, _06553_, _06552_);
  and _51258_ (_06555_, _06554_, _34796_);
  or _51259_ (_06556_, _06555_, _06551_);
  or _51260_ (_06557_, _06556_, _34790_);
  or _51261_ (_06558_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or _51262_ (_06559_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and _51263_ (_06560_, _06559_, _06558_);
  and _51264_ (_06561_, _06560_, _34581_);
  or _51265_ (_06562_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or _51266_ (_06563_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and _51267_ (_06564_, _06563_, _06562_);
  and _51268_ (_06565_, _06564_, _34796_);
  or _51269_ (_06566_, _06565_, _06561_);
  or _51270_ (_06567_, _06566_, _34772_);
  and _51271_ (_06568_, _06567_, _34719_);
  and _51272_ (_06569_, _06568_, _06557_);
  or _51273_ (_06570_, _06569_, _06547_);
  and _51274_ (_06571_, _06570_, _34700_);
  or _51275_ (_06572_, _06571_, _06525_);
  and _51276_ (_06573_, _06572_, _34840_);
  or _51277_ (_06574_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or _51278_ (_06575_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and _51279_ (_06576_, _06575_, _06574_);
  and _51280_ (_06577_, _06576_, _34581_);
  or _51281_ (_06578_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or _51282_ (_06579_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  and _51283_ (_06580_, _06579_, _06578_);
  and _51284_ (_06581_, _06580_, _34796_);
  or _51285_ (_06582_, _06581_, _06577_);
  and _51286_ (_06583_, _06582_, _34790_);
  or _51287_ (_06584_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or _51288_ (_06585_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and _51289_ (_06586_, _06585_, _06584_);
  and _51290_ (_06587_, _06586_, _34581_);
  or _51291_ (_06588_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or _51292_ (_06589_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  and _51293_ (_06590_, _06589_, _06588_);
  and _51294_ (_06591_, _06590_, _34796_);
  or _51295_ (_06592_, _06591_, _06587_);
  and _51296_ (_06593_, _06592_, _34772_);
  or _51297_ (_06594_, _06593_, _06583_);
  and _51298_ (_06595_, _06594_, _34719_);
  and _51299_ (_06596_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and _51300_ (_06597_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or _51301_ (_06598_, _06597_, _06596_);
  and _51302_ (_06599_, _06598_, _34581_);
  and _51303_ (_06600_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  and _51304_ (_06601_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or _51305_ (_06602_, _06601_, _06600_);
  and _51306_ (_06603_, _06602_, _34796_);
  or _51307_ (_06604_, _06603_, _06599_);
  and _51308_ (_06605_, _06604_, _34790_);
  and _51309_ (_06606_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and _51310_ (_06607_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or _51311_ (_06608_, _06607_, _06606_);
  and _51312_ (_06609_, _06608_, _34581_);
  and _51313_ (_06610_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  and _51314_ (_06611_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or _51315_ (_06612_, _06611_, _06610_);
  and _51316_ (_06613_, _06612_, _34796_);
  or _51317_ (_06614_, _06613_, _06609_);
  and _51318_ (_06615_, _06614_, _34772_);
  or _51319_ (_06616_, _06615_, _06605_);
  and _51320_ (_06617_, _06616_, _34803_);
  or _51321_ (_06618_, _06617_, _06595_);
  and _51322_ (_06619_, _06618_, _34700_);
  or _51323_ (_06620_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or _51324_ (_06621_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  and _51325_ (_06622_, _06621_, _34796_);
  and _51326_ (_06623_, _06622_, _06620_);
  or _51327_ (_06624_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or _51328_ (_06625_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and _51329_ (_06626_, _06625_, _34581_);
  and _51330_ (_06627_, _06626_, _06624_);
  or _51331_ (_06628_, _06627_, _06623_);
  and _51332_ (_06629_, _06628_, _34790_);
  or _51333_ (_06630_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or _51334_ (_06631_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  and _51335_ (_06632_, _06631_, _34796_);
  and _51336_ (_06633_, _06632_, _06630_);
  or _51337_ (_06634_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or _51338_ (_06635_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  and _51339_ (_06636_, _06635_, _34581_);
  and _51340_ (_06637_, _06636_, _06634_);
  or _51341_ (_06638_, _06637_, _06633_);
  and _51342_ (_06639_, _06638_, _34772_);
  or _51343_ (_06640_, _06639_, _06629_);
  and _51344_ (_06641_, _06640_, _34719_);
  and _51345_ (_06642_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  and _51346_ (_06643_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or _51347_ (_06644_, _06643_, _06642_);
  and _51348_ (_06645_, _06644_, _34581_);
  and _51349_ (_06646_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  and _51350_ (_06647_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or _51351_ (_06648_, _06647_, _06646_);
  and _51352_ (_06649_, _06648_, _34796_);
  or _51353_ (_06650_, _06649_, _06645_);
  and _51354_ (_06651_, _06650_, _34790_);
  and _51355_ (_06652_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and _51356_ (_06653_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or _51357_ (_06654_, _06653_, _06652_);
  and _51358_ (_06655_, _06654_, _34581_);
  and _51359_ (_06656_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  and _51360_ (_06657_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or _51361_ (_06658_, _06657_, _06656_);
  and _51362_ (_06659_, _06658_, _34796_);
  or _51363_ (_06660_, _06659_, _06655_);
  and _51364_ (_06661_, _06660_, _34772_);
  or _51365_ (_06662_, _06661_, _06651_);
  and _51366_ (_06663_, _06662_, _34803_);
  or _51367_ (_06664_, _06663_, _06641_);
  and _51368_ (_06665_, _06664_, _34789_);
  or _51369_ (_06666_, _06665_, _06619_);
  and _51370_ (_06667_, _06666_, _34638_);
  or _51371_ (_06668_, _06667_, _06573_);
  or _51372_ (_06669_, _06668_, _34985_);
  and _51373_ (_06670_, _06669_, _06479_);
  or _51374_ (_06671_, _06670_, _34346_);
  and _51375_ (_06672_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and _51376_ (_06673_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or _51377_ (_06674_, _06673_, _06672_);
  and _51378_ (_06675_, _06674_, _34796_);
  and _51379_ (_06676_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and _51380_ (_06677_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or _51381_ (_06678_, _06677_, _06676_);
  and _51382_ (_06679_, _06678_, _34581_);
  or _51383_ (_06680_, _06679_, _06675_);
  or _51384_ (_06681_, _06680_, _34790_);
  and _51385_ (_06682_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and _51386_ (_06683_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or _51387_ (_06684_, _06683_, _06682_);
  and _51388_ (_06685_, _06684_, _34796_);
  and _51389_ (_06686_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and _51390_ (_06687_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or _51391_ (_06688_, _06687_, _06686_);
  and _51392_ (_06689_, _06688_, _34581_);
  or _51393_ (_06690_, _06689_, _06685_);
  or _51394_ (_06691_, _06690_, _34772_);
  and _51395_ (_06692_, _06691_, _34803_);
  and _51396_ (_06693_, _06692_, _06681_);
  or _51397_ (_06694_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or _51398_ (_06695_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and _51399_ (_06696_, _06695_, _34581_);
  and _51400_ (_06697_, _06696_, _06694_);
  or _51401_ (_06698_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or _51402_ (_06699_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and _51403_ (_06700_, _06699_, _34796_);
  and _51404_ (_06701_, _06700_, _06698_);
  or _51405_ (_06702_, _06701_, _06697_);
  or _51406_ (_06703_, _06702_, _34790_);
  or _51407_ (_06704_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or _51408_ (_06705_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and _51409_ (_06706_, _06705_, _34581_);
  and _51410_ (_06707_, _06706_, _06704_);
  or _51411_ (_06708_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or _51412_ (_06709_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and _51413_ (_06710_, _06709_, _34796_);
  and _51414_ (_06711_, _06710_, _06708_);
  or _51415_ (_06712_, _06711_, _06707_);
  or _51416_ (_06713_, _06712_, _34772_);
  and _51417_ (_06714_, _06713_, _34719_);
  and _51418_ (_06715_, _06714_, _06703_);
  or _51419_ (_06716_, _06715_, _06693_);
  and _51420_ (_06717_, _06716_, _34789_);
  and _51421_ (_06718_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and _51422_ (_06719_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or _51423_ (_06720_, _06719_, _34581_);
  or _51424_ (_06721_, _06720_, _06718_);
  and _51425_ (_06722_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and _51426_ (_06723_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or _51427_ (_06724_, _06723_, _34796_);
  or _51428_ (_06725_, _06724_, _06722_);
  and _51429_ (_06726_, _06725_, _06721_);
  or _51430_ (_06727_, _06726_, _34790_);
  and _51431_ (_06728_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and _51432_ (_06729_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or _51433_ (_06730_, _06729_, _34581_);
  or _51434_ (_06731_, _06730_, _06728_);
  and _51435_ (_06732_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and _51436_ (_06733_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or _51437_ (_06734_, _06733_, _34796_);
  or _51438_ (_06735_, _06734_, _06732_);
  and _51439_ (_06736_, _06735_, _06731_);
  or _51440_ (_06737_, _06736_, _34772_);
  and _51441_ (_06738_, _06737_, _34803_);
  and _51442_ (_06739_, _06738_, _06727_);
  or _51443_ (_06740_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or _51444_ (_06741_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and _51445_ (_06742_, _06741_, _06740_);
  or _51446_ (_06743_, _06742_, _34796_);
  or _51447_ (_06744_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or _51448_ (_06745_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and _51449_ (_06746_, _06745_, _06744_);
  or _51450_ (_06747_, _06746_, _34581_);
  and _51451_ (_06748_, _06747_, _06743_);
  or _51452_ (_06749_, _06748_, _34790_);
  or _51453_ (_06750_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or _51454_ (_06751_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and _51455_ (_06752_, _06751_, _06750_);
  or _51456_ (_06753_, _06752_, _34796_);
  or _51457_ (_06754_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or _51458_ (_06755_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and _51459_ (_06756_, _06755_, _06754_);
  or _51460_ (_06757_, _06756_, _34581_);
  and _51461_ (_06758_, _06757_, _06753_);
  or _51462_ (_06759_, _06758_, _34772_);
  and _51463_ (_06760_, _06759_, _34719_);
  and _51464_ (_06761_, _06760_, _06749_);
  or _51465_ (_06762_, _06761_, _06739_);
  and _51466_ (_06763_, _06762_, _34700_);
  or _51467_ (_06764_, _06763_, _06717_);
  and _51468_ (_06765_, _06764_, _34840_);
  and _51469_ (_06766_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  and _51470_ (_06767_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  or _51471_ (_06768_, _06767_, _06766_);
  and _51472_ (_06769_, _06768_, _34581_);
  and _51473_ (_06770_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  and _51474_ (_06771_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  or _51475_ (_06772_, _06771_, _06770_);
  and _51476_ (_06773_, _06772_, _34796_);
  or _51477_ (_06774_, _06773_, _06769_);
  and _51478_ (_06775_, _06774_, _34772_);
  and _51479_ (_06776_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  and _51480_ (_06777_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  or _51481_ (_06778_, _06777_, _06776_);
  and _51482_ (_06779_, _06778_, _34581_);
  and _51483_ (_06780_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  and _51484_ (_06781_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  or _51485_ (_06782_, _06781_, _06780_);
  and _51486_ (_06783_, _06782_, _34796_);
  or _51487_ (_06784_, _06783_, _06779_);
  and _51488_ (_06785_, _06784_, _34790_);
  or _51489_ (_06786_, _06785_, _06775_);
  and _51490_ (_06787_, _06786_, _34803_);
  or _51491_ (_06788_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  or _51492_ (_06789_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  and _51493_ (_06790_, _06789_, _06788_);
  and _51494_ (_06791_, _06790_, _34581_);
  or _51495_ (_06792_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  or _51496_ (_06793_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  and _51497_ (_06794_, _06793_, _06792_);
  and _51498_ (_06795_, _06794_, _34796_);
  or _51499_ (_06796_, _06795_, _06791_);
  and _51500_ (_06797_, _06796_, _34772_);
  or _51501_ (_06798_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  or _51502_ (_06799_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  and _51503_ (_06800_, _06799_, _06798_);
  and _51504_ (_06801_, _06800_, _34581_);
  or _51505_ (_06802_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  or _51506_ (_06803_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  and _51507_ (_06804_, _06803_, _06802_);
  and _51508_ (_06805_, _06804_, _34796_);
  or _51509_ (_06806_, _06805_, _06801_);
  and _51510_ (_06807_, _06806_, _34790_);
  or _51511_ (_06808_, _06807_, _06797_);
  and _51512_ (_06809_, _06808_, _34719_);
  or _51513_ (_06810_, _06809_, _06787_);
  and _51514_ (_06811_, _06810_, _34789_);
  and _51515_ (_06812_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and _51516_ (_06813_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or _51517_ (_06814_, _06813_, _06812_);
  and _51518_ (_06815_, _06814_, _34581_);
  and _51519_ (_06816_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and _51520_ (_06817_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or _51521_ (_06818_, _06817_, _06816_);
  and _51522_ (_06819_, _06818_, _34796_);
  or _51523_ (_06820_, _06819_, _06815_);
  and _51524_ (_06821_, _06820_, _34772_);
  and _51525_ (_06822_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and _51526_ (_06823_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or _51527_ (_06824_, _06823_, _06822_);
  and _51528_ (_06825_, _06824_, _34581_);
  and _51529_ (_06826_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and _51530_ (_06827_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or _51531_ (_06828_, _06827_, _06826_);
  and _51532_ (_06829_, _06828_, _34796_);
  or _51533_ (_06830_, _06829_, _06825_);
  and _51534_ (_06831_, _06830_, _34790_);
  or _51535_ (_06832_, _06831_, _06821_);
  and _51536_ (_06833_, _06832_, _34803_);
  or _51537_ (_06834_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or _51538_ (_06835_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and _51539_ (_06836_, _06835_, _06834_);
  and _51540_ (_06837_, _06836_, _34581_);
  or _51541_ (_06838_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or _51542_ (_06839_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and _51543_ (_06840_, _06839_, _06838_);
  and _51544_ (_06841_, _06840_, _34796_);
  or _51545_ (_06842_, _06841_, _06837_);
  and _51546_ (_06843_, _06842_, _34772_);
  or _51547_ (_06844_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or _51548_ (_06845_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and _51549_ (_06846_, _06845_, _06844_);
  and _51550_ (_06847_, _06846_, _34581_);
  or _51551_ (_06848_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or _51552_ (_06849_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and _51553_ (_06850_, _06849_, _06848_);
  and _51554_ (_06851_, _06850_, _34796_);
  or _51555_ (_06852_, _06851_, _06847_);
  and _51556_ (_06853_, _06852_, _34790_);
  or _51557_ (_06854_, _06853_, _06843_);
  and _51558_ (_06855_, _06854_, _34719_);
  or _51559_ (_06856_, _06855_, _06833_);
  and _51560_ (_06857_, _06856_, _34700_);
  or _51561_ (_06858_, _06857_, _06811_);
  and _51562_ (_06859_, _06858_, _34638_);
  or _51563_ (_06860_, _06859_, _06765_);
  or _51564_ (_06861_, _06860_, _34692_);
  and _51565_ (_06862_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and _51566_ (_06863_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or _51567_ (_06864_, _06863_, _06862_);
  and _51568_ (_06865_, _06864_, _34581_);
  and _51569_ (_06866_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and _51570_ (_06867_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or _51571_ (_06868_, _06867_, _06866_);
  and _51572_ (_06869_, _06868_, _34796_);
  or _51573_ (_06870_, _06869_, _06865_);
  or _51574_ (_06871_, _06870_, _34790_);
  and _51575_ (_06872_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and _51576_ (_06873_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or _51577_ (_06874_, _06873_, _06872_);
  and _51578_ (_06875_, _06874_, _34581_);
  and _51579_ (_06876_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and _51580_ (_06877_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or _51581_ (_06878_, _06877_, _06876_);
  and _51582_ (_06879_, _06878_, _34796_);
  or _51583_ (_06880_, _06879_, _06875_);
  or _51584_ (_06881_, _06880_, _34772_);
  and _51585_ (_06882_, _06881_, _34803_);
  and _51586_ (_06883_, _06882_, _06871_);
  or _51587_ (_06884_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or _51588_ (_06885_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and _51589_ (_06886_, _06885_, _34796_);
  and _51590_ (_06887_, _06886_, _06884_);
  or _51591_ (_06888_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or _51592_ (_06889_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and _51593_ (_06890_, _06889_, _34581_);
  and _51594_ (_06891_, _06890_, _06888_);
  or _51595_ (_06892_, _06891_, _06887_);
  or _51596_ (_06893_, _06892_, _34790_);
  or _51597_ (_06894_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or _51598_ (_06895_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and _51599_ (_06896_, _06895_, _34796_);
  and _51600_ (_06897_, _06896_, _06894_);
  or _51601_ (_06898_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or _51602_ (_06899_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and _51603_ (_06900_, _06899_, _34581_);
  and _51604_ (_06901_, _06900_, _06898_);
  or _51605_ (_06902_, _06901_, _06897_);
  or _51606_ (_06903_, _06902_, _34772_);
  and _51607_ (_06904_, _06903_, _34719_);
  and _51608_ (_06905_, _06904_, _06893_);
  or _51609_ (_06906_, _06905_, _06883_);
  and _51610_ (_06907_, _06906_, _34789_);
  and _51611_ (_06908_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and _51612_ (_06909_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or _51613_ (_06910_, _06909_, _06908_);
  and _51614_ (_06911_, _06910_, _34581_);
  and _51615_ (_06912_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and _51616_ (_06913_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or _51617_ (_06914_, _06913_, _06912_);
  and _51618_ (_06915_, _06914_, _34796_);
  or _51619_ (_06916_, _06915_, _06911_);
  or _51620_ (_06917_, _06916_, _34790_);
  and _51621_ (_06918_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and _51622_ (_06919_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or _51623_ (_06920_, _06919_, _06918_);
  and _51624_ (_06921_, _06920_, _34581_);
  and _51625_ (_06922_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and _51626_ (_06923_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or _51627_ (_06924_, _06923_, _06922_);
  and _51628_ (_06925_, _06924_, _34796_);
  or _51629_ (_06926_, _06925_, _06921_);
  or _51630_ (_06927_, _06926_, _34772_);
  and _51631_ (_06928_, _06927_, _34803_);
  and _51632_ (_06929_, _06928_, _06917_);
  or _51633_ (_06930_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or _51634_ (_06931_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and _51635_ (_06932_, _06931_, _06930_);
  and _51636_ (_06933_, _06932_, _34581_);
  or _51637_ (_06934_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or _51638_ (_06935_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and _51639_ (_06936_, _06935_, _06934_);
  and _51640_ (_06937_, _06936_, _34796_);
  or _51641_ (_06938_, _06937_, _06933_);
  or _51642_ (_06939_, _06938_, _34790_);
  or _51643_ (_06940_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or _51644_ (_06941_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and _51645_ (_06942_, _06941_, _06940_);
  and _51646_ (_06943_, _06942_, _34581_);
  or _51647_ (_06944_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or _51648_ (_06945_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and _51649_ (_06946_, _06945_, _06944_);
  and _51650_ (_06947_, _06946_, _34796_);
  or _51651_ (_06948_, _06947_, _06943_);
  or _51652_ (_06949_, _06948_, _34772_);
  and _51653_ (_06950_, _06949_, _34719_);
  and _51654_ (_06951_, _06950_, _06939_);
  or _51655_ (_06952_, _06951_, _06929_);
  and _51656_ (_06953_, _06952_, _34700_);
  or _51657_ (_06954_, _06953_, _06907_);
  and _51658_ (_06955_, _06954_, _34840_);
  or _51659_ (_06956_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or _51660_ (_06957_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and _51661_ (_06958_, _06957_, _06956_);
  and _51662_ (_06959_, _06958_, _34581_);
  or _51663_ (_06960_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or _51664_ (_06961_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and _51665_ (_06962_, _06961_, _06960_);
  and _51666_ (_06963_, _06962_, _34796_);
  or _51667_ (_06964_, _06963_, _06959_);
  and _51668_ (_06965_, _06964_, _34790_);
  or _51669_ (_06966_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or _51670_ (_06967_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and _51671_ (_06968_, _06967_, _06966_);
  and _51672_ (_06969_, _06968_, _34581_);
  or _51673_ (_06970_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or _51674_ (_06971_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and _51675_ (_06972_, _06971_, _06970_);
  and _51676_ (_06973_, _06972_, _34796_);
  or _51677_ (_06974_, _06973_, _06969_);
  and _51678_ (_06975_, _06974_, _34772_);
  or _51679_ (_06976_, _06975_, _06965_);
  and _51680_ (_06977_, _06976_, _34719_);
  and _51681_ (_06978_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and _51682_ (_06979_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or _51683_ (_06980_, _06979_, _06978_);
  and _51684_ (_06981_, _06980_, _34581_);
  and _51685_ (_06982_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and _51686_ (_06983_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or _51687_ (_06984_, _06983_, _06982_);
  and _51688_ (_06985_, _06984_, _34796_);
  or _51689_ (_06986_, _06985_, _06981_);
  and _51690_ (_06987_, _06986_, _34790_);
  and _51691_ (_06988_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and _51692_ (_06989_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or _51693_ (_06990_, _06989_, _06988_);
  and _51694_ (_06991_, _06990_, _34581_);
  and _51695_ (_06992_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and _51696_ (_06993_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or _51697_ (_06994_, _06993_, _06992_);
  and _51698_ (_06995_, _06994_, _34796_);
  or _51699_ (_06996_, _06995_, _06991_);
  and _51700_ (_06997_, _06996_, _34772_);
  or _51701_ (_06998_, _06997_, _06987_);
  and _51702_ (_06999_, _06998_, _34803_);
  or _51703_ (_07000_, _06999_, _06977_);
  and _51704_ (_07001_, _07000_, _34700_);
  or _51705_ (_07002_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or _51706_ (_07003_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and _51707_ (_07004_, _07003_, _34796_);
  and _51708_ (_07005_, _07004_, _07002_);
  or _51709_ (_07006_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or _51710_ (_07007_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and _51711_ (_07008_, _07007_, _34581_);
  and _51712_ (_07009_, _07008_, _07006_);
  or _51713_ (_07010_, _07009_, _07005_);
  and _51714_ (_07011_, _07010_, _34790_);
  or _51715_ (_07012_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or _51716_ (_07013_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and _51717_ (_07014_, _07013_, _34796_);
  and _51718_ (_07015_, _07014_, _07012_);
  or _51719_ (_07016_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or _51720_ (_07017_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and _51721_ (_07018_, _07017_, _34581_);
  and _51722_ (_07019_, _07018_, _07016_);
  or _51723_ (_07020_, _07019_, _07015_);
  and _51724_ (_07021_, _07020_, _34772_);
  or _51725_ (_07022_, _07021_, _07011_);
  and _51726_ (_07023_, _07022_, _34719_);
  and _51727_ (_07024_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and _51728_ (_07025_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or _51729_ (_07026_, _07025_, _07024_);
  and _51730_ (_07027_, _07026_, _34581_);
  and _51731_ (_07028_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and _51732_ (_07029_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or _51733_ (_07030_, _07029_, _07028_);
  and _51734_ (_07031_, _07030_, _34796_);
  or _51735_ (_07032_, _07031_, _07027_);
  and _51736_ (_07033_, _07032_, _34790_);
  and _51737_ (_07034_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and _51738_ (_07035_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or _51739_ (_07036_, _07035_, _07034_);
  and _51740_ (_07037_, _07036_, _34581_);
  and _51741_ (_07038_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and _51742_ (_07039_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or _51743_ (_07040_, _07039_, _07038_);
  and _51744_ (_07041_, _07040_, _34796_);
  or _51745_ (_07042_, _07041_, _07037_);
  and _51746_ (_07043_, _07042_, _34772_);
  or _51747_ (_07044_, _07043_, _07033_);
  and _51748_ (_07045_, _07044_, _34803_);
  or _51749_ (_07046_, _07045_, _07023_);
  and _51750_ (_07047_, _07046_, _34789_);
  or _51751_ (_07048_, _07047_, _07001_);
  and _51752_ (_07049_, _07048_, _34638_);
  or _51753_ (_07050_, _07049_, _06955_);
  or _51754_ (_07051_, _07050_, _34985_);
  and _51755_ (_07052_, _07051_, _06861_);
  or _51756_ (_07053_, _07052_, _35178_);
  and _51757_ (_07054_, _07053_, _06671_);
  or _51758_ (_07055_, _07054_, _34788_);
  or _51759_ (_07056_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and _51760_ (_07057_, _07056_, _38997_);
  and _51761_ (_38984_[1], _07057_, _07055_);
  and _51762_ (_07058_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and _51763_ (_07059_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or _51764_ (_07060_, _07059_, _07058_);
  and _51765_ (_07061_, _07060_, _34581_);
  and _51766_ (_07062_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and _51767_ (_07063_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or _51768_ (_07064_, _07063_, _07062_);
  and _51769_ (_07065_, _07064_, _34796_);
  or _51770_ (_07066_, _07065_, _07061_);
  or _51771_ (_07067_, _07066_, _34790_);
  and _51772_ (_07068_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and _51773_ (_07069_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or _51774_ (_07070_, _07069_, _07068_);
  and _51775_ (_07071_, _07070_, _34581_);
  and _51776_ (_07072_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and _51777_ (_07073_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or _51778_ (_07074_, _07073_, _07072_);
  and _51779_ (_07075_, _07074_, _34796_);
  or _51780_ (_07076_, _07075_, _07071_);
  or _51781_ (_07077_, _07076_, _34772_);
  and _51782_ (_07078_, _07077_, _34803_);
  and _51783_ (_07079_, _07078_, _07067_);
  or _51784_ (_07080_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or _51785_ (_07081_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and _51786_ (_07082_, _07081_, _07080_);
  and _51787_ (_07083_, _07082_, _34581_);
  or _51788_ (_07084_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or _51789_ (_07085_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and _51790_ (_07086_, _07085_, _07084_);
  and _51791_ (_07087_, _07086_, _34796_);
  or _51792_ (_07088_, _07087_, _07083_);
  or _51793_ (_07089_, _07088_, _34790_);
  or _51794_ (_07090_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or _51795_ (_07091_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and _51796_ (_07092_, _07091_, _07090_);
  and _51797_ (_07093_, _07092_, _34581_);
  or _51798_ (_07094_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or _51799_ (_07095_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and _51800_ (_07096_, _07095_, _07094_);
  and _51801_ (_07097_, _07096_, _34796_);
  or _51802_ (_07098_, _07097_, _07093_);
  or _51803_ (_07099_, _07098_, _34772_);
  and _51804_ (_07100_, _07099_, _34719_);
  and _51805_ (_07101_, _07100_, _07089_);
  or _51806_ (_07102_, _07101_, _07079_);
  and _51807_ (_07103_, _07102_, _34700_);
  and _51808_ (_07104_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and _51809_ (_07105_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or _51810_ (_07106_, _07105_, _07104_);
  and _51811_ (_07107_, _07106_, _34581_);
  and _51812_ (_07108_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and _51813_ (_07109_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or _51814_ (_07110_, _07109_, _07108_);
  and _51815_ (_07111_, _07110_, _34796_);
  or _51816_ (_07112_, _07111_, _07107_);
  or _51817_ (_07113_, _07112_, _34790_);
  and _51818_ (_07114_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and _51819_ (_07115_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or _51820_ (_07116_, _07115_, _07114_);
  and _51821_ (_07117_, _07116_, _34581_);
  and _51822_ (_07118_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and _51823_ (_07119_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or _51824_ (_07120_, _07119_, _07118_);
  and _51825_ (_07121_, _07120_, _34796_);
  or _51826_ (_07122_, _07121_, _07117_);
  or _51827_ (_07123_, _07122_, _34772_);
  and _51828_ (_07124_, _07123_, _34803_);
  and _51829_ (_07125_, _07124_, _07113_);
  or _51830_ (_07126_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or _51831_ (_07127_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  and _51832_ (_07128_, _07127_, _34796_);
  and _51833_ (_07129_, _07128_, _07126_);
  or _51834_ (_07130_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or _51835_ (_07131_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  and _51836_ (_07132_, _07131_, _34581_);
  and _51837_ (_07133_, _07132_, _07130_);
  or _51838_ (_07134_, _07133_, _07129_);
  or _51839_ (_07135_, _07134_, _34790_);
  or _51840_ (_07136_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or _51841_ (_07137_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and _51842_ (_07138_, _07137_, _34796_);
  and _51843_ (_07139_, _07138_, _07136_);
  or _51844_ (_07140_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or _51845_ (_07141_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and _51846_ (_07142_, _07141_, _34581_);
  and _51847_ (_07143_, _07142_, _07140_);
  or _51848_ (_07144_, _07143_, _07139_);
  or _51849_ (_07145_, _07144_, _34772_);
  and _51850_ (_07146_, _07145_, _34719_);
  and _51851_ (_07147_, _07146_, _07135_);
  or _51852_ (_07148_, _07147_, _07125_);
  and _51853_ (_07149_, _07148_, _34789_);
  or _51854_ (_07150_, _07149_, _07103_);
  and _51855_ (_07151_, _07150_, _34840_);
  and _51856_ (_07152_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and _51857_ (_07153_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or _51858_ (_07154_, _07153_, _07152_);
  and _51859_ (_07155_, _07154_, _34581_);
  and _51860_ (_07156_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and _51861_ (_07157_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or _51862_ (_07158_, _07157_, _07156_);
  and _51863_ (_07159_, _07158_, _34796_);
  or _51864_ (_07160_, _07159_, _07155_);
  and _51865_ (_07161_, _07160_, _34772_);
  and _51866_ (_07162_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and _51867_ (_07163_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _51868_ (_07164_, _07163_, _07162_);
  and _51869_ (_07165_, _07164_, _34581_);
  and _51870_ (_07166_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and _51871_ (_07167_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or _51872_ (_07168_, _07167_, _07166_);
  and _51873_ (_07169_, _07168_, _34796_);
  or _51874_ (_07170_, _07169_, _07165_);
  and _51875_ (_07171_, _07170_, _34790_);
  or _51876_ (_07172_, _07171_, _07161_);
  and _51877_ (_07173_, _07172_, _34803_);
  or _51878_ (_07174_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or _51879_ (_07175_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and _51880_ (_07176_, _07175_, _34796_);
  and _51881_ (_07177_, _07176_, _07174_);
  or _51882_ (_07178_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or _51883_ (_07179_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and _51884_ (_07180_, _07179_, _34581_);
  and _51885_ (_07181_, _07180_, _07178_);
  or _51886_ (_07182_, _07181_, _07177_);
  and _51887_ (_07183_, _07182_, _34772_);
  or _51888_ (_07184_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or _51889_ (_07185_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and _51890_ (_07186_, _07185_, _34796_);
  and _51891_ (_07187_, _07186_, _07184_);
  or _51892_ (_07188_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or _51893_ (_07189_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and _51894_ (_07190_, _07189_, _34581_);
  and _51895_ (_07191_, _07190_, _07188_);
  or _51896_ (_07192_, _07191_, _07187_);
  and _51897_ (_07193_, _07192_, _34790_);
  or _51898_ (_07194_, _07193_, _07183_);
  and _51899_ (_07195_, _07194_, _34719_);
  or _51900_ (_07196_, _07195_, _07173_);
  and _51901_ (_07197_, _07196_, _34789_);
  and _51902_ (_07198_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and _51903_ (_07199_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or _51904_ (_07200_, _07199_, _07198_);
  and _51905_ (_07201_, _07200_, _34581_);
  and _51906_ (_07202_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  and _51907_ (_07203_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or _51908_ (_07204_, _07203_, _07202_);
  and _51909_ (_07205_, _07204_, _34796_);
  or _51910_ (_07206_, _07205_, _07201_);
  and _51911_ (_07207_, _07206_, _34772_);
  and _51912_ (_07208_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and _51913_ (_07209_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or _51914_ (_07210_, _07209_, _07208_);
  and _51915_ (_07211_, _07210_, _34581_);
  and _51916_ (_07212_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and _51917_ (_07213_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or _51918_ (_07214_, _07213_, _07212_);
  and _51919_ (_07215_, _07214_, _34796_);
  or _51920_ (_07216_, _07215_, _07211_);
  and _51921_ (_07217_, _07216_, _34790_);
  or _51922_ (_07218_, _07217_, _07207_);
  and _51923_ (_07219_, _07218_, _34803_);
  or _51924_ (_07220_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or _51925_ (_07221_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and _51926_ (_07222_, _07221_, _07220_);
  and _51927_ (_07223_, _07222_, _34581_);
  or _51928_ (_07224_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or _51929_ (_07225_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and _51930_ (_07226_, _07225_, _07224_);
  and _51931_ (_07227_, _07226_, _34796_);
  or _51932_ (_07228_, _07227_, _07223_);
  and _51933_ (_07229_, _07228_, _34772_);
  or _51934_ (_07230_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or _51935_ (_07231_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and _51936_ (_07232_, _07231_, _07230_);
  and _51937_ (_07233_, _07232_, _34581_);
  or _51938_ (_07234_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or _51939_ (_07235_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and _51940_ (_07236_, _07235_, _07234_);
  and _51941_ (_07237_, _07236_, _34796_);
  or _51942_ (_07238_, _07237_, _07233_);
  and _51943_ (_07239_, _07238_, _34790_);
  or _51944_ (_07240_, _07239_, _07229_);
  and _51945_ (_07241_, _07240_, _34719_);
  or _51946_ (_07242_, _07241_, _07219_);
  and _51947_ (_07243_, _07242_, _34700_);
  or _51948_ (_07244_, _07243_, _07197_);
  and _51949_ (_07245_, _07244_, _34638_);
  or _51950_ (_07246_, _07245_, _07151_);
  or _51951_ (_07247_, _07246_, _34692_);
  and _51952_ (_07248_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and _51953_ (_07249_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or _51954_ (_07250_, _07249_, _07248_);
  and _51955_ (_07251_, _07250_, _34581_);
  and _51956_ (_07252_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and _51957_ (_07253_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or _51958_ (_07254_, _07253_, _07252_);
  and _51959_ (_07255_, _07254_, _34796_);
  or _51960_ (_07256_, _07255_, _07251_);
  or _51961_ (_07257_, _07256_, _34790_);
  and _51962_ (_07258_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and _51963_ (_07259_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or _51964_ (_07260_, _07259_, _07258_);
  and _51965_ (_07261_, _07260_, _34581_);
  and _51966_ (_07262_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and _51967_ (_07263_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or _51968_ (_07264_, _07263_, _07262_);
  and _51969_ (_07265_, _07264_, _34796_);
  or _51970_ (_07266_, _07265_, _07261_);
  or _51971_ (_07267_, _07266_, _34772_);
  and _51972_ (_07268_, _07267_, _34803_);
  and _51973_ (_07269_, _07268_, _07257_);
  or _51974_ (_07270_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or _51975_ (_07271_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and _51976_ (_07272_, _07271_, _34796_);
  and _51977_ (_07273_, _07272_, _07270_);
  or _51978_ (_07274_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or _51979_ (_07275_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and _51980_ (_07276_, _07275_, _34581_);
  and _51981_ (_07277_, _07276_, _07274_);
  or _51982_ (_07278_, _07277_, _07273_);
  or _51983_ (_07279_, _07278_, _34790_);
  or _51984_ (_07280_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or _51985_ (_07281_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and _51986_ (_07282_, _07281_, _34796_);
  and _51987_ (_07283_, _07282_, _07280_);
  or _51988_ (_07284_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or _51989_ (_07285_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  and _51990_ (_07286_, _07285_, _34581_);
  and _51991_ (_07287_, _07286_, _07284_);
  or _51992_ (_07288_, _07287_, _07283_);
  or _51993_ (_07289_, _07288_, _34772_);
  and _51994_ (_07290_, _07289_, _34719_);
  and _51995_ (_07291_, _07290_, _07279_);
  or _51996_ (_07292_, _07291_, _07269_);
  and _51997_ (_07293_, _07292_, _34789_);
  and _51998_ (_07294_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and _51999_ (_07295_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or _52000_ (_07296_, _07295_, _07294_);
  and _52001_ (_07297_, _07296_, _34581_);
  and _52002_ (_07298_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and _52003_ (_07299_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or _52004_ (_07300_, _07299_, _07298_);
  and _52005_ (_07301_, _07300_, _34796_);
  or _52006_ (_07302_, _07301_, _07297_);
  or _52007_ (_07303_, _07302_, _34790_);
  and _52008_ (_07304_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and _52009_ (_07305_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or _52010_ (_07306_, _07305_, _07304_);
  and _52011_ (_07307_, _07306_, _34581_);
  and _52012_ (_07308_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and _52013_ (_07309_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or _52014_ (_07310_, _07309_, _07308_);
  and _52015_ (_07311_, _07310_, _34796_);
  or _52016_ (_07312_, _07311_, _07307_);
  or _52017_ (_07313_, _07312_, _34772_);
  and _52018_ (_07314_, _07313_, _34803_);
  and _52019_ (_07315_, _07314_, _07303_);
  or _52020_ (_07316_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or _52021_ (_07317_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and _52022_ (_07318_, _07317_, _07316_);
  and _52023_ (_07319_, _07318_, _34581_);
  or _52024_ (_07320_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or _52025_ (_07321_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and _52026_ (_07322_, _07321_, _07320_);
  and _52027_ (_07323_, _07322_, _34796_);
  or _52028_ (_07324_, _07323_, _07319_);
  or _52029_ (_07325_, _07324_, _34790_);
  or _52030_ (_07326_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or _52031_ (_07327_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and _52032_ (_07328_, _07327_, _07326_);
  and _52033_ (_07329_, _07328_, _34581_);
  or _52034_ (_07330_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or _52035_ (_07331_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and _52036_ (_07332_, _07331_, _07330_);
  and _52037_ (_07333_, _07332_, _34796_);
  or _52038_ (_07334_, _07333_, _07329_);
  or _52039_ (_07335_, _07334_, _34772_);
  and _52040_ (_07336_, _07335_, _34719_);
  and _52041_ (_07337_, _07336_, _07325_);
  or _52042_ (_07338_, _07337_, _07315_);
  and _52043_ (_07339_, _07338_, _34700_);
  or _52044_ (_07340_, _07339_, _07293_);
  and _52045_ (_07341_, _07340_, _34840_);
  or _52046_ (_07342_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or _52047_ (_07343_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and _52048_ (_07344_, _07343_, _07342_);
  and _52049_ (_07345_, _07344_, _34581_);
  or _52050_ (_07346_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or _52051_ (_07347_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  and _52052_ (_07348_, _07347_, _07346_);
  and _52053_ (_07349_, _07348_, _34796_);
  or _52054_ (_07350_, _07349_, _07345_);
  and _52055_ (_07351_, _07350_, _34790_);
  or _52056_ (_07352_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or _52057_ (_07353_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and _52058_ (_07354_, _07353_, _07352_);
  and _52059_ (_07355_, _07354_, _34581_);
  or _52060_ (_07356_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or _52061_ (_07357_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and _52062_ (_07358_, _07357_, _07356_);
  and _52063_ (_07359_, _07358_, _34796_);
  or _52064_ (_07360_, _07359_, _07355_);
  and _52065_ (_07361_, _07360_, _34772_);
  or _52066_ (_07362_, _07361_, _07351_);
  and _52067_ (_07363_, _07362_, _34719_);
  and _52068_ (_07364_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and _52069_ (_07365_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or _52070_ (_07366_, _07365_, _07364_);
  and _52071_ (_07367_, _07366_, _34581_);
  and _52072_ (_07368_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and _52073_ (_07369_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or _52074_ (_07370_, _07369_, _07368_);
  and _52075_ (_07371_, _07370_, _34796_);
  or _52076_ (_07372_, _07371_, _07367_);
  and _52077_ (_07373_, _07372_, _34790_);
  and _52078_ (_07374_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and _52079_ (_07375_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or _52080_ (_07376_, _07375_, _07374_);
  and _52081_ (_07377_, _07376_, _34581_);
  and _52082_ (_07378_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and _52083_ (_07379_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or _52084_ (_07380_, _07379_, _07378_);
  and _52085_ (_07381_, _07380_, _34796_);
  or _52086_ (_07382_, _07381_, _07377_);
  and _52087_ (_07383_, _07382_, _34772_);
  or _52088_ (_07384_, _07383_, _07373_);
  and _52089_ (_07385_, _07384_, _34803_);
  or _52090_ (_07386_, _07385_, _07363_);
  and _52091_ (_07387_, _07386_, _34700_);
  or _52092_ (_07388_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or _52093_ (_07389_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  and _52094_ (_07390_, _07389_, _34796_);
  and _52095_ (_07391_, _07390_, _07388_);
  or _52096_ (_07392_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or _52097_ (_07393_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and _52098_ (_07394_, _07393_, _34581_);
  and _52099_ (_07395_, _07394_, _07392_);
  or _52100_ (_07396_, _07395_, _07391_);
  and _52101_ (_07397_, _07396_, _34790_);
  or _52102_ (_07398_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or _52103_ (_07399_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  and _52104_ (_07400_, _07399_, _34796_);
  and _52105_ (_07401_, _07400_, _07398_);
  or _52106_ (_07402_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or _52107_ (_07403_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and _52108_ (_07404_, _07403_, _34581_);
  and _52109_ (_07405_, _07404_, _07402_);
  or _52110_ (_07406_, _07405_, _07401_);
  and _52111_ (_07407_, _07406_, _34772_);
  or _52112_ (_07408_, _07407_, _07397_);
  and _52113_ (_07409_, _07408_, _34719_);
  and _52114_ (_07410_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and _52115_ (_07411_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or _52116_ (_07412_, _07411_, _07410_);
  and _52117_ (_07413_, _07412_, _34581_);
  and _52118_ (_07414_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  and _52119_ (_07415_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or _52120_ (_07416_, _07415_, _07414_);
  and _52121_ (_07417_, _07416_, _34796_);
  or _52122_ (_07418_, _07417_, _07413_);
  and _52123_ (_07419_, _07418_, _34790_);
  and _52124_ (_07420_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  and _52125_ (_07421_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or _52126_ (_07422_, _07421_, _07420_);
  and _52127_ (_07423_, _07422_, _34581_);
  and _52128_ (_07424_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and _52129_ (_07425_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or _52130_ (_07426_, _07425_, _07424_);
  and _52131_ (_07427_, _07426_, _34796_);
  or _52132_ (_07428_, _07427_, _07423_);
  and _52133_ (_07429_, _07428_, _34772_);
  or _52134_ (_07430_, _07429_, _07419_);
  and _52135_ (_07431_, _07430_, _34803_);
  or _52136_ (_07432_, _07431_, _07409_);
  and _52137_ (_07433_, _07432_, _34789_);
  or _52138_ (_07434_, _07433_, _07387_);
  and _52139_ (_07435_, _07434_, _34638_);
  or _52140_ (_07436_, _07435_, _07341_);
  or _52141_ (_07437_, _07436_, _34985_);
  and _52142_ (_07438_, _07437_, _07247_);
  or _52143_ (_07439_, _07438_, _34346_);
  and _52144_ (_07440_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and _52145_ (_07441_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or _52146_ (_07442_, _07441_, _07440_);
  and _52147_ (_07443_, _07442_, _34796_);
  and _52148_ (_07444_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and _52149_ (_07445_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or _52150_ (_07446_, _07445_, _07444_);
  and _52151_ (_07447_, _07446_, _34581_);
  or _52152_ (_07448_, _07447_, _07443_);
  or _52153_ (_07449_, _07448_, _34790_);
  and _52154_ (_07450_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and _52155_ (_07451_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or _52156_ (_07452_, _07451_, _07450_);
  and _52157_ (_07453_, _07452_, _34796_);
  and _52158_ (_07454_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and _52159_ (_07455_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or _52160_ (_07456_, _07455_, _07454_);
  and _52161_ (_07457_, _07456_, _34581_);
  or _52162_ (_07458_, _07457_, _07453_);
  or _52163_ (_07459_, _07458_, _34772_);
  and _52164_ (_07460_, _07459_, _34803_);
  and _52165_ (_07461_, _07460_, _07449_);
  or _52166_ (_07462_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or _52167_ (_07463_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and _52168_ (_07464_, _07463_, _34581_);
  and _52169_ (_07465_, _07464_, _07462_);
  or _52170_ (_07466_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or _52171_ (_07467_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and _52172_ (_07468_, _07467_, _34796_);
  and _52173_ (_07469_, _07468_, _07466_);
  or _52174_ (_07470_, _07469_, _07465_);
  or _52175_ (_07471_, _07470_, _34790_);
  or _52176_ (_07472_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or _52177_ (_07473_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and _52178_ (_07474_, _07473_, _34581_);
  and _52179_ (_07475_, _07474_, _07472_);
  or _52180_ (_07476_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or _52181_ (_07477_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and _52182_ (_07478_, _07477_, _34796_);
  and _52183_ (_07479_, _07478_, _07476_);
  or _52184_ (_07480_, _07479_, _07475_);
  or _52185_ (_07481_, _07480_, _34772_);
  and _52186_ (_07482_, _07481_, _34719_);
  and _52187_ (_07483_, _07482_, _07471_);
  or _52188_ (_07484_, _07483_, _07461_);
  and _52189_ (_07485_, _07484_, _34789_);
  and _52190_ (_07486_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and _52191_ (_07487_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or _52192_ (_07488_, _07487_, _34581_);
  or _52193_ (_07489_, _07488_, _07486_);
  and _52194_ (_07490_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and _52195_ (_07491_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or _52196_ (_07492_, _07491_, _34796_);
  or _52197_ (_07493_, _07492_, _07490_);
  and _52198_ (_07494_, _07493_, _07489_);
  or _52199_ (_07495_, _07494_, _34790_);
  and _52200_ (_07496_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and _52201_ (_07497_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or _52202_ (_07498_, _07497_, _34581_);
  or _52203_ (_07499_, _07498_, _07496_);
  and _52204_ (_07500_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and _52205_ (_07501_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or _52206_ (_07502_, _07501_, _34796_);
  or _52207_ (_07503_, _07502_, _07500_);
  and _52208_ (_07504_, _07503_, _07499_);
  or _52209_ (_07505_, _07504_, _34772_);
  and _52210_ (_07506_, _07505_, _34803_);
  and _52211_ (_07507_, _07506_, _07495_);
  or _52212_ (_07508_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or _52213_ (_07509_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and _52214_ (_07510_, _07509_, _07508_);
  or _52215_ (_07511_, _07510_, _34796_);
  or _52216_ (_07512_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or _52217_ (_07513_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and _52218_ (_07514_, _07513_, _07512_);
  or _52219_ (_07515_, _07514_, _34581_);
  and _52220_ (_07516_, _07515_, _07511_);
  or _52221_ (_07517_, _07516_, _34790_);
  or _52222_ (_07518_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or _52223_ (_07519_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and _52224_ (_07520_, _07519_, _07518_);
  or _52225_ (_07521_, _07520_, _34796_);
  or _52226_ (_07522_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or _52227_ (_07523_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and _52228_ (_07524_, _07523_, _07522_);
  or _52229_ (_07525_, _07524_, _34581_);
  and _52230_ (_07526_, _07525_, _07521_);
  or _52231_ (_07527_, _07526_, _34772_);
  and _52232_ (_07528_, _07527_, _34719_);
  and _52233_ (_07529_, _07528_, _07517_);
  or _52234_ (_07530_, _07529_, _07507_);
  and _52235_ (_07531_, _07530_, _34700_);
  or _52236_ (_07532_, _07531_, _07485_);
  and _52237_ (_07533_, _07532_, _34840_);
  and _52238_ (_07534_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  and _52239_ (_07535_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  or _52240_ (_07536_, _07535_, _07534_);
  and _52241_ (_07537_, _07536_, _34581_);
  and _52242_ (_07538_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  and _52243_ (_07539_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  or _52244_ (_07540_, _07539_, _07538_);
  and _52245_ (_07541_, _07540_, _34796_);
  or _52246_ (_07542_, _07541_, _07537_);
  and _52247_ (_07543_, _07542_, _34772_);
  and _52248_ (_07544_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  and _52249_ (_07545_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  or _52250_ (_07546_, _07545_, _07544_);
  and _52251_ (_07547_, _07546_, _34581_);
  and _52252_ (_07548_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  and _52253_ (_07549_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  or _52254_ (_07550_, _07549_, _07548_);
  and _52255_ (_07551_, _07550_, _34796_);
  or _52256_ (_07552_, _07551_, _07547_);
  and _52257_ (_07553_, _07552_, _34790_);
  or _52258_ (_07554_, _07553_, _07543_);
  and _52259_ (_07555_, _07554_, _34803_);
  or _52260_ (_07556_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  or _52261_ (_07557_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  and _52262_ (_07558_, _07557_, _07556_);
  and _52263_ (_07559_, _07558_, _34581_);
  or _52264_ (_07560_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  or _52265_ (_07561_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  and _52266_ (_07562_, _07561_, _07560_);
  and _52267_ (_07563_, _07562_, _34796_);
  or _52268_ (_07564_, _07563_, _07559_);
  and _52269_ (_07565_, _07564_, _34772_);
  or _52270_ (_07566_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  or _52271_ (_07567_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  and _52272_ (_07568_, _07567_, _07566_);
  and _52273_ (_07569_, _07568_, _34581_);
  or _52274_ (_07570_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  or _52275_ (_07571_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  and _52276_ (_07572_, _07571_, _07570_);
  and _52277_ (_07573_, _07572_, _34796_);
  or _52278_ (_07574_, _07573_, _07569_);
  and _52279_ (_07575_, _07574_, _34790_);
  or _52280_ (_07576_, _07575_, _07565_);
  and _52281_ (_07577_, _07576_, _34719_);
  or _52282_ (_07578_, _07577_, _07555_);
  and _52283_ (_07579_, _07578_, _34789_);
  and _52284_ (_07580_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and _52285_ (_07581_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or _52286_ (_07582_, _07581_, _07580_);
  and _52287_ (_07583_, _07582_, _34581_);
  and _52288_ (_07584_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and _52289_ (_07585_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or _52290_ (_07586_, _07585_, _07584_);
  and _52291_ (_07587_, _07586_, _34796_);
  or _52292_ (_07588_, _07587_, _07583_);
  and _52293_ (_07589_, _07588_, _34772_);
  and _52294_ (_07590_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and _52295_ (_07591_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or _52296_ (_07592_, _07591_, _07590_);
  and _52297_ (_07593_, _07592_, _34581_);
  and _52298_ (_07594_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and _52299_ (_07595_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or _52300_ (_07596_, _07595_, _07594_);
  and _52301_ (_07597_, _07596_, _34796_);
  or _52302_ (_07598_, _07597_, _07593_);
  and _52303_ (_07599_, _07598_, _34790_);
  or _52304_ (_07600_, _07599_, _07589_);
  and _52305_ (_07601_, _07600_, _34803_);
  or _52306_ (_07602_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or _52307_ (_07603_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and _52308_ (_07604_, _07603_, _07602_);
  and _52309_ (_07605_, _07604_, _34581_);
  or _52310_ (_07606_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or _52311_ (_07607_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and _52312_ (_07608_, _07607_, _07606_);
  and _52313_ (_07609_, _07608_, _34796_);
  or _52314_ (_07610_, _07609_, _07605_);
  and _52315_ (_07611_, _07610_, _34772_);
  or _52316_ (_07612_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or _52317_ (_07613_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and _52318_ (_07614_, _07613_, _07612_);
  and _52319_ (_07615_, _07614_, _34581_);
  or _52320_ (_07616_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or _52321_ (_07617_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and _52322_ (_07618_, _07617_, _07616_);
  and _52323_ (_07619_, _07618_, _34796_);
  or _52324_ (_07620_, _07619_, _07615_);
  and _52325_ (_07621_, _07620_, _34790_);
  or _52326_ (_07622_, _07621_, _07611_);
  and _52327_ (_07623_, _07622_, _34719_);
  or _52328_ (_07624_, _07623_, _07601_);
  and _52329_ (_07625_, _07624_, _34700_);
  or _52330_ (_07626_, _07625_, _07579_);
  and _52331_ (_07627_, _07626_, _34638_);
  or _52332_ (_07628_, _07627_, _07533_);
  or _52333_ (_07629_, _07628_, _34692_);
  and _52334_ (_07630_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and _52335_ (_07631_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or _52336_ (_07632_, _07631_, _07630_);
  and _52337_ (_07633_, _07632_, _34581_);
  and _52338_ (_07634_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and _52339_ (_07635_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or _52340_ (_07636_, _07635_, _07634_);
  and _52341_ (_07637_, _07636_, _34796_);
  or _52342_ (_07638_, _07637_, _07633_);
  or _52343_ (_07639_, _07638_, _34790_);
  and _52344_ (_07640_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and _52345_ (_07641_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or _52346_ (_07642_, _07641_, _07640_);
  and _52347_ (_07643_, _07642_, _34581_);
  and _52348_ (_07644_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and _52349_ (_07645_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or _52350_ (_07646_, _07645_, _07644_);
  and _52351_ (_07647_, _07646_, _34796_);
  or _52352_ (_07648_, _07647_, _07643_);
  or _52353_ (_07649_, _07648_, _34772_);
  and _52354_ (_07650_, _07649_, _34803_);
  and _52355_ (_07651_, _07650_, _07639_);
  or _52356_ (_07652_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or _52357_ (_07653_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and _52358_ (_07654_, _07653_, _34796_);
  and _52359_ (_07655_, _07654_, _07652_);
  or _52360_ (_07656_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or _52361_ (_07657_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and _52362_ (_07658_, _07657_, _34581_);
  and _52363_ (_07659_, _07658_, _07656_);
  or _52364_ (_07660_, _07659_, _07655_);
  or _52365_ (_07661_, _07660_, _34790_);
  or _52366_ (_07662_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or _52367_ (_07663_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and _52368_ (_07664_, _07663_, _34796_);
  and _52369_ (_07665_, _07664_, _07662_);
  or _52370_ (_07666_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or _52371_ (_07667_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and _52372_ (_07668_, _07667_, _34581_);
  and _52373_ (_07669_, _07668_, _07666_);
  or _52374_ (_07670_, _07669_, _07665_);
  or _52375_ (_07671_, _07670_, _34772_);
  and _52376_ (_07672_, _07671_, _34719_);
  and _52377_ (_07673_, _07672_, _07661_);
  or _52378_ (_07674_, _07673_, _07651_);
  and _52379_ (_07675_, _07674_, _34789_);
  and _52380_ (_07676_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and _52381_ (_07677_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or _52382_ (_07678_, _07677_, _07676_);
  and _52383_ (_07679_, _07678_, _34581_);
  and _52384_ (_07680_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and _52385_ (_07681_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or _52386_ (_07682_, _07681_, _07680_);
  and _52387_ (_07683_, _07682_, _34796_);
  or _52388_ (_07684_, _07683_, _07679_);
  or _52389_ (_07685_, _07684_, _34790_);
  and _52390_ (_07686_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and _52391_ (_07687_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or _52392_ (_07688_, _07687_, _07686_);
  and _52393_ (_07689_, _07688_, _34581_);
  and _52394_ (_07690_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and _52395_ (_07691_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or _52396_ (_07692_, _07691_, _07690_);
  and _52397_ (_07693_, _07692_, _34796_);
  or _52398_ (_07694_, _07693_, _07689_);
  or _52399_ (_07695_, _07694_, _34772_);
  and _52400_ (_07696_, _07695_, _34803_);
  and _52401_ (_07697_, _07696_, _07685_);
  or _52402_ (_07698_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or _52403_ (_07699_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and _52404_ (_07700_, _07699_, _07698_);
  and _52405_ (_07701_, _07700_, _34581_);
  or _52406_ (_07702_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or _52407_ (_07703_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and _52408_ (_07704_, _07703_, _07702_);
  and _52409_ (_07705_, _07704_, _34796_);
  or _52410_ (_07706_, _07705_, _07701_);
  or _52411_ (_07707_, _07706_, _34790_);
  or _52412_ (_07708_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or _52413_ (_07709_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and _52414_ (_07710_, _07709_, _07708_);
  and _52415_ (_07711_, _07710_, _34581_);
  or _52416_ (_07712_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or _52417_ (_07713_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and _52418_ (_07714_, _07713_, _07712_);
  and _52419_ (_07715_, _07714_, _34796_);
  or _52420_ (_07716_, _07715_, _07711_);
  or _52421_ (_07717_, _07716_, _34772_);
  and _52422_ (_07718_, _07717_, _34719_);
  and _52423_ (_07719_, _07718_, _07707_);
  or _52424_ (_07720_, _07719_, _07697_);
  and _52425_ (_07721_, _07720_, _34700_);
  or _52426_ (_07722_, _07721_, _07675_);
  and _52427_ (_07723_, _07722_, _34840_);
  or _52428_ (_07724_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or _52429_ (_07725_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and _52430_ (_07726_, _07725_, _07724_);
  and _52431_ (_07727_, _07726_, _34581_);
  or _52432_ (_07728_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or _52433_ (_07729_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and _52434_ (_07730_, _07729_, _07728_);
  and _52435_ (_07731_, _07730_, _34796_);
  or _52436_ (_07732_, _07731_, _07727_);
  and _52437_ (_07733_, _07732_, _34790_);
  or _52438_ (_07734_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or _52439_ (_07735_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and _52440_ (_07736_, _07735_, _07734_);
  and _52441_ (_07737_, _07736_, _34581_);
  or _52442_ (_07738_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or _52443_ (_07739_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and _52444_ (_07740_, _07739_, _07738_);
  and _52445_ (_07741_, _07740_, _34796_);
  or _52446_ (_07742_, _07741_, _07737_);
  and _52447_ (_07743_, _07742_, _34772_);
  or _52448_ (_07744_, _07743_, _07733_);
  and _52449_ (_07745_, _07744_, _34719_);
  and _52450_ (_07746_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and _52451_ (_07747_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or _52452_ (_07748_, _07747_, _07746_);
  and _52453_ (_07749_, _07748_, _34581_);
  and _52454_ (_07750_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and _52455_ (_07751_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or _52456_ (_07752_, _07751_, _07750_);
  and _52457_ (_07753_, _07752_, _34796_);
  or _52458_ (_07754_, _07753_, _07749_);
  and _52459_ (_07755_, _07754_, _34790_);
  and _52460_ (_07756_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and _52461_ (_07757_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or _52462_ (_07758_, _07757_, _07756_);
  and _52463_ (_07759_, _07758_, _34581_);
  and _52464_ (_07760_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and _52465_ (_07761_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or _52466_ (_07762_, _07761_, _07760_);
  and _52467_ (_07763_, _07762_, _34796_);
  or _52468_ (_07764_, _07763_, _07759_);
  and _52469_ (_07765_, _07764_, _34772_);
  or _52470_ (_07766_, _07765_, _07755_);
  and _52471_ (_07767_, _07766_, _34803_);
  or _52472_ (_07768_, _07767_, _07745_);
  and _52473_ (_07769_, _07768_, _34700_);
  or _52474_ (_07770_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or _52475_ (_07771_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and _52476_ (_07772_, _07771_, _34796_);
  and _52477_ (_07773_, _07772_, _07770_);
  or _52478_ (_07774_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or _52479_ (_07775_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and _52480_ (_07776_, _07775_, _34581_);
  and _52481_ (_07777_, _07776_, _07774_);
  or _52482_ (_07778_, _07777_, _07773_);
  and _52483_ (_07779_, _07778_, _34790_);
  or _52484_ (_07780_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or _52485_ (_07781_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and _52486_ (_07782_, _07781_, _34796_);
  and _52487_ (_07783_, _07782_, _07780_);
  or _52488_ (_07784_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or _52489_ (_07785_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and _52490_ (_07786_, _07785_, _34581_);
  and _52491_ (_07787_, _07786_, _07784_);
  or _52492_ (_07788_, _07787_, _07783_);
  and _52493_ (_07789_, _07788_, _34772_);
  or _52494_ (_07790_, _07789_, _07779_);
  and _52495_ (_07791_, _07790_, _34719_);
  and _52496_ (_07792_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and _52497_ (_07793_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or _52498_ (_07794_, _07793_, _07792_);
  and _52499_ (_07795_, _07794_, _34581_);
  and _52500_ (_07796_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and _52501_ (_07797_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or _52502_ (_07798_, _07797_, _07796_);
  and _52503_ (_07799_, _07798_, _34796_);
  or _52504_ (_07800_, _07799_, _07795_);
  and _52505_ (_07801_, _07800_, _34790_);
  and _52506_ (_07802_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and _52507_ (_07803_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or _52508_ (_07804_, _07803_, _07802_);
  and _52509_ (_07805_, _07804_, _34581_);
  and _52510_ (_07806_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and _52511_ (_07807_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or _52512_ (_07808_, _07807_, _07806_);
  and _52513_ (_07809_, _07808_, _34796_);
  or _52514_ (_07810_, _07809_, _07805_);
  and _52515_ (_07811_, _07810_, _34772_);
  or _52516_ (_07812_, _07811_, _07801_);
  and _52517_ (_07813_, _07812_, _34803_);
  or _52518_ (_07814_, _07813_, _07791_);
  and _52519_ (_07815_, _07814_, _34789_);
  or _52520_ (_07816_, _07815_, _07769_);
  and _52521_ (_07817_, _07816_, _34638_);
  or _52522_ (_07818_, _07817_, _07723_);
  or _52523_ (_07819_, _07818_, _34985_);
  and _52524_ (_07820_, _07819_, _07629_);
  or _52525_ (_07821_, _07820_, _35178_);
  and _52526_ (_07822_, _07821_, _07439_);
  or _52527_ (_07823_, _07822_, _34788_);
  or _52528_ (_07824_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and _52529_ (_07825_, _07824_, _38997_);
  and _52530_ (_38984_[2], _07825_, _07823_);
  and _52531_ (_07826_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and _52532_ (_07827_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or _52533_ (_07828_, _07827_, _07826_);
  and _52534_ (_07829_, _07828_, _34796_);
  and _52535_ (_07830_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and _52536_ (_07831_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or _52537_ (_07832_, _07831_, _07830_);
  and _52538_ (_07833_, _07832_, _34581_);
  or _52539_ (_07834_, _07833_, _07829_);
  or _52540_ (_07835_, _07834_, _34790_);
  and _52541_ (_07836_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and _52542_ (_07837_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or _52543_ (_07838_, _07837_, _07836_);
  and _52544_ (_07839_, _07838_, _34796_);
  and _52545_ (_07840_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  and _52546_ (_07841_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or _52547_ (_07842_, _07841_, _07840_);
  and _52548_ (_07843_, _07842_, _34581_);
  or _52549_ (_07844_, _07843_, _07839_);
  or _52550_ (_07845_, _07844_, _34772_);
  and _52551_ (_07846_, _07845_, _34803_);
  and _52552_ (_07847_, _07846_, _07835_);
  or _52553_ (_07848_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or _52554_ (_07849_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and _52555_ (_07850_, _07849_, _34581_);
  and _52556_ (_07851_, _07850_, _07848_);
  or _52557_ (_07852_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or _52558_ (_07853_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and _52559_ (_07854_, _07853_, _34796_);
  and _52560_ (_07855_, _07854_, _07852_);
  or _52561_ (_07856_, _07855_, _07851_);
  or _52562_ (_07857_, _07856_, _34790_);
  or _52563_ (_07858_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or _52564_ (_07859_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and _52565_ (_07860_, _07859_, _34581_);
  and _52566_ (_07861_, _07860_, _07858_);
  or _52567_ (_07862_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or _52568_ (_07863_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  and _52569_ (_07864_, _07863_, _34796_);
  and _52570_ (_07865_, _07864_, _07862_);
  or _52571_ (_07866_, _07865_, _07861_);
  or _52572_ (_07867_, _07866_, _34772_);
  and _52573_ (_07868_, _07867_, _34719_);
  and _52574_ (_07869_, _07868_, _07857_);
  or _52575_ (_07870_, _07869_, _07847_);
  or _52576_ (_07871_, _07870_, _34700_);
  and _52577_ (_07872_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and _52578_ (_07873_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or _52579_ (_07874_, _07873_, _34581_);
  or _52580_ (_07875_, _07874_, _07872_);
  and _52581_ (_07876_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and _52582_ (_07877_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or _52583_ (_07878_, _07877_, _34796_);
  or _52584_ (_07879_, _07878_, _07876_);
  and _52585_ (_07880_, _07879_, _07875_);
  or _52586_ (_07881_, _07880_, _34790_);
  and _52587_ (_07882_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  and _52588_ (_07883_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or _52589_ (_07884_, _07883_, _34581_);
  or _52590_ (_07885_, _07884_, _07882_);
  and _52591_ (_07886_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and _52592_ (_07887_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or _52593_ (_07888_, _07887_, _34796_);
  or _52594_ (_07889_, _07888_, _07886_);
  and _52595_ (_07890_, _07889_, _07885_);
  or _52596_ (_07891_, _07890_, _34772_);
  and _52597_ (_07892_, _07891_, _34803_);
  and _52598_ (_07893_, _07892_, _07881_);
  or _52599_ (_07894_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or _52600_ (_07895_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  and _52601_ (_07896_, _07895_, _07894_);
  or _52602_ (_07897_, _07896_, _34796_);
  or _52603_ (_07898_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or _52604_ (_07899_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and _52605_ (_07900_, _07899_, _07898_);
  or _52606_ (_07901_, _07900_, _34581_);
  and _52607_ (_07902_, _07901_, _07897_);
  or _52608_ (_07903_, _07902_, _34790_);
  or _52609_ (_07904_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or _52610_ (_07905_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and _52611_ (_07906_, _07905_, _07904_);
  or _52612_ (_07907_, _07906_, _34796_);
  or _52613_ (_07908_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or _52614_ (_07909_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and _52615_ (_07910_, _07909_, _07908_);
  or _52616_ (_07911_, _07910_, _34581_);
  and _52617_ (_07912_, _07911_, _07907_);
  or _52618_ (_07913_, _07912_, _34772_);
  and _52619_ (_07914_, _07913_, _34719_);
  and _52620_ (_07915_, _07914_, _07903_);
  or _52621_ (_07916_, _07915_, _07893_);
  or _52622_ (_07917_, _07916_, _34789_);
  and _52623_ (_07918_, _07917_, _34840_);
  and _52624_ (_07919_, _07918_, _07871_);
  and _52625_ (_07920_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and _52626_ (_07921_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or _52627_ (_07922_, _07921_, _07920_);
  and _52628_ (_07923_, _07922_, _34581_);
  and _52629_ (_07924_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and _52630_ (_07925_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _52631_ (_07926_, _07925_, _07924_);
  and _52632_ (_07927_, _07926_, _34796_);
  or _52633_ (_07928_, _07927_, _07923_);
  and _52634_ (_07929_, _07928_, _34772_);
  and _52635_ (_07930_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and _52636_ (_07931_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or _52637_ (_07932_, _07931_, _07930_);
  and _52638_ (_07933_, _07932_, _34581_);
  and _52639_ (_07934_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and _52640_ (_07935_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _52641_ (_07936_, _07935_, _07934_);
  and _52642_ (_07937_, _07936_, _34796_);
  or _52643_ (_07938_, _07937_, _07933_);
  and _52644_ (_07939_, _07938_, _34790_);
  or _52645_ (_07940_, _07939_, _07929_);
  and _52646_ (_07941_, _07940_, _34803_);
  or _52647_ (_07942_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or _52648_ (_07943_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and _52649_ (_07944_, _07943_, _07942_);
  and _52650_ (_07945_, _07944_, _34581_);
  or _52651_ (_07946_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or _52652_ (_07947_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and _52653_ (_07948_, _07947_, _07946_);
  and _52654_ (_07949_, _07948_, _34796_);
  or _52655_ (_07950_, _07949_, _07945_);
  and _52656_ (_07951_, _07950_, _34772_);
  or _52657_ (_07952_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or _52658_ (_07953_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and _52659_ (_07954_, _07953_, _07952_);
  and _52660_ (_07955_, _07954_, _34581_);
  or _52661_ (_07956_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or _52662_ (_07957_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and _52663_ (_07958_, _07957_, _07956_);
  and _52664_ (_07959_, _07958_, _34796_);
  or _52665_ (_07960_, _07959_, _07955_);
  and _52666_ (_07961_, _07960_, _34790_);
  or _52667_ (_07962_, _07961_, _07951_);
  and _52668_ (_07963_, _07962_, _34719_);
  or _52669_ (_07964_, _07963_, _07941_);
  and _52670_ (_07965_, _07964_, _34789_);
  and _52671_ (_07966_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and _52672_ (_07967_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or _52673_ (_07968_, _07967_, _07966_);
  and _52674_ (_07969_, _07968_, _34581_);
  and _52675_ (_07970_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and _52676_ (_07971_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or _52677_ (_07972_, _07971_, _07970_);
  and _52678_ (_07973_, _07972_, _34796_);
  or _52679_ (_07974_, _07973_, _07969_);
  and _52680_ (_07975_, _07974_, _34772_);
  and _52681_ (_07976_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and _52682_ (_07977_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or _52683_ (_07978_, _07977_, _07976_);
  and _52684_ (_07979_, _07978_, _34581_);
  and _52685_ (_07980_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  and _52686_ (_07981_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or _52687_ (_07982_, _07981_, _07980_);
  and _52688_ (_07983_, _07982_, _34796_);
  or _52689_ (_07984_, _07983_, _07979_);
  and _52690_ (_07985_, _07984_, _34790_);
  or _52691_ (_07986_, _07985_, _07975_);
  and _52692_ (_07987_, _07986_, _34803_);
  or _52693_ (_07988_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or _52694_ (_07989_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  and _52695_ (_07990_, _07989_, _07988_);
  and _52696_ (_07991_, _07990_, _34581_);
  or _52697_ (_07992_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or _52698_ (_07993_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and _52699_ (_07994_, _07993_, _07992_);
  and _52700_ (_07995_, _07994_, _34796_);
  or _52701_ (_07996_, _07995_, _07991_);
  and _52702_ (_07997_, _07996_, _34772_);
  or _52703_ (_07998_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or _52704_ (_07999_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and _52705_ (_08000_, _07999_, _07998_);
  and _52706_ (_08001_, _08000_, _34581_);
  or _52707_ (_08002_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or _52708_ (_08003_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and _52709_ (_08004_, _08003_, _08002_);
  and _52710_ (_08005_, _08004_, _34796_);
  or _52711_ (_08006_, _08005_, _08001_);
  and _52712_ (_08007_, _08006_, _34790_);
  or _52713_ (_08008_, _08007_, _07997_);
  and _52714_ (_08009_, _08008_, _34719_);
  or _52715_ (_08010_, _08009_, _07987_);
  and _52716_ (_08011_, _08010_, _34700_);
  or _52717_ (_08012_, _08011_, _07965_);
  and _52718_ (_08013_, _08012_, _34638_);
  or _52719_ (_08014_, _08013_, _07919_);
  or _52720_ (_08015_, _08014_, _34692_);
  and _52721_ (_08016_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and _52722_ (_08017_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or _52723_ (_08018_, _08017_, _08016_);
  and _52724_ (_08019_, _08018_, _34581_);
  and _52725_ (_08020_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  and _52726_ (_08021_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or _52727_ (_08022_, _08021_, _08020_);
  and _52728_ (_08023_, _08022_, _34796_);
  or _52729_ (_08024_, _08023_, _08019_);
  or _52730_ (_08025_, _08024_, _34790_);
  and _52731_ (_08026_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and _52732_ (_08027_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or _52733_ (_08028_, _08027_, _08026_);
  and _52734_ (_08029_, _08028_, _34581_);
  and _52735_ (_08030_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and _52736_ (_08031_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or _52737_ (_08032_, _08031_, _08030_);
  and _52738_ (_08033_, _08032_, _34796_);
  or _52739_ (_08034_, _08033_, _08029_);
  or _52740_ (_08035_, _08034_, _34772_);
  and _52741_ (_08036_, _08035_, _34803_);
  and _52742_ (_08037_, _08036_, _08025_);
  or _52743_ (_08038_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or _52744_ (_08039_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  and _52745_ (_08040_, _08039_, _34796_);
  and _52746_ (_08041_, _08040_, _08038_);
  or _52747_ (_08042_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or _52748_ (_08043_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and _52749_ (_08044_, _08043_, _34581_);
  and _52750_ (_08045_, _08044_, _08042_);
  or _52751_ (_08046_, _08045_, _08041_);
  or _52752_ (_08047_, _08046_, _34790_);
  or _52753_ (_08048_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or _52754_ (_08049_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  and _52755_ (_08050_, _08049_, _34796_);
  and _52756_ (_08051_, _08050_, _08048_);
  or _52757_ (_08052_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or _52758_ (_08053_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and _52759_ (_08054_, _08053_, _34581_);
  and _52760_ (_08055_, _08054_, _08052_);
  or _52761_ (_08056_, _08055_, _08051_);
  or _52762_ (_08057_, _08056_, _34772_);
  and _52763_ (_08058_, _08057_, _34719_);
  and _52764_ (_08059_, _08058_, _08047_);
  or _52765_ (_08060_, _08059_, _08037_);
  and _52766_ (_08061_, _08060_, _34789_);
  and _52767_ (_08062_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and _52768_ (_08063_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or _52769_ (_08064_, _08063_, _08062_);
  and _52770_ (_08065_, _08064_, _34581_);
  and _52771_ (_08066_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and _52772_ (_08067_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or _52773_ (_08068_, _08067_, _08066_);
  and _52774_ (_08069_, _08068_, _34796_);
  or _52775_ (_08070_, _08069_, _08065_);
  or _52776_ (_08071_, _08070_, _34790_);
  and _52777_ (_08072_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and _52778_ (_08073_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or _52779_ (_08074_, _08073_, _08072_);
  and _52780_ (_08075_, _08074_, _34581_);
  and _52781_ (_08076_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and _52782_ (_08077_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or _52783_ (_08078_, _08077_, _08076_);
  and _52784_ (_08079_, _08078_, _34796_);
  or _52785_ (_08080_, _08079_, _08075_);
  or _52786_ (_08081_, _08080_, _34772_);
  and _52787_ (_08082_, _08081_, _34803_);
  and _52788_ (_08083_, _08082_, _08071_);
  or _52789_ (_08084_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or _52790_ (_08085_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and _52791_ (_08086_, _08085_, _08084_);
  and _52792_ (_08087_, _08086_, _34581_);
  or _52793_ (_08088_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or _52794_ (_08089_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and _52795_ (_08090_, _08089_, _08088_);
  and _52796_ (_08091_, _08090_, _34796_);
  or _52797_ (_08092_, _08091_, _08087_);
  or _52798_ (_08093_, _08092_, _34790_);
  or _52799_ (_08094_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or _52800_ (_08095_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and _52801_ (_08096_, _08095_, _08094_);
  and _52802_ (_08097_, _08096_, _34581_);
  or _52803_ (_08098_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or _52804_ (_08099_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and _52805_ (_08100_, _08099_, _08098_);
  and _52806_ (_08101_, _08100_, _34796_);
  or _52807_ (_08102_, _08101_, _08097_);
  or _52808_ (_08103_, _08102_, _34772_);
  and _52809_ (_08104_, _08103_, _34719_);
  and _52810_ (_08105_, _08104_, _08093_);
  or _52811_ (_08106_, _08105_, _08083_);
  and _52812_ (_08107_, _08106_, _34700_);
  or _52813_ (_08108_, _08107_, _08061_);
  and _52814_ (_08109_, _08108_, _34840_);
  or _52815_ (_08110_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or _52816_ (_08111_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and _52817_ (_08112_, _08111_, _08110_);
  and _52818_ (_08113_, _08112_, _34581_);
  or _52819_ (_08114_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or _52820_ (_08115_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  and _52821_ (_08116_, _08115_, _08114_);
  and _52822_ (_08117_, _08116_, _34796_);
  or _52823_ (_08118_, _08117_, _08113_);
  and _52824_ (_08119_, _08118_, _34790_);
  or _52825_ (_08120_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or _52826_ (_08121_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and _52827_ (_08122_, _08121_, _08120_);
  and _52828_ (_08123_, _08122_, _34581_);
  or _52829_ (_08124_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or _52830_ (_08125_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and _52831_ (_08126_, _08125_, _08124_);
  and _52832_ (_08127_, _08126_, _34796_);
  or _52833_ (_08128_, _08127_, _08123_);
  and _52834_ (_08129_, _08128_, _34772_);
  or _52835_ (_08130_, _08129_, _08119_);
  and _52836_ (_08131_, _08130_, _34719_);
  and _52837_ (_08132_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  and _52838_ (_08133_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or _52839_ (_08134_, _08133_, _08132_);
  and _52840_ (_08135_, _08134_, _34581_);
  and _52841_ (_08136_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and _52842_ (_08137_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or _52843_ (_08138_, _08137_, _08136_);
  and _52844_ (_08139_, _08138_, _34796_);
  or _52845_ (_08140_, _08139_, _08135_);
  and _52846_ (_08141_, _08140_, _34790_);
  and _52847_ (_08142_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and _52848_ (_08143_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or _52849_ (_08144_, _08143_, _08142_);
  and _52850_ (_08145_, _08144_, _34581_);
  and _52851_ (_08146_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and _52852_ (_08147_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or _52853_ (_08148_, _08147_, _08146_);
  and _52854_ (_08149_, _08148_, _34796_);
  or _52855_ (_08150_, _08149_, _08145_);
  and _52856_ (_08151_, _08150_, _34772_);
  or _52857_ (_08152_, _08151_, _08141_);
  and _52858_ (_08153_, _08152_, _34803_);
  or _52859_ (_08154_, _08153_, _08131_);
  and _52860_ (_08155_, _08154_, _34700_);
  or _52861_ (_08156_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or _52862_ (_08157_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  and _52863_ (_08158_, _08157_, _34796_);
  and _52864_ (_08159_, _08158_, _08156_);
  or _52865_ (_08160_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or _52866_ (_08161_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  and _52867_ (_08162_, _08161_, _34581_);
  and _52868_ (_08163_, _08162_, _08160_);
  or _52869_ (_08164_, _08163_, _08159_);
  and _52870_ (_08165_, _08164_, _34790_);
  or _52871_ (_08166_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or _52872_ (_08167_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and _52873_ (_08168_, _08167_, _34796_);
  and _52874_ (_08169_, _08168_, _08166_);
  or _52875_ (_08170_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or _52876_ (_08171_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  and _52877_ (_08172_, _08171_, _34581_);
  and _52878_ (_08173_, _08172_, _08170_);
  or _52879_ (_08174_, _08173_, _08169_);
  and _52880_ (_08175_, _08174_, _34772_);
  or _52881_ (_08176_, _08175_, _08165_);
  and _52882_ (_08177_, _08176_, _34719_);
  and _52883_ (_08178_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  and _52884_ (_08179_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or _52885_ (_08180_, _08179_, _08178_);
  and _52886_ (_08181_, _08180_, _34581_);
  and _52887_ (_08182_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and _52888_ (_08183_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or _52889_ (_08184_, _08183_, _08182_);
  and _52890_ (_08185_, _08184_, _34796_);
  or _52891_ (_08186_, _08185_, _08181_);
  and _52892_ (_08187_, _08186_, _34790_);
  and _52893_ (_08188_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  and _52894_ (_08189_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or _52895_ (_08190_, _08189_, _08188_);
  and _52896_ (_08191_, _08190_, _34581_);
  and _52897_ (_08192_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and _52898_ (_08193_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or _52899_ (_08194_, _08193_, _08192_);
  and _52900_ (_08195_, _08194_, _34796_);
  or _52901_ (_08196_, _08195_, _08191_);
  and _52902_ (_08197_, _08196_, _34772_);
  or _52903_ (_08198_, _08197_, _08187_);
  and _52904_ (_08199_, _08198_, _34803_);
  or _52905_ (_08200_, _08199_, _08177_);
  and _52906_ (_08201_, _08200_, _34789_);
  or _52907_ (_08202_, _08201_, _08155_);
  and _52908_ (_08203_, _08202_, _34638_);
  or _52909_ (_08204_, _08203_, _08109_);
  or _52910_ (_08205_, _08204_, _34985_);
  and _52911_ (_08206_, _08205_, _08015_);
  or _52912_ (_08207_, _08206_, _34346_);
  and _52913_ (_08208_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and _52914_ (_08209_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or _52915_ (_08210_, _08209_, _08208_);
  and _52916_ (_08211_, _08210_, _34581_);
  and _52917_ (_08212_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and _52918_ (_08213_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or _52919_ (_08214_, _08213_, _08212_);
  and _52920_ (_08215_, _08214_, _34796_);
  or _52921_ (_08216_, _08215_, _08211_);
  or _52922_ (_08217_, _08216_, _34790_);
  and _52923_ (_08218_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and _52924_ (_08219_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or _52925_ (_08220_, _08219_, _08218_);
  and _52926_ (_08221_, _08220_, _34581_);
  and _52927_ (_08222_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and _52928_ (_08223_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or _52929_ (_08224_, _08223_, _08222_);
  and _52930_ (_08225_, _08224_, _34796_);
  or _52931_ (_08226_, _08225_, _08221_);
  or _52932_ (_08227_, _08226_, _34772_);
  and _52933_ (_08228_, _08227_, _34803_);
  and _52934_ (_08229_, _08228_, _08217_);
  or _52935_ (_08230_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or _52936_ (_08231_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and _52937_ (_08232_, _08231_, _08230_);
  and _52938_ (_08233_, _08232_, _34581_);
  or _52939_ (_08234_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or _52940_ (_08235_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and _52941_ (_08236_, _08235_, _08234_);
  and _52942_ (_08237_, _08236_, _34796_);
  or _52943_ (_08238_, _08237_, _08233_);
  or _52944_ (_08239_, _08238_, _34790_);
  or _52945_ (_08240_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or _52946_ (_08241_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and _52947_ (_08242_, _08241_, _08240_);
  and _52948_ (_08243_, _08242_, _34581_);
  or _52949_ (_08244_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or _52950_ (_08245_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and _52951_ (_08246_, _08245_, _08244_);
  and _52952_ (_08247_, _08246_, _34796_);
  or _52953_ (_08248_, _08247_, _08243_);
  or _52954_ (_08249_, _08248_, _34772_);
  and _52955_ (_08250_, _08249_, _34719_);
  and _52956_ (_08251_, _08250_, _08239_);
  or _52957_ (_08252_, _08251_, _08229_);
  and _52958_ (_08253_, _08252_, _34700_);
  and _52959_ (_08254_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and _52960_ (_08255_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or _52961_ (_08256_, _08255_, _08254_);
  and _52962_ (_08257_, _08256_, _34581_);
  and _52963_ (_08258_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and _52964_ (_08259_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or _52965_ (_08260_, _08259_, _08258_);
  and _52966_ (_08261_, _08260_, _34796_);
  or _52967_ (_08262_, _08261_, _08257_);
  or _52968_ (_08263_, _08262_, _34790_);
  and _52969_ (_08264_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and _52970_ (_08265_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or _52971_ (_08266_, _08265_, _08264_);
  and _52972_ (_08267_, _08266_, _34581_);
  and _52973_ (_08268_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and _52974_ (_08269_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or _52975_ (_08270_, _08269_, _08268_);
  and _52976_ (_08271_, _08270_, _34796_);
  or _52977_ (_08272_, _08271_, _08267_);
  or _52978_ (_08273_, _08272_, _34772_);
  and _52979_ (_08274_, _08273_, _34803_);
  and _52980_ (_08275_, _08274_, _08263_);
  or _52981_ (_08276_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or _52982_ (_08277_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and _52983_ (_08278_, _08277_, _34796_);
  and _52984_ (_08279_, _08278_, _08276_);
  or _52985_ (_08280_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or _52986_ (_08281_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and _52987_ (_08282_, _08281_, _34581_);
  and _52988_ (_08283_, _08282_, _08280_);
  or _52989_ (_08284_, _08283_, _08279_);
  or _52990_ (_08285_, _08284_, _34790_);
  or _52991_ (_08286_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or _52992_ (_08287_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and _52993_ (_08288_, _08287_, _34796_);
  and _52994_ (_08289_, _08288_, _08286_);
  or _52995_ (_08290_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or _52996_ (_08291_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and _52997_ (_08292_, _08291_, _34581_);
  and _52998_ (_08293_, _08292_, _08290_);
  or _52999_ (_08294_, _08293_, _08289_);
  or _53000_ (_08295_, _08294_, _34772_);
  and _53001_ (_08296_, _08295_, _34719_);
  and _53002_ (_08297_, _08296_, _08285_);
  or _53003_ (_08298_, _08297_, _08275_);
  and _53004_ (_08299_, _08298_, _34789_);
  or _53005_ (_08300_, _08299_, _08253_);
  and _53006_ (_08301_, _08300_, _34840_);
  and _53007_ (_08302_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and _53008_ (_08303_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or _53009_ (_08304_, _08303_, _08302_);
  and _53010_ (_08305_, _08304_, _34581_);
  and _53011_ (_08306_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and _53012_ (_08307_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or _53013_ (_08308_, _08307_, _08306_);
  and _53014_ (_08309_, _08308_, _34796_);
  or _53015_ (_08310_, _08309_, _08305_);
  and _53016_ (_08311_, _08310_, _34772_);
  and _53017_ (_08312_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and _53018_ (_08313_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or _53019_ (_08314_, _08313_, _08312_);
  and _53020_ (_08315_, _08314_, _34581_);
  and _53021_ (_08316_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and _53022_ (_08317_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or _53023_ (_08318_, _08317_, _08316_);
  and _53024_ (_08319_, _08318_, _34796_);
  or _53025_ (_08320_, _08319_, _08315_);
  and _53026_ (_08321_, _08320_, _34790_);
  or _53027_ (_08322_, _08321_, _08311_);
  and _53028_ (_08323_, _08322_, _34803_);
  or _53029_ (_08324_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or _53030_ (_08325_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and _53031_ (_08326_, _08325_, _34796_);
  and _53032_ (_08327_, _08326_, _08324_);
  or _53033_ (_08328_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or _53034_ (_08329_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and _53035_ (_08330_, _08329_, _34581_);
  and _53036_ (_08331_, _08330_, _08328_);
  or _53037_ (_08332_, _08331_, _08327_);
  and _53038_ (_08333_, _08332_, _34772_);
  or _53039_ (_08334_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or _53040_ (_08335_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and _53041_ (_08336_, _08335_, _34796_);
  and _53042_ (_08337_, _08336_, _08334_);
  or _53043_ (_08338_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or _53044_ (_08339_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and _53045_ (_08340_, _08339_, _34581_);
  and _53046_ (_08341_, _08340_, _08338_);
  or _53047_ (_08342_, _08341_, _08337_);
  and _53048_ (_08343_, _08342_, _34790_);
  or _53049_ (_08344_, _08343_, _08333_);
  and _53050_ (_08345_, _08344_, _34719_);
  or _53051_ (_08346_, _08345_, _08323_);
  and _53052_ (_08347_, _08346_, _34789_);
  and _53053_ (_08348_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and _53054_ (_08349_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or _53055_ (_08350_, _08349_, _08348_);
  and _53056_ (_08351_, _08350_, _34581_);
  and _53057_ (_08352_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and _53058_ (_08353_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or _53059_ (_08354_, _08353_, _08352_);
  and _53060_ (_08355_, _08354_, _34796_);
  or _53061_ (_08356_, _08355_, _08351_);
  and _53062_ (_08357_, _08356_, _34772_);
  and _53063_ (_08358_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and _53064_ (_08359_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or _53065_ (_08360_, _08359_, _08358_);
  and _53066_ (_08361_, _08360_, _34581_);
  and _53067_ (_08362_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and _53068_ (_08363_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or _53069_ (_08364_, _08363_, _08362_);
  and _53070_ (_08365_, _08364_, _34796_);
  or _53071_ (_08366_, _08365_, _08361_);
  and _53072_ (_08367_, _08366_, _34790_);
  or _53073_ (_08368_, _08367_, _08357_);
  and _53074_ (_08369_, _08368_, _34803_);
  or _53075_ (_08370_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or _53076_ (_08371_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and _53077_ (_08372_, _08371_, _08370_);
  and _53078_ (_08373_, _08372_, _34581_);
  or _53079_ (_08374_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or _53080_ (_08375_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and _53081_ (_08376_, _08375_, _08374_);
  and _53082_ (_08377_, _08376_, _34796_);
  or _53083_ (_08378_, _08377_, _08373_);
  and _53084_ (_08379_, _08378_, _34772_);
  or _53085_ (_08380_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or _53086_ (_08381_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and _53087_ (_08382_, _08381_, _08380_);
  and _53088_ (_08383_, _08382_, _34581_);
  or _53089_ (_08384_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or _53090_ (_08385_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and _53091_ (_08386_, _08385_, _08384_);
  and _53092_ (_08387_, _08386_, _34796_);
  or _53093_ (_08388_, _08387_, _08383_);
  and _53094_ (_08389_, _08388_, _34790_);
  or _53095_ (_08390_, _08389_, _08379_);
  and _53096_ (_08391_, _08390_, _34719_);
  or _53097_ (_08392_, _08391_, _08369_);
  and _53098_ (_08393_, _08392_, _34700_);
  or _53099_ (_08394_, _08393_, _08347_);
  and _53100_ (_08395_, _08394_, _34638_);
  or _53101_ (_08396_, _08395_, _08301_);
  or _53102_ (_08397_, _08396_, _34692_);
  and _53103_ (_08398_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and _53104_ (_08399_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or _53105_ (_08400_, _08399_, _08398_);
  and _53106_ (_08401_, _08400_, _34581_);
  and _53107_ (_08402_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and _53108_ (_08403_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or _53109_ (_08404_, _08403_, _08402_);
  and _53110_ (_08405_, _08404_, _34796_);
  or _53111_ (_08406_, _08405_, _08401_);
  or _53112_ (_08407_, _08406_, _34790_);
  and _53113_ (_08408_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and _53114_ (_08409_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or _53115_ (_08410_, _08409_, _08408_);
  and _53116_ (_08411_, _08410_, _34581_);
  and _53117_ (_08412_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and _53118_ (_08413_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or _53119_ (_08414_, _08413_, _08412_);
  and _53120_ (_08415_, _08414_, _34796_);
  or _53121_ (_08416_, _08415_, _08411_);
  or _53122_ (_08417_, _08416_, _34772_);
  and _53123_ (_08418_, _08417_, _34803_);
  and _53124_ (_08419_, _08418_, _08407_);
  or _53125_ (_08420_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or _53126_ (_08421_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and _53127_ (_08422_, _08421_, _34796_);
  and _53128_ (_08423_, _08422_, _08420_);
  or _53129_ (_08424_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or _53130_ (_08425_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and _53131_ (_08426_, _08425_, _34581_);
  and _53132_ (_08427_, _08426_, _08424_);
  or _53133_ (_08428_, _08427_, _08423_);
  or _53134_ (_08429_, _08428_, _34790_);
  or _53135_ (_08430_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or _53136_ (_08431_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and _53137_ (_08432_, _08431_, _34796_);
  and _53138_ (_08433_, _08432_, _08430_);
  or _53139_ (_08434_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or _53140_ (_08435_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and _53141_ (_08436_, _08435_, _34581_);
  and _53142_ (_08437_, _08436_, _08434_);
  or _53143_ (_08438_, _08437_, _08433_);
  or _53144_ (_08439_, _08438_, _34772_);
  and _53145_ (_08440_, _08439_, _34719_);
  and _53146_ (_08441_, _08440_, _08429_);
  or _53147_ (_08442_, _08441_, _08419_);
  and _53148_ (_08443_, _08442_, _34789_);
  and _53149_ (_08444_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and _53150_ (_08445_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or _53151_ (_08446_, _08445_, _08444_);
  and _53152_ (_08447_, _08446_, _34581_);
  and _53153_ (_08448_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and _53154_ (_08449_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or _53155_ (_08450_, _08449_, _08448_);
  and _53156_ (_08451_, _08450_, _34796_);
  or _53157_ (_08452_, _08451_, _08447_);
  or _53158_ (_08453_, _08452_, _34790_);
  and _53159_ (_08454_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and _53160_ (_08455_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or _53161_ (_08456_, _08455_, _08454_);
  and _53162_ (_08457_, _08456_, _34581_);
  and _53163_ (_08458_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and _53164_ (_08459_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or _53165_ (_08460_, _08459_, _08458_);
  and _53166_ (_08461_, _08460_, _34796_);
  or _53167_ (_08462_, _08461_, _08457_);
  or _53168_ (_08463_, _08462_, _34772_);
  and _53169_ (_08464_, _08463_, _34803_);
  and _53170_ (_08465_, _08464_, _08453_);
  or _53171_ (_08466_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or _53172_ (_08467_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and _53173_ (_08468_, _08467_, _08466_);
  and _53174_ (_08469_, _08468_, _34581_);
  or _53175_ (_08470_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or _53176_ (_08471_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and _53177_ (_08472_, _08471_, _08470_);
  and _53178_ (_08473_, _08472_, _34796_);
  or _53179_ (_08474_, _08473_, _08469_);
  or _53180_ (_08475_, _08474_, _34790_);
  or _53181_ (_08476_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or _53182_ (_08477_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and _53183_ (_08478_, _08477_, _08476_);
  and _53184_ (_08479_, _08478_, _34581_);
  or _53185_ (_08480_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or _53186_ (_08481_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and _53187_ (_08482_, _08481_, _08480_);
  and _53188_ (_08483_, _08482_, _34796_);
  or _53189_ (_08484_, _08483_, _08479_);
  or _53190_ (_08485_, _08484_, _34772_);
  and _53191_ (_08486_, _08485_, _34719_);
  and _53192_ (_08487_, _08486_, _08475_);
  or _53193_ (_08488_, _08487_, _08465_);
  and _53194_ (_08489_, _08488_, _34700_);
  or _53195_ (_08490_, _08489_, _08443_);
  and _53196_ (_08491_, _08490_, _34840_);
  or _53197_ (_08492_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or _53198_ (_08493_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and _53199_ (_08494_, _08493_, _08492_);
  and _53200_ (_08495_, _08494_, _34581_);
  or _53201_ (_08496_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or _53202_ (_08497_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and _53203_ (_08498_, _08497_, _08496_);
  and _53204_ (_08499_, _08498_, _34796_);
  or _53205_ (_08500_, _08499_, _08495_);
  and _53206_ (_08501_, _08500_, _34790_);
  or _53207_ (_08502_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or _53208_ (_08503_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and _53209_ (_08504_, _08503_, _08502_);
  and _53210_ (_08505_, _08504_, _34581_);
  or _53211_ (_08506_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or _53212_ (_08507_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and _53213_ (_08508_, _08507_, _08506_);
  and _53214_ (_08509_, _08508_, _34796_);
  or _53215_ (_08510_, _08509_, _08505_);
  and _53216_ (_08511_, _08510_, _34772_);
  or _53217_ (_08512_, _08511_, _08501_);
  and _53218_ (_08513_, _08512_, _34719_);
  and _53219_ (_08514_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and _53220_ (_08515_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or _53221_ (_08516_, _08515_, _08514_);
  and _53222_ (_08517_, _08516_, _34581_);
  and _53223_ (_08518_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and _53224_ (_08519_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or _53225_ (_08520_, _08519_, _08518_);
  and _53226_ (_08521_, _08520_, _34796_);
  or _53227_ (_08522_, _08521_, _08517_);
  and _53228_ (_08523_, _08522_, _34790_);
  and _53229_ (_08524_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and _53230_ (_08525_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or _53231_ (_08526_, _08525_, _08524_);
  and _53232_ (_08527_, _08526_, _34581_);
  and _53233_ (_08528_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and _53234_ (_08529_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or _53235_ (_08530_, _08529_, _08528_);
  and _53236_ (_08531_, _08530_, _34796_);
  or _53237_ (_08532_, _08531_, _08527_);
  and _53238_ (_08533_, _08532_, _34772_);
  or _53239_ (_08534_, _08533_, _08523_);
  and _53240_ (_08535_, _08534_, _34803_);
  or _53241_ (_08536_, _08535_, _08513_);
  and _53242_ (_08537_, _08536_, _34700_);
  or _53243_ (_08538_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or _53244_ (_08539_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and _53245_ (_08540_, _08539_, _34796_);
  and _53246_ (_08541_, _08540_, _08538_);
  or _53247_ (_08542_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or _53248_ (_08543_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and _53249_ (_08544_, _08543_, _34581_);
  and _53250_ (_08545_, _08544_, _08542_);
  or _53251_ (_08546_, _08545_, _08541_);
  and _53252_ (_08547_, _08546_, _34790_);
  or _53253_ (_08548_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or _53254_ (_08549_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and _53255_ (_08550_, _08549_, _34796_);
  and _53256_ (_08551_, _08550_, _08548_);
  or _53257_ (_08552_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or _53258_ (_08553_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and _53259_ (_08554_, _08553_, _34581_);
  and _53260_ (_08555_, _08554_, _08552_);
  or _53261_ (_08556_, _08555_, _08551_);
  and _53262_ (_08557_, _08556_, _34772_);
  or _53263_ (_08558_, _08557_, _08547_);
  and _53264_ (_08559_, _08558_, _34719_);
  and _53265_ (_08560_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and _53266_ (_08561_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or _53267_ (_08562_, _08561_, _08560_);
  and _53268_ (_08563_, _08562_, _34581_);
  and _53269_ (_08564_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and _53270_ (_08565_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or _53271_ (_08566_, _08565_, _08564_);
  and _53272_ (_08567_, _08566_, _34796_);
  or _53273_ (_08568_, _08567_, _08563_);
  and _53274_ (_08569_, _08568_, _34790_);
  and _53275_ (_08570_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and _53276_ (_08571_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or _53277_ (_08572_, _08571_, _08570_);
  and _53278_ (_08573_, _08572_, _34581_);
  and _53279_ (_08574_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and _53280_ (_08575_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or _53281_ (_08576_, _08575_, _08574_);
  and _53282_ (_08577_, _08576_, _34796_);
  or _53283_ (_08578_, _08577_, _08573_);
  and _53284_ (_08579_, _08578_, _34772_);
  or _53285_ (_08580_, _08579_, _08569_);
  and _53286_ (_08581_, _08580_, _34803_);
  or _53287_ (_08582_, _08581_, _08559_);
  and _53288_ (_08583_, _08582_, _34789_);
  or _53289_ (_08584_, _08583_, _08537_);
  and _53290_ (_08585_, _08584_, _34638_);
  or _53291_ (_08586_, _08585_, _08491_);
  or _53292_ (_08587_, _08586_, _34985_);
  and _53293_ (_08588_, _08587_, _08397_);
  or _53294_ (_08589_, _08588_, _35178_);
  and _53295_ (_08590_, _08589_, _08207_);
  or _53296_ (_08591_, _08590_, _34788_);
  or _53297_ (_08592_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and _53298_ (_08593_, _08592_, _38997_);
  and _53299_ (_38984_[3], _08593_, _08591_);
  and _53300_ (_08594_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and _53301_ (_08595_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or _53302_ (_08596_, _08595_, _08594_);
  and _53303_ (_08597_, _08596_, _34581_);
  and _53304_ (_08598_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and _53305_ (_08599_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or _53306_ (_08600_, _08599_, _08598_);
  and _53307_ (_08601_, _08600_, _34796_);
  or _53308_ (_08602_, _08601_, _08597_);
  or _53309_ (_08603_, _08602_, _34790_);
  and _53310_ (_08604_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and _53311_ (_08605_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or _53312_ (_08606_, _08605_, _08604_);
  and _53313_ (_08607_, _08606_, _34581_);
  and _53314_ (_08608_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  and _53315_ (_08609_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or _53316_ (_08610_, _08609_, _08608_);
  and _53317_ (_08611_, _08610_, _34796_);
  or _53318_ (_08612_, _08611_, _08607_);
  or _53319_ (_08613_, _08612_, _34772_);
  and _53320_ (_08614_, _08613_, _34803_);
  and _53321_ (_08615_, _08614_, _08603_);
  or _53322_ (_08616_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or _53323_ (_08617_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and _53324_ (_08618_, _08617_, _08616_);
  and _53325_ (_08619_, _08618_, _34581_);
  or _53326_ (_08620_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or _53327_ (_08621_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  and _53328_ (_08622_, _08621_, _08620_);
  and _53329_ (_08623_, _08622_, _34796_);
  or _53330_ (_08624_, _08623_, _08619_);
  or _53331_ (_08625_, _08624_, _34790_);
  or _53332_ (_08626_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or _53333_ (_08627_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and _53334_ (_08628_, _08627_, _08626_);
  and _53335_ (_08629_, _08628_, _34581_);
  or _53336_ (_08630_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or _53337_ (_08631_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and _53338_ (_08632_, _08631_, _08630_);
  and _53339_ (_08633_, _08632_, _34796_);
  or _53340_ (_08634_, _08633_, _08629_);
  or _53341_ (_08635_, _08634_, _34772_);
  and _53342_ (_08636_, _08635_, _34719_);
  and _53343_ (_08637_, _08636_, _08625_);
  or _53344_ (_08638_, _08637_, _08615_);
  or _53345_ (_08639_, _08638_, _34789_);
  and _53346_ (_08640_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and _53347_ (_08641_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or _53348_ (_08642_, _08641_, _08640_);
  and _53349_ (_08643_, _08642_, _34581_);
  and _53350_ (_08644_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  and _53351_ (_08645_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or _53352_ (_08646_, _08645_, _08644_);
  and _53353_ (_08647_, _08646_, _34796_);
  or _53354_ (_08648_, _08647_, _08643_);
  or _53355_ (_08649_, _08648_, _34790_);
  and _53356_ (_08650_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and _53357_ (_08651_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or _53358_ (_08652_, _08651_, _08650_);
  and _53359_ (_08653_, _08652_, _34581_);
  and _53360_ (_08654_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and _53361_ (_08655_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or _53362_ (_08656_, _08655_, _08654_);
  and _53363_ (_08657_, _08656_, _34796_);
  or _53364_ (_08658_, _08657_, _08653_);
  or _53365_ (_08659_, _08658_, _34772_);
  and _53366_ (_08660_, _08659_, _34803_);
  and _53367_ (_08661_, _08660_, _08649_);
  or _53368_ (_08662_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or _53369_ (_08663_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and _53370_ (_08664_, _08663_, _34796_);
  and _53371_ (_08665_, _08664_, _08662_);
  or _53372_ (_08666_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or _53373_ (_08667_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and _53374_ (_08668_, _08667_, _34581_);
  and _53375_ (_08669_, _08668_, _08666_);
  or _53376_ (_08670_, _08669_, _08665_);
  or _53377_ (_08671_, _08670_, _34790_);
  or _53378_ (_08672_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or _53379_ (_08673_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and _53380_ (_08674_, _08673_, _34796_);
  and _53381_ (_08675_, _08674_, _08672_);
  or _53382_ (_08676_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or _53383_ (_08677_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  and _53384_ (_08678_, _08677_, _34581_);
  and _53385_ (_08679_, _08678_, _08676_);
  or _53386_ (_08680_, _08679_, _08675_);
  or _53387_ (_08681_, _08680_, _34772_);
  and _53388_ (_08682_, _08681_, _34719_);
  and _53389_ (_08683_, _08682_, _08671_);
  or _53390_ (_08684_, _08683_, _08661_);
  or _53391_ (_08685_, _08684_, _34700_);
  and _53392_ (_08686_, _08685_, _34840_);
  and _53393_ (_08687_, _08686_, _08639_);
  and _53394_ (_08688_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and _53395_ (_08689_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or _53396_ (_08690_, _08689_, _08688_);
  and _53397_ (_08691_, _08690_, _34581_);
  and _53398_ (_08692_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and _53399_ (_08693_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or _53400_ (_08694_, _08693_, _08692_);
  and _53401_ (_08695_, _08694_, _34796_);
  or _53402_ (_08696_, _08695_, _08691_);
  and _53403_ (_08697_, _08696_, _34772_);
  and _53404_ (_08698_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and _53405_ (_08699_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _53406_ (_08700_, _08699_, _08698_);
  and _53407_ (_08701_, _08700_, _34581_);
  and _53408_ (_08702_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and _53409_ (_08703_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or _53410_ (_08704_, _08703_, _08702_);
  and _53411_ (_08705_, _08704_, _34796_);
  or _53412_ (_08706_, _08705_, _08701_);
  and _53413_ (_08707_, _08706_, _34790_);
  or _53414_ (_08708_, _08707_, _34719_);
  or _53415_ (_08709_, _08708_, _08697_);
  or _53416_ (_08710_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _53417_ (_08711_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and _53418_ (_08712_, _08711_, _34796_);
  and _53419_ (_08713_, _08712_, _08710_);
  or _53420_ (_08714_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or _53421_ (_08715_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and _53422_ (_08716_, _08715_, _34581_);
  and _53423_ (_08717_, _08716_, _08714_);
  or _53424_ (_08718_, _08717_, _08713_);
  and _53425_ (_08719_, _08718_, _34772_);
  or _53426_ (_08720_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _53427_ (_08721_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and _53428_ (_08722_, _08721_, _34796_);
  and _53429_ (_08723_, _08722_, _08720_);
  or _53430_ (_08724_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or _53431_ (_08725_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and _53432_ (_08726_, _08725_, _34581_);
  and _53433_ (_08727_, _08726_, _08724_);
  or _53434_ (_08728_, _08727_, _08723_);
  and _53435_ (_08729_, _08728_, _34790_);
  or _53436_ (_08730_, _08729_, _34803_);
  or _53437_ (_08731_, _08730_, _08719_);
  and _53438_ (_08732_, _08731_, _08709_);
  or _53439_ (_08733_, _08732_, _34700_);
  and _53440_ (_08734_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and _53441_ (_08735_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or _53442_ (_08736_, _08735_, _08734_);
  and _53443_ (_08737_, _08736_, _34581_);
  and _53444_ (_08738_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and _53445_ (_08739_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or _53446_ (_08740_, _08739_, _08738_);
  and _53447_ (_08741_, _08740_, _34796_);
  or _53448_ (_08742_, _08741_, _08737_);
  and _53449_ (_08743_, _08742_, _34772_);
  and _53450_ (_08744_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and _53451_ (_08745_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or _53452_ (_08746_, _08745_, _08744_);
  and _53453_ (_08747_, _08746_, _34581_);
  and _53454_ (_08748_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and _53455_ (_08749_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or _53456_ (_08750_, _08749_, _08748_);
  and _53457_ (_08751_, _08750_, _34796_);
  or _53458_ (_08752_, _08751_, _08747_);
  and _53459_ (_08753_, _08752_, _34790_);
  or _53460_ (_08754_, _08753_, _34719_);
  or _53461_ (_08755_, _08754_, _08743_);
  or _53462_ (_08756_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or _53463_ (_08757_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and _53464_ (_08758_, _08757_, _08756_);
  and _53465_ (_08759_, _08758_, _34581_);
  or _53466_ (_08760_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or _53467_ (_08761_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and _53468_ (_08762_, _08761_, _08760_);
  and _53469_ (_08763_, _08762_, _34796_);
  or _53470_ (_08764_, _08763_, _08759_);
  and _53471_ (_08765_, _08764_, _34772_);
  or _53472_ (_08766_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or _53473_ (_08767_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and _53474_ (_08768_, _08767_, _08766_);
  and _53475_ (_08769_, _08768_, _34581_);
  or _53476_ (_08770_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or _53477_ (_08771_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and _53478_ (_08772_, _08771_, _08770_);
  and _53479_ (_08773_, _08772_, _34796_);
  or _53480_ (_08774_, _08773_, _08769_);
  and _53481_ (_08775_, _08774_, _34790_);
  or _53482_ (_08776_, _08775_, _34803_);
  or _53483_ (_08777_, _08776_, _08765_);
  and _53484_ (_08778_, _08777_, _08755_);
  or _53485_ (_08779_, _08778_, _34789_);
  and _53486_ (_08780_, _08779_, _34638_);
  and _53487_ (_08781_, _08780_, _08733_);
  or _53488_ (_08782_, _08781_, _08687_);
  or _53489_ (_08783_, _08782_, _34692_);
  and _53490_ (_08784_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  and _53491_ (_08785_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or _53492_ (_08786_, _08785_, _08784_);
  and _53493_ (_08787_, _08786_, _34581_);
  and _53494_ (_08788_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  and _53495_ (_08789_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  or _53496_ (_08790_, _08789_, _08788_);
  and _53497_ (_08791_, _08790_, _34796_);
  or _53498_ (_08792_, _08791_, _08787_);
  and _53499_ (_08793_, _08792_, _34772_);
  and _53500_ (_08794_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  and _53501_ (_08795_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  or _53502_ (_08796_, _08795_, _08794_);
  and _53503_ (_08797_, _08796_, _34581_);
  and _53504_ (_08798_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  and _53505_ (_08799_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or _53506_ (_08800_, _08799_, _08798_);
  and _53507_ (_08801_, _08800_, _34796_);
  or _53508_ (_08802_, _08801_, _08797_);
  and _53509_ (_08803_, _08802_, _34790_);
  or _53510_ (_08804_, _08803_, _34719_);
  or _53511_ (_08805_, _08804_, _08793_);
  or _53512_ (_08806_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or _53513_ (_08807_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  and _53514_ (_08808_, _08807_, _08806_);
  and _53515_ (_08809_, _08808_, _34581_);
  or _53516_ (_08810_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or _53517_ (_08811_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  and _53518_ (_08812_, _08811_, _08810_);
  and _53519_ (_08813_, _08812_, _34796_);
  or _53520_ (_08814_, _08813_, _08809_);
  and _53521_ (_08815_, _08814_, _34772_);
  or _53522_ (_08816_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  or _53523_ (_08817_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  and _53524_ (_08818_, _08817_, _08816_);
  and _53525_ (_08819_, _08818_, _34581_);
  or _53526_ (_08820_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or _53527_ (_08821_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  and _53528_ (_08822_, _08821_, _08820_);
  and _53529_ (_08823_, _08822_, _34796_);
  or _53530_ (_08824_, _08823_, _08819_);
  and _53531_ (_08825_, _08824_, _34790_);
  or _53532_ (_08826_, _08825_, _34803_);
  or _53533_ (_08827_, _08826_, _08815_);
  and _53534_ (_08828_, _08827_, _08805_);
  or _53535_ (_08829_, _08828_, _34700_);
  and _53536_ (_08830_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and _53537_ (_08831_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or _53538_ (_08832_, _08831_, _08830_);
  and _53539_ (_08833_, _08832_, _34581_);
  and _53540_ (_08834_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and _53541_ (_08835_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or _53542_ (_08836_, _08835_, _08834_);
  and _53543_ (_08837_, _08836_, _34796_);
  or _53544_ (_08838_, _08837_, _08833_);
  and _53545_ (_08839_, _08838_, _34772_);
  and _53546_ (_08840_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and _53547_ (_08841_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or _53548_ (_08842_, _08841_, _08840_);
  and _53549_ (_08843_, _08842_, _34581_);
  and _53550_ (_08844_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and _53551_ (_08845_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or _53552_ (_08846_, _08845_, _08844_);
  and _53553_ (_08847_, _08846_, _34796_);
  or _53554_ (_08848_, _08847_, _08843_);
  and _53555_ (_08849_, _08848_, _34790_);
  or _53556_ (_08850_, _08849_, _34719_);
  or _53557_ (_08851_, _08850_, _08839_);
  or _53558_ (_08852_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or _53559_ (_08853_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and _53560_ (_08854_, _08853_, _08852_);
  and _53561_ (_08855_, _08854_, _34581_);
  or _53562_ (_08856_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or _53563_ (_08857_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  and _53564_ (_08858_, _08857_, _08856_);
  and _53565_ (_08859_, _08858_, _34796_);
  or _53566_ (_08860_, _08859_, _08855_);
  and _53567_ (_08861_, _08860_, _34772_);
  or _53568_ (_08862_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or _53569_ (_08863_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  and _53570_ (_08864_, _08863_, _08862_);
  and _53571_ (_08865_, _08864_, _34581_);
  or _53572_ (_08866_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or _53573_ (_08867_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and _53574_ (_08868_, _08867_, _08866_);
  and _53575_ (_08869_, _08868_, _34796_);
  or _53576_ (_08870_, _08869_, _08865_);
  and _53577_ (_08871_, _08870_, _34790_);
  or _53578_ (_08872_, _08871_, _34803_);
  or _53579_ (_08873_, _08872_, _08861_);
  and _53580_ (_08874_, _08873_, _08851_);
  or _53581_ (_08875_, _08874_, _34789_);
  and _53582_ (_08876_, _08875_, _34638_);
  and _53583_ (_08877_, _08876_, _08829_);
  and _53584_ (_08878_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and _53585_ (_08879_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or _53586_ (_08880_, _08879_, _08878_);
  and _53587_ (_08881_, _08880_, _34796_);
  and _53588_ (_08882_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  and _53589_ (_08883_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or _53590_ (_08884_, _08883_, _08882_);
  and _53591_ (_08885_, _08884_, _34581_);
  or _53592_ (_08886_, _08885_, _08881_);
  or _53593_ (_08887_, _08886_, _34790_);
  and _53594_ (_08888_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and _53595_ (_08889_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or _53596_ (_08890_, _08889_, _08888_);
  and _53597_ (_08891_, _08890_, _34796_);
  and _53598_ (_08892_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and _53599_ (_08893_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or _53600_ (_08894_, _08893_, _08892_);
  and _53601_ (_08895_, _08894_, _34581_);
  or _53602_ (_08896_, _08895_, _08891_);
  or _53603_ (_08897_, _08896_, _34772_);
  and _53604_ (_08898_, _08897_, _34803_);
  and _53605_ (_08899_, _08898_, _08887_);
  or _53606_ (_08900_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or _53607_ (_08901_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and _53608_ (_08902_, _08901_, _34581_);
  and _53609_ (_08903_, _08902_, _08900_);
  or _53610_ (_08904_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or _53611_ (_08905_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and _53612_ (_08906_, _08905_, _34796_);
  and _53613_ (_08907_, _08906_, _08904_);
  or _53614_ (_08908_, _08907_, _08903_);
  or _53615_ (_08909_, _08908_, _34790_);
  or _53616_ (_08910_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or _53617_ (_08911_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  and _53618_ (_08912_, _08911_, _34581_);
  and _53619_ (_08913_, _08912_, _08910_);
  or _53620_ (_08914_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or _53621_ (_08915_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and _53622_ (_08916_, _08915_, _34796_);
  and _53623_ (_08917_, _08916_, _08914_);
  or _53624_ (_08918_, _08917_, _08913_);
  or _53625_ (_08919_, _08918_, _34772_);
  and _53626_ (_08920_, _08919_, _34719_);
  and _53627_ (_08921_, _08920_, _08909_);
  or _53628_ (_08922_, _08921_, _08899_);
  and _53629_ (_08923_, _08922_, _34789_);
  and _53630_ (_08924_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and _53631_ (_08925_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or _53632_ (_08926_, _08925_, _34581_);
  or _53633_ (_08927_, _08926_, _08924_);
  and _53634_ (_08928_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and _53635_ (_08929_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or _53636_ (_08930_, _08929_, _34796_);
  or _53637_ (_08931_, _08930_, _08928_);
  and _53638_ (_08932_, _08931_, _08927_);
  or _53639_ (_08933_, _08932_, _34790_);
  and _53640_ (_08934_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and _53641_ (_08935_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or _53642_ (_08936_, _08935_, _34581_);
  or _53643_ (_08937_, _08936_, _08934_);
  and _53644_ (_08938_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and _53645_ (_08939_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or _53646_ (_08940_, _08939_, _34796_);
  or _53647_ (_08941_, _08940_, _08938_);
  and _53648_ (_08942_, _08941_, _08937_);
  or _53649_ (_08943_, _08942_, _34772_);
  and _53650_ (_08944_, _08943_, _34803_);
  and _53651_ (_08945_, _08944_, _08933_);
  or _53652_ (_08946_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or _53653_ (_08947_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and _53654_ (_08948_, _08947_, _08946_);
  or _53655_ (_08949_, _08948_, _34796_);
  or _53656_ (_08950_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or _53657_ (_08951_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and _53658_ (_08952_, _08951_, _08950_);
  or _53659_ (_08953_, _08952_, _34581_);
  and _53660_ (_08954_, _08953_, _08949_);
  or _53661_ (_08955_, _08954_, _34790_);
  or _53662_ (_08956_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or _53663_ (_08957_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and _53664_ (_08958_, _08957_, _08956_);
  or _53665_ (_08959_, _08958_, _34796_);
  or _53666_ (_08960_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or _53667_ (_08961_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and _53668_ (_08962_, _08961_, _08960_);
  or _53669_ (_08963_, _08962_, _34581_);
  and _53670_ (_08964_, _08963_, _08959_);
  or _53671_ (_08965_, _08964_, _34772_);
  and _53672_ (_08966_, _08965_, _34719_);
  and _53673_ (_08967_, _08966_, _08955_);
  or _53674_ (_08968_, _08967_, _08945_);
  and _53675_ (_08969_, _08968_, _34700_);
  or _53676_ (_08970_, _08969_, _08923_);
  and _53677_ (_08971_, _08970_, _34840_);
  or _53678_ (_08972_, _08971_, _08877_);
  or _53679_ (_08973_, _08972_, _34985_);
  and _53680_ (_08974_, _08973_, _08783_);
  or _53681_ (_08975_, _08974_, _34346_);
  and _53682_ (_08976_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and _53683_ (_08977_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or _53684_ (_08978_, _08977_, _08976_);
  and _53685_ (_08979_, _08978_, _34581_);
  and _53686_ (_08980_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and _53687_ (_08981_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or _53688_ (_08982_, _08981_, _08980_);
  and _53689_ (_08983_, _08982_, _34796_);
  or _53690_ (_08984_, _08983_, _08979_);
  or _53691_ (_08985_, _08984_, _34790_);
  and _53692_ (_08986_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and _53693_ (_08987_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or _53694_ (_08988_, _08987_, _08986_);
  and _53695_ (_08989_, _08988_, _34581_);
  and _53696_ (_08990_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and _53697_ (_08991_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or _53698_ (_08992_, _08991_, _08990_);
  and _53699_ (_08993_, _08992_, _34796_);
  or _53700_ (_08994_, _08993_, _08989_);
  or _53701_ (_08995_, _08994_, _34772_);
  and _53702_ (_08996_, _08995_, _34803_);
  and _53703_ (_08997_, _08996_, _08985_);
  or _53704_ (_08998_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or _53705_ (_08999_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and _53706_ (_09000_, _08999_, _08998_);
  and _53707_ (_09001_, _09000_, _34581_);
  or _53708_ (_09002_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or _53709_ (_09003_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and _53710_ (_09004_, _09003_, _09002_);
  and _53711_ (_09005_, _09004_, _34796_);
  or _53712_ (_09006_, _09005_, _09001_);
  or _53713_ (_09007_, _09006_, _34790_);
  or _53714_ (_09008_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or _53715_ (_09009_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and _53716_ (_09010_, _09009_, _09008_);
  and _53717_ (_09011_, _09010_, _34581_);
  or _53718_ (_09012_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or _53719_ (_09013_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and _53720_ (_09014_, _09013_, _09012_);
  and _53721_ (_09015_, _09014_, _34796_);
  or _53722_ (_09016_, _09015_, _09011_);
  or _53723_ (_09017_, _09016_, _34772_);
  and _53724_ (_09018_, _09017_, _34719_);
  and _53725_ (_09019_, _09018_, _09007_);
  or _53726_ (_09020_, _09019_, _08997_);
  and _53727_ (_09021_, _09020_, _34700_);
  and _53728_ (_09022_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and _53729_ (_09023_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or _53730_ (_09024_, _09023_, _09022_);
  and _53731_ (_09025_, _09024_, _34581_);
  and _53732_ (_09026_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and _53733_ (_09027_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or _53734_ (_09028_, _09027_, _09026_);
  and _53735_ (_09029_, _09028_, _34796_);
  or _53736_ (_09030_, _09029_, _09025_);
  or _53737_ (_09031_, _09030_, _34790_);
  and _53738_ (_09032_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and _53739_ (_09033_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or _53740_ (_09034_, _09033_, _09032_);
  and _53741_ (_09035_, _09034_, _34581_);
  and _53742_ (_09036_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and _53743_ (_09037_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or _53744_ (_09038_, _09037_, _09036_);
  and _53745_ (_09039_, _09038_, _34796_);
  or _53746_ (_09040_, _09039_, _09035_);
  or _53747_ (_09041_, _09040_, _34772_);
  and _53748_ (_09042_, _09041_, _34803_);
  and _53749_ (_09043_, _09042_, _09031_);
  or _53750_ (_09044_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or _53751_ (_09045_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and _53752_ (_09046_, _09045_, _34796_);
  and _53753_ (_09047_, _09046_, _09044_);
  or _53754_ (_09048_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or _53755_ (_09049_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and _53756_ (_09050_, _09049_, _34581_);
  and _53757_ (_09051_, _09050_, _09048_);
  or _53758_ (_09052_, _09051_, _09047_);
  or _53759_ (_09053_, _09052_, _34790_);
  or _53760_ (_09054_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or _53761_ (_09055_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and _53762_ (_09056_, _09055_, _34796_);
  and _53763_ (_09057_, _09056_, _09054_);
  or _53764_ (_09058_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or _53765_ (_09059_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and _53766_ (_09060_, _09059_, _34581_);
  and _53767_ (_09061_, _09060_, _09058_);
  or _53768_ (_09062_, _09061_, _09057_);
  or _53769_ (_09063_, _09062_, _34772_);
  and _53770_ (_09064_, _09063_, _34719_);
  and _53771_ (_09065_, _09064_, _09053_);
  or _53772_ (_09066_, _09065_, _09043_);
  and _53773_ (_09067_, _09066_, _34789_);
  or _53774_ (_09068_, _09067_, _09021_);
  and _53775_ (_09069_, _09068_, _34840_);
  and _53776_ (_09070_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and _53777_ (_09071_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or _53778_ (_09072_, _09071_, _09070_);
  and _53779_ (_09073_, _09072_, _34581_);
  and _53780_ (_09074_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and _53781_ (_09075_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or _53782_ (_09076_, _09075_, _09074_);
  and _53783_ (_09077_, _09076_, _34796_);
  or _53784_ (_09078_, _09077_, _09073_);
  and _53785_ (_09079_, _09078_, _34772_);
  and _53786_ (_09080_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and _53787_ (_09081_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or _53788_ (_09082_, _09081_, _09080_);
  and _53789_ (_09083_, _09082_, _34581_);
  and _53790_ (_09084_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and _53791_ (_09085_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or _53792_ (_09086_, _09085_, _09084_);
  and _53793_ (_09087_, _09086_, _34796_);
  or _53794_ (_09088_, _09087_, _09083_);
  and _53795_ (_09089_, _09088_, _34790_);
  or _53796_ (_09090_, _09089_, _09079_);
  and _53797_ (_09091_, _09090_, _34803_);
  or _53798_ (_09092_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or _53799_ (_09093_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and _53800_ (_09094_, _09093_, _34796_);
  and _53801_ (_09095_, _09094_, _09092_);
  or _53802_ (_09096_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or _53803_ (_09097_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and _53804_ (_09098_, _09097_, _34581_);
  and _53805_ (_09099_, _09098_, _09096_);
  or _53806_ (_09100_, _09099_, _09095_);
  and _53807_ (_09101_, _09100_, _34772_);
  or _53808_ (_09102_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or _53809_ (_09103_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and _53810_ (_09104_, _09103_, _34796_);
  and _53811_ (_09105_, _09104_, _09102_);
  or _53812_ (_09106_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or _53813_ (_09107_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and _53814_ (_09108_, _09107_, _34581_);
  and _53815_ (_09109_, _09108_, _09106_);
  or _53816_ (_09110_, _09109_, _09105_);
  and _53817_ (_09111_, _09110_, _34790_);
  or _53818_ (_09112_, _09111_, _09101_);
  and _53819_ (_09113_, _09112_, _34719_);
  or _53820_ (_09114_, _09113_, _09091_);
  and _53821_ (_09115_, _09114_, _34789_);
  and _53822_ (_09116_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and _53823_ (_09117_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or _53824_ (_09118_, _09117_, _09116_);
  and _53825_ (_09119_, _09118_, _34581_);
  and _53826_ (_09120_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and _53827_ (_09121_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or _53828_ (_09122_, _09121_, _09120_);
  and _53829_ (_09123_, _09122_, _34796_);
  or _53830_ (_09124_, _09123_, _09119_);
  and _53831_ (_09125_, _09124_, _34772_);
  and _53832_ (_09126_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and _53833_ (_09127_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or _53834_ (_09128_, _09127_, _09126_);
  and _53835_ (_09129_, _09128_, _34581_);
  and _53836_ (_09130_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and _53837_ (_09131_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or _53838_ (_09132_, _09131_, _09130_);
  and _53839_ (_09133_, _09132_, _34796_);
  or _53840_ (_09134_, _09133_, _09129_);
  and _53841_ (_09135_, _09134_, _34790_);
  or _53842_ (_09136_, _09135_, _09125_);
  and _53843_ (_09137_, _09136_, _34803_);
  or _53844_ (_09138_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or _53845_ (_09139_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and _53846_ (_09140_, _09139_, _09138_);
  and _53847_ (_09141_, _09140_, _34581_);
  or _53848_ (_09142_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or _53849_ (_09143_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and _53850_ (_09144_, _09143_, _09142_);
  and _53851_ (_09145_, _09144_, _34796_);
  or _53852_ (_09146_, _09145_, _09141_);
  and _53853_ (_09147_, _09146_, _34772_);
  or _53854_ (_09148_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or _53855_ (_09149_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and _53856_ (_09150_, _09149_, _09148_);
  and _53857_ (_09151_, _09150_, _34581_);
  or _53858_ (_09152_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or _53859_ (_09153_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and _53860_ (_09154_, _09153_, _09152_);
  and _53861_ (_09155_, _09154_, _34796_);
  or _53862_ (_09156_, _09155_, _09151_);
  and _53863_ (_09157_, _09156_, _34790_);
  or _53864_ (_09158_, _09157_, _09147_);
  and _53865_ (_09159_, _09158_, _34719_);
  or _53866_ (_09160_, _09159_, _09137_);
  and _53867_ (_09161_, _09160_, _34700_);
  or _53868_ (_09162_, _09161_, _09115_);
  and _53869_ (_09163_, _09162_, _34638_);
  or _53870_ (_09164_, _09163_, _09069_);
  or _53871_ (_09165_, _09164_, _34692_);
  and _53872_ (_09166_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and _53873_ (_09167_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or _53874_ (_09168_, _09167_, _09166_);
  and _53875_ (_09169_, _09168_, _34581_);
  and _53876_ (_09170_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and _53877_ (_09171_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or _53878_ (_09172_, _09171_, _09170_);
  and _53879_ (_09173_, _09172_, _34796_);
  or _53880_ (_09174_, _09173_, _09169_);
  or _53881_ (_09175_, _09174_, _34790_);
  and _53882_ (_09176_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and _53883_ (_09177_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or _53884_ (_09178_, _09177_, _09176_);
  and _53885_ (_09179_, _09178_, _34581_);
  and _53886_ (_09180_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and _53887_ (_09181_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or _53888_ (_09182_, _09181_, _09180_);
  and _53889_ (_09183_, _09182_, _34796_);
  or _53890_ (_09184_, _09183_, _09179_);
  or _53891_ (_09185_, _09184_, _34772_);
  and _53892_ (_09186_, _09185_, _34803_);
  and _53893_ (_09187_, _09186_, _09175_);
  or _53894_ (_09188_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or _53895_ (_09189_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and _53896_ (_09190_, _09189_, _34796_);
  and _53897_ (_09191_, _09190_, _09188_);
  or _53898_ (_09192_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or _53899_ (_09193_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and _53900_ (_09194_, _09193_, _34581_);
  and _53901_ (_09195_, _09194_, _09192_);
  or _53902_ (_09196_, _09195_, _09191_);
  or _53903_ (_09197_, _09196_, _34790_);
  or _53904_ (_09198_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or _53905_ (_09199_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and _53906_ (_09200_, _09199_, _34796_);
  and _53907_ (_09201_, _09200_, _09198_);
  or _53908_ (_09202_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or _53909_ (_09203_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and _53910_ (_09204_, _09203_, _34581_);
  and _53911_ (_09205_, _09204_, _09202_);
  or _53912_ (_09206_, _09205_, _09201_);
  or _53913_ (_09207_, _09206_, _34772_);
  and _53914_ (_09208_, _09207_, _34719_);
  and _53915_ (_09209_, _09208_, _09197_);
  or _53916_ (_09210_, _09209_, _09187_);
  and _53917_ (_09211_, _09210_, _34789_);
  and _53918_ (_09212_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and _53919_ (_09213_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or _53920_ (_09214_, _09213_, _09212_);
  and _53921_ (_09215_, _09214_, _34581_);
  and _53922_ (_09216_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and _53923_ (_09217_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or _53924_ (_09218_, _09217_, _09216_);
  and _53925_ (_09219_, _09218_, _34796_);
  or _53926_ (_09220_, _09219_, _09215_);
  or _53927_ (_09221_, _09220_, _34790_);
  and _53928_ (_09222_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and _53929_ (_09223_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or _53930_ (_09224_, _09223_, _09222_);
  and _53931_ (_09225_, _09224_, _34581_);
  and _53932_ (_09226_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and _53933_ (_09227_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or _53934_ (_09228_, _09227_, _09226_);
  and _53935_ (_09229_, _09228_, _34796_);
  or _53936_ (_09230_, _09229_, _09225_);
  or _53937_ (_09231_, _09230_, _34772_);
  and _53938_ (_09232_, _09231_, _34803_);
  and _53939_ (_09233_, _09232_, _09221_);
  or _53940_ (_09234_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or _53941_ (_09235_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and _53942_ (_09236_, _09235_, _09234_);
  and _53943_ (_09237_, _09236_, _34581_);
  or _53944_ (_09238_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or _53945_ (_09239_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and _53946_ (_09240_, _09239_, _09238_);
  and _53947_ (_09241_, _09240_, _34796_);
  or _53948_ (_09242_, _09241_, _09237_);
  or _53949_ (_09243_, _09242_, _34790_);
  or _53950_ (_09244_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or _53951_ (_09245_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and _53952_ (_09246_, _09245_, _09244_);
  and _53953_ (_09247_, _09246_, _34581_);
  or _53954_ (_09248_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or _53955_ (_09249_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and _53956_ (_09250_, _09249_, _09248_);
  and _53957_ (_09251_, _09250_, _34796_);
  or _53958_ (_09252_, _09251_, _09247_);
  or _53959_ (_09253_, _09252_, _34772_);
  and _53960_ (_09254_, _09253_, _34719_);
  and _53961_ (_09255_, _09254_, _09243_);
  or _53962_ (_09256_, _09255_, _09233_);
  and _53963_ (_09257_, _09256_, _34700_);
  or _53964_ (_09258_, _09257_, _09211_);
  and _53965_ (_09259_, _09258_, _34840_);
  or _53966_ (_09260_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or _53967_ (_09261_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and _53968_ (_09262_, _09261_, _09260_);
  and _53969_ (_09263_, _09262_, _34581_);
  or _53970_ (_09264_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or _53971_ (_09265_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and _53972_ (_09266_, _09265_, _09264_);
  and _53973_ (_09267_, _09266_, _34796_);
  or _53974_ (_09268_, _09267_, _09263_);
  and _53975_ (_09269_, _09268_, _34790_);
  or _53976_ (_09270_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or _53977_ (_09271_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and _53978_ (_09272_, _09271_, _09270_);
  and _53979_ (_09273_, _09272_, _34581_);
  or _53980_ (_09274_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or _53981_ (_09275_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and _53982_ (_09276_, _09275_, _09274_);
  and _53983_ (_09277_, _09276_, _34796_);
  or _53984_ (_09278_, _09277_, _09273_);
  and _53985_ (_09279_, _09278_, _34772_);
  or _53986_ (_09280_, _09279_, _09269_);
  and _53987_ (_09281_, _09280_, _34719_);
  and _53988_ (_09282_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and _53989_ (_09283_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or _53990_ (_09284_, _09283_, _09282_);
  and _53991_ (_09285_, _09284_, _34581_);
  and _53992_ (_09286_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and _53993_ (_09287_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or _53994_ (_09288_, _09287_, _09286_);
  and _53995_ (_09289_, _09288_, _34796_);
  or _53996_ (_09290_, _09289_, _09285_);
  and _53997_ (_09291_, _09290_, _34790_);
  and _53998_ (_09292_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and _53999_ (_09293_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or _54000_ (_09294_, _09293_, _09292_);
  and _54001_ (_09295_, _09294_, _34581_);
  and _54002_ (_09296_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and _54003_ (_09297_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or _54004_ (_09298_, _09297_, _09296_);
  and _54005_ (_09299_, _09298_, _34796_);
  or _54006_ (_09300_, _09299_, _09295_);
  and _54007_ (_09301_, _09300_, _34772_);
  or _54008_ (_09302_, _09301_, _09291_);
  and _54009_ (_09303_, _09302_, _34803_);
  or _54010_ (_09304_, _09303_, _09281_);
  and _54011_ (_09305_, _09304_, _34700_);
  or _54012_ (_09306_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or _54013_ (_09307_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and _54014_ (_09308_, _09307_, _34796_);
  and _54015_ (_09309_, _09308_, _09306_);
  or _54016_ (_09310_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or _54017_ (_09311_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and _54018_ (_09312_, _09311_, _34581_);
  and _54019_ (_09313_, _09312_, _09310_);
  or _54020_ (_09314_, _09313_, _09309_);
  and _54021_ (_09315_, _09314_, _34790_);
  or _54022_ (_09316_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or _54023_ (_09317_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and _54024_ (_09318_, _09317_, _34796_);
  and _54025_ (_09319_, _09318_, _09316_);
  or _54026_ (_09320_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or _54027_ (_09321_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and _54028_ (_09322_, _09321_, _34581_);
  and _54029_ (_09323_, _09322_, _09320_);
  or _54030_ (_09324_, _09323_, _09319_);
  and _54031_ (_09325_, _09324_, _34772_);
  or _54032_ (_09326_, _09325_, _09315_);
  and _54033_ (_09327_, _09326_, _34719_);
  and _54034_ (_09328_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and _54035_ (_09329_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or _54036_ (_09330_, _09329_, _09328_);
  and _54037_ (_09331_, _09330_, _34581_);
  and _54038_ (_09332_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and _54039_ (_09333_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or _54040_ (_09334_, _09333_, _09332_);
  and _54041_ (_09335_, _09334_, _34796_);
  or _54042_ (_09336_, _09335_, _09331_);
  and _54043_ (_09337_, _09336_, _34790_);
  and _54044_ (_09338_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and _54045_ (_09339_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or _54046_ (_09340_, _09339_, _09338_);
  and _54047_ (_09341_, _09340_, _34581_);
  and _54048_ (_09342_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and _54049_ (_09343_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or _54050_ (_09344_, _09343_, _09342_);
  and _54051_ (_09345_, _09344_, _34796_);
  or _54052_ (_09346_, _09345_, _09341_);
  and _54053_ (_09347_, _09346_, _34772_);
  or _54054_ (_09348_, _09347_, _09337_);
  and _54055_ (_09349_, _09348_, _34803_);
  or _54056_ (_09350_, _09349_, _09327_);
  and _54057_ (_09351_, _09350_, _34789_);
  or _54058_ (_09352_, _09351_, _09305_);
  and _54059_ (_09353_, _09352_, _34638_);
  or _54060_ (_09354_, _09353_, _09259_);
  or _54061_ (_09355_, _09354_, _34985_);
  and _54062_ (_09356_, _09355_, _09165_);
  or _54063_ (_09357_, _09356_, _35178_);
  and _54064_ (_09358_, _09357_, _08975_);
  or _54065_ (_09359_, _09358_, _34788_);
  or _54066_ (_09360_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and _54067_ (_09361_, _09360_, _38997_);
  and _54068_ (_38984_[4], _09361_, _09359_);
  and _54069_ (_09362_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and _54070_ (_09363_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or _54071_ (_09364_, _09363_, _09362_);
  and _54072_ (_09365_, _09364_, _34581_);
  and _54073_ (_09366_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and _54074_ (_09367_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or _54075_ (_09368_, _09367_, _09366_);
  and _54076_ (_09369_, _09368_, _34796_);
  or _54077_ (_09370_, _09369_, _09365_);
  or _54078_ (_09371_, _09370_, _34790_);
  and _54079_ (_09372_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and _54080_ (_09373_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or _54081_ (_09374_, _09373_, _09372_);
  and _54082_ (_09375_, _09374_, _34581_);
  and _54083_ (_09376_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  and _54084_ (_09377_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or _54085_ (_09378_, _09377_, _09376_);
  and _54086_ (_09379_, _09378_, _34796_);
  or _54087_ (_09380_, _09379_, _09375_);
  or _54088_ (_09381_, _09380_, _34772_);
  and _54089_ (_09382_, _09381_, _34803_);
  and _54090_ (_09383_, _09382_, _09371_);
  or _54091_ (_09384_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or _54092_ (_09385_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and _54093_ (_09386_, _09385_, _09384_);
  and _54094_ (_09387_, _09386_, _34581_);
  or _54095_ (_09388_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or _54096_ (_09389_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and _54097_ (_09390_, _09389_, _09388_);
  and _54098_ (_09391_, _09390_, _34796_);
  or _54099_ (_09392_, _09391_, _09387_);
  or _54100_ (_09393_, _09392_, _34790_);
  or _54101_ (_09394_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or _54102_ (_09395_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and _54103_ (_09396_, _09395_, _09394_);
  and _54104_ (_09397_, _09396_, _34581_);
  or _54105_ (_09398_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or _54106_ (_09399_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and _54107_ (_09400_, _09399_, _09398_);
  and _54108_ (_09401_, _09400_, _34796_);
  or _54109_ (_09402_, _09401_, _09397_);
  or _54110_ (_09403_, _09402_, _34772_);
  and _54111_ (_09404_, _09403_, _34719_);
  and _54112_ (_09405_, _09404_, _09393_);
  or _54113_ (_09406_, _09405_, _09383_);
  and _54114_ (_09407_, _09406_, _34700_);
  and _54115_ (_09408_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and _54116_ (_09409_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or _54117_ (_09410_, _09409_, _09408_);
  and _54118_ (_09411_, _09410_, _34581_);
  and _54119_ (_09412_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and _54120_ (_09413_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or _54121_ (_09414_, _09413_, _09412_);
  and _54122_ (_09415_, _09414_, _34796_);
  or _54123_ (_09416_, _09415_, _09411_);
  or _54124_ (_09417_, _09416_, _34790_);
  and _54125_ (_09418_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and _54126_ (_09419_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or _54127_ (_09420_, _09419_, _09418_);
  and _54128_ (_09421_, _09420_, _34581_);
  and _54129_ (_09422_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and _54130_ (_09423_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or _54131_ (_09424_, _09423_, _09422_);
  and _54132_ (_09425_, _09424_, _34796_);
  or _54133_ (_09426_, _09425_, _09421_);
  or _54134_ (_09427_, _09426_, _34772_);
  and _54135_ (_09428_, _09427_, _34803_);
  and _54136_ (_09429_, _09428_, _09417_);
  or _54137_ (_09430_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or _54138_ (_09431_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  and _54139_ (_09432_, _09431_, _34796_);
  and _54140_ (_09433_, _09432_, _09430_);
  or _54141_ (_09434_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or _54142_ (_09435_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and _54143_ (_09436_, _09435_, _34581_);
  and _54144_ (_09437_, _09436_, _09434_);
  or _54145_ (_09438_, _09437_, _09433_);
  or _54146_ (_09439_, _09438_, _34790_);
  or _54147_ (_09440_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or _54148_ (_09441_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  and _54149_ (_09442_, _09441_, _34796_);
  and _54150_ (_09443_, _09442_, _09440_);
  or _54151_ (_09444_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or _54152_ (_09445_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and _54153_ (_09446_, _09445_, _34581_);
  and _54154_ (_09447_, _09446_, _09444_);
  or _54155_ (_09448_, _09447_, _09443_);
  or _54156_ (_09449_, _09448_, _34772_);
  and _54157_ (_09450_, _09449_, _34719_);
  and _54158_ (_09451_, _09450_, _09439_);
  or _54159_ (_09452_, _09451_, _09429_);
  and _54160_ (_09453_, _09452_, _34789_);
  or _54161_ (_09454_, _09453_, _09407_);
  and _54162_ (_09455_, _09454_, _34840_);
  and _54163_ (_09456_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and _54164_ (_09457_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or _54165_ (_09458_, _09457_, _09456_);
  and _54166_ (_09459_, _09458_, _34581_);
  and _54167_ (_09460_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and _54168_ (_09461_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or _54169_ (_09462_, _09461_, _09460_);
  and _54170_ (_09463_, _09462_, _34796_);
  or _54171_ (_09464_, _09463_, _09459_);
  and _54172_ (_09465_, _09464_, _34772_);
  and _54173_ (_09466_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and _54174_ (_09467_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _54175_ (_09468_, _09467_, _09466_);
  and _54176_ (_09469_, _09468_, _34581_);
  and _54177_ (_09470_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and _54178_ (_09471_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or _54179_ (_09472_, _09471_, _09470_);
  and _54180_ (_09473_, _09472_, _34796_);
  or _54181_ (_09474_, _09473_, _09469_);
  and _54182_ (_09475_, _09474_, _34790_);
  or _54183_ (_09476_, _09475_, _09465_);
  and _54184_ (_09477_, _09476_, _34803_);
  or _54185_ (_09478_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or _54186_ (_09479_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and _54187_ (_09480_, _09479_, _34796_);
  and _54188_ (_09481_, _09480_, _09478_);
  or _54189_ (_09482_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or _54190_ (_09483_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and _54191_ (_09484_, _09483_, _34581_);
  and _54192_ (_09485_, _09484_, _09482_);
  or _54193_ (_09486_, _09485_, _09481_);
  and _54194_ (_09487_, _09486_, _34772_);
  or _54195_ (_09488_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or _54196_ (_09489_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and _54197_ (_09490_, _09489_, _34796_);
  and _54198_ (_09491_, _09490_, _09488_);
  or _54199_ (_09492_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or _54200_ (_09493_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and _54201_ (_09494_, _09493_, _34581_);
  and _54202_ (_09495_, _09494_, _09492_);
  or _54203_ (_09496_, _09495_, _09491_);
  and _54204_ (_09497_, _09496_, _34790_);
  or _54205_ (_09498_, _09497_, _09487_);
  and _54206_ (_09499_, _09498_, _34719_);
  or _54207_ (_09500_, _09499_, _09477_);
  and _54208_ (_09501_, _09500_, _34789_);
  and _54209_ (_09502_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and _54210_ (_09503_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or _54211_ (_09504_, _09503_, _09502_);
  and _54212_ (_09505_, _09504_, _34581_);
  and _54213_ (_09506_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and _54214_ (_09507_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or _54215_ (_09508_, _09507_, _09506_);
  and _54216_ (_09509_, _09508_, _34796_);
  or _54217_ (_09510_, _09509_, _09505_);
  and _54218_ (_09511_, _09510_, _34772_);
  and _54219_ (_09512_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and _54220_ (_09513_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or _54221_ (_09514_, _09513_, _09512_);
  and _54222_ (_09515_, _09514_, _34581_);
  and _54223_ (_09516_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  and _54224_ (_09517_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or _54225_ (_09518_, _09517_, _09516_);
  and _54226_ (_09519_, _09518_, _34796_);
  or _54227_ (_09520_, _09519_, _09515_);
  and _54228_ (_09521_, _09520_, _34790_);
  or _54229_ (_09522_, _09521_, _09511_);
  and _54230_ (_09523_, _09522_, _34803_);
  or _54231_ (_09524_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or _54232_ (_09525_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  and _54233_ (_09526_, _09525_, _09524_);
  and _54234_ (_09527_, _09526_, _34581_);
  or _54235_ (_09528_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or _54236_ (_09529_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and _54237_ (_09530_, _09529_, _09528_);
  and _54238_ (_09531_, _09530_, _34796_);
  or _54239_ (_09532_, _09531_, _09527_);
  and _54240_ (_09533_, _09532_, _34772_);
  or _54241_ (_09534_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or _54242_ (_09535_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  and _54243_ (_09536_, _09535_, _09534_);
  and _54244_ (_09537_, _09536_, _34581_);
  or _54245_ (_09538_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or _54246_ (_09539_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and _54247_ (_09540_, _09539_, _09538_);
  and _54248_ (_09541_, _09540_, _34796_);
  or _54249_ (_09542_, _09541_, _09537_);
  and _54250_ (_09543_, _09542_, _34790_);
  or _54251_ (_09544_, _09543_, _09533_);
  and _54252_ (_09545_, _09544_, _34719_);
  or _54253_ (_09546_, _09545_, _09523_);
  and _54254_ (_09547_, _09546_, _34700_);
  or _54255_ (_09548_, _09547_, _09501_);
  and _54256_ (_09549_, _09548_, _34638_);
  or _54257_ (_09550_, _09549_, _09455_);
  or _54258_ (_09551_, _09550_, _34692_);
  and _54259_ (_09552_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and _54260_ (_09553_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or _54261_ (_09554_, _09553_, _09552_);
  and _54262_ (_09555_, _09554_, _34581_);
  and _54263_ (_09556_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and _54264_ (_09557_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or _54265_ (_09558_, _09557_, _09556_);
  and _54266_ (_09559_, _09558_, _34796_);
  or _54267_ (_09560_, _09559_, _09555_);
  or _54268_ (_09561_, _09560_, _34790_);
  and _54269_ (_09562_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and _54270_ (_09563_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or _54271_ (_09564_, _09563_, _09562_);
  and _54272_ (_09565_, _09564_, _34581_);
  and _54273_ (_09566_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and _54274_ (_09567_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or _54275_ (_09568_, _09567_, _09566_);
  and _54276_ (_09569_, _09568_, _34796_);
  or _54277_ (_09570_, _09569_, _09565_);
  or _54278_ (_09571_, _09570_, _34772_);
  and _54279_ (_09572_, _09571_, _34803_);
  and _54280_ (_09573_, _09572_, _09561_);
  or _54281_ (_09574_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or _54282_ (_09575_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and _54283_ (_09576_, _09575_, _34796_);
  and _54284_ (_09577_, _09576_, _09574_);
  or _54285_ (_09578_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or _54286_ (_09579_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and _54287_ (_09580_, _09579_, _34581_);
  and _54288_ (_09581_, _09580_, _09578_);
  or _54289_ (_09582_, _09581_, _09577_);
  or _54290_ (_09583_, _09582_, _34790_);
  or _54291_ (_09584_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or _54292_ (_09585_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  and _54293_ (_09586_, _09585_, _34796_);
  and _54294_ (_09587_, _09586_, _09584_);
  or _54295_ (_09588_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or _54296_ (_09589_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  and _54297_ (_09590_, _09589_, _34581_);
  and _54298_ (_09591_, _09590_, _09588_);
  or _54299_ (_09592_, _09591_, _09587_);
  or _54300_ (_09593_, _09592_, _34772_);
  and _54301_ (_09594_, _09593_, _34719_);
  and _54302_ (_09595_, _09594_, _09583_);
  or _54303_ (_09596_, _09595_, _09573_);
  and _54304_ (_09597_, _09596_, _34789_);
  and _54305_ (_09598_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and _54306_ (_09599_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or _54307_ (_09600_, _09599_, _09598_);
  and _54308_ (_09601_, _09600_, _34581_);
  and _54309_ (_09602_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and _54310_ (_09603_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or _54311_ (_09604_, _09603_, _09602_);
  and _54312_ (_09605_, _09604_, _34796_);
  or _54313_ (_09606_, _09605_, _09601_);
  or _54314_ (_09607_, _09606_, _34790_);
  and _54315_ (_09608_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and _54316_ (_09609_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or _54317_ (_09610_, _09609_, _09608_);
  and _54318_ (_09611_, _09610_, _34581_);
  and _54319_ (_09612_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and _54320_ (_09613_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or _54321_ (_09614_, _09613_, _09612_);
  and _54322_ (_09615_, _09614_, _34796_);
  or _54323_ (_09616_, _09615_, _09611_);
  or _54324_ (_09617_, _09616_, _34772_);
  and _54325_ (_09618_, _09617_, _34803_);
  and _54326_ (_09619_, _09618_, _09607_);
  or _54327_ (_09620_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or _54328_ (_09621_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and _54329_ (_09622_, _09621_, _09620_);
  and _54330_ (_09623_, _09622_, _34581_);
  or _54331_ (_09624_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or _54332_ (_09625_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and _54333_ (_09626_, _09625_, _09624_);
  and _54334_ (_09627_, _09626_, _34796_);
  or _54335_ (_09628_, _09627_, _09623_);
  or _54336_ (_09629_, _09628_, _34790_);
  or _54337_ (_09630_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or _54338_ (_09631_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and _54339_ (_09632_, _09631_, _09630_);
  and _54340_ (_09633_, _09632_, _34581_);
  or _54341_ (_09634_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or _54342_ (_09635_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and _54343_ (_09636_, _09635_, _09634_);
  and _54344_ (_09637_, _09636_, _34796_);
  or _54345_ (_09638_, _09637_, _09633_);
  or _54346_ (_09639_, _09638_, _34772_);
  and _54347_ (_09640_, _09639_, _34719_);
  and _54348_ (_09641_, _09640_, _09629_);
  or _54349_ (_09642_, _09641_, _09619_);
  and _54350_ (_09643_, _09642_, _34700_);
  or _54351_ (_09644_, _09643_, _09597_);
  and _54352_ (_09645_, _09644_, _34840_);
  or _54353_ (_09646_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or _54354_ (_09647_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  and _54355_ (_09648_, _09647_, _09646_);
  and _54356_ (_09649_, _09648_, _34581_);
  or _54357_ (_09650_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or _54358_ (_09651_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and _54359_ (_09652_, _09651_, _09650_);
  and _54360_ (_09653_, _09652_, _34796_);
  or _54361_ (_09654_, _09653_, _09649_);
  and _54362_ (_09655_, _09654_, _34790_);
  or _54363_ (_09656_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or _54364_ (_09657_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and _54365_ (_09658_, _09657_, _09656_);
  and _54366_ (_09659_, _09658_, _34581_);
  or _54367_ (_09660_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or _54368_ (_09661_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and _54369_ (_09662_, _09661_, _09660_);
  and _54370_ (_09663_, _09662_, _34796_);
  or _54371_ (_09664_, _09663_, _09659_);
  and _54372_ (_09665_, _09664_, _34772_);
  or _54373_ (_09666_, _09665_, _09655_);
  and _54374_ (_09667_, _09666_, _34719_);
  and _54375_ (_09668_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  and _54376_ (_09669_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or _54377_ (_09670_, _09669_, _09668_);
  and _54378_ (_09671_, _09670_, _34581_);
  and _54379_ (_09672_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  and _54380_ (_09673_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or _54381_ (_09674_, _09673_, _09672_);
  and _54382_ (_09675_, _09674_, _34796_);
  or _54383_ (_09676_, _09675_, _09671_);
  and _54384_ (_09677_, _09676_, _34790_);
  and _54385_ (_09678_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  and _54386_ (_09679_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or _54387_ (_09680_, _09679_, _09678_);
  and _54388_ (_09681_, _09680_, _34581_);
  and _54389_ (_09682_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and _54390_ (_09683_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or _54391_ (_09684_, _09683_, _09682_);
  and _54392_ (_09685_, _09684_, _34796_);
  or _54393_ (_09686_, _09685_, _09681_);
  and _54394_ (_09687_, _09686_, _34772_);
  or _54395_ (_09688_, _09687_, _09677_);
  and _54396_ (_09689_, _09688_, _34803_);
  or _54397_ (_09690_, _09689_, _09667_);
  and _54398_ (_09691_, _09690_, _34700_);
  or _54399_ (_09692_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or _54400_ (_09693_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and _54401_ (_09694_, _09693_, _34796_);
  and _54402_ (_09695_, _09694_, _09692_);
  or _54403_ (_09696_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or _54404_ (_09697_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and _54405_ (_09698_, _09697_, _34581_);
  and _54406_ (_09699_, _09698_, _09696_);
  or _54407_ (_09700_, _09699_, _09695_);
  and _54408_ (_09701_, _09700_, _34790_);
  or _54409_ (_09702_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or _54410_ (_09703_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and _54411_ (_09704_, _09703_, _34796_);
  and _54412_ (_09705_, _09704_, _09702_);
  or _54413_ (_09706_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or _54414_ (_09707_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  and _54415_ (_09708_, _09707_, _34581_);
  and _54416_ (_09709_, _09708_, _09706_);
  or _54417_ (_09710_, _09709_, _09705_);
  and _54418_ (_09711_, _09710_, _34772_);
  or _54419_ (_09712_, _09711_, _09701_);
  and _54420_ (_09713_, _09712_, _34719_);
  and _54421_ (_09714_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  and _54422_ (_09715_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or _54423_ (_09716_, _09715_, _09714_);
  and _54424_ (_09717_, _09716_, _34581_);
  and _54425_ (_09718_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and _54426_ (_09719_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or _54427_ (_09720_, _09719_, _09718_);
  and _54428_ (_09721_, _09720_, _34796_);
  or _54429_ (_09722_, _09721_, _09717_);
  and _54430_ (_09723_, _09722_, _34790_);
  and _54431_ (_09724_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and _54432_ (_09725_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or _54433_ (_09726_, _09725_, _09724_);
  and _54434_ (_09727_, _09726_, _34581_);
  and _54435_ (_09728_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and _54436_ (_09729_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or _54437_ (_09730_, _09729_, _09728_);
  and _54438_ (_09731_, _09730_, _34796_);
  or _54439_ (_09732_, _09731_, _09727_);
  and _54440_ (_09733_, _09732_, _34772_);
  or _54441_ (_09734_, _09733_, _09723_);
  and _54442_ (_09735_, _09734_, _34803_);
  or _54443_ (_09736_, _09735_, _09713_);
  and _54444_ (_09737_, _09736_, _34789_);
  or _54445_ (_09738_, _09737_, _09691_);
  and _54446_ (_09739_, _09738_, _34638_);
  or _54447_ (_09740_, _09739_, _09645_);
  or _54448_ (_09741_, _09740_, _34985_);
  and _54449_ (_09742_, _09741_, _09551_);
  or _54450_ (_09743_, _09742_, _34346_);
  and _54451_ (_09744_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and _54452_ (_09745_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or _54453_ (_09746_, _09745_, _09744_);
  and _54454_ (_09747_, _09746_, _34581_);
  and _54455_ (_09748_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and _54456_ (_09749_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or _54457_ (_09750_, _09749_, _09748_);
  and _54458_ (_09751_, _09750_, _34796_);
  or _54459_ (_09752_, _09751_, _09747_);
  and _54460_ (_09753_, _09752_, _34772_);
  and _54461_ (_09754_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and _54462_ (_09755_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or _54463_ (_09756_, _09755_, _09754_);
  and _54464_ (_09757_, _09756_, _34581_);
  and _54465_ (_09758_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and _54466_ (_09759_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or _54467_ (_09760_, _09759_, _09758_);
  and _54468_ (_09761_, _09760_, _34796_);
  or _54469_ (_09762_, _09761_, _09757_);
  and _54470_ (_09763_, _09762_, _34790_);
  or _54471_ (_09764_, _09763_, _09753_);
  and _54472_ (_09765_, _09764_, _34803_);
  or _54473_ (_09766_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or _54474_ (_09767_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and _54475_ (_09768_, _09767_, _34796_);
  and _54476_ (_09769_, _09768_, _09766_);
  or _54477_ (_09770_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or _54478_ (_09771_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and _54479_ (_09772_, _09771_, _34581_);
  and _54480_ (_09773_, _09772_, _09770_);
  or _54481_ (_09774_, _09773_, _09769_);
  and _54482_ (_09775_, _09774_, _34772_);
  or _54483_ (_09776_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or _54484_ (_09777_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and _54485_ (_09778_, _09777_, _34796_);
  and _54486_ (_09779_, _09778_, _09776_);
  or _54487_ (_09780_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or _54488_ (_09781_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and _54489_ (_09782_, _09781_, _34581_);
  and _54490_ (_09783_, _09782_, _09780_);
  or _54491_ (_09784_, _09783_, _09779_);
  and _54492_ (_09785_, _09784_, _34790_);
  or _54493_ (_09786_, _09785_, _09775_);
  and _54494_ (_09787_, _09786_, _34719_);
  or _54495_ (_09788_, _09787_, _09765_);
  and _54496_ (_09789_, _09788_, _34789_);
  and _54497_ (_09790_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and _54498_ (_09791_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or _54499_ (_09792_, _09791_, _09790_);
  and _54500_ (_09793_, _09792_, _34581_);
  and _54501_ (_09794_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and _54502_ (_09795_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or _54503_ (_09796_, _09795_, _09794_);
  and _54504_ (_09797_, _09796_, _34796_);
  or _54505_ (_09798_, _09797_, _09793_);
  and _54506_ (_09799_, _09798_, _34772_);
  and _54507_ (_09800_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and _54508_ (_09801_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or _54509_ (_09802_, _09801_, _09800_);
  and _54510_ (_09803_, _09802_, _34581_);
  and _54511_ (_09804_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and _54512_ (_09805_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or _54513_ (_09806_, _09805_, _09804_);
  and _54514_ (_09807_, _09806_, _34796_);
  or _54515_ (_09808_, _09807_, _09803_);
  and _54516_ (_09809_, _09808_, _34790_);
  or _54517_ (_09810_, _09809_, _09799_);
  and _54518_ (_09811_, _09810_, _34803_);
  or _54519_ (_09812_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or _54520_ (_09813_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and _54521_ (_09814_, _09813_, _09812_);
  and _54522_ (_09815_, _09814_, _34581_);
  or _54523_ (_09816_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or _54524_ (_09817_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and _54525_ (_09818_, _09817_, _09816_);
  and _54526_ (_09819_, _09818_, _34796_);
  or _54527_ (_09820_, _09819_, _09815_);
  and _54528_ (_09821_, _09820_, _34772_);
  or _54529_ (_09822_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or _54530_ (_09823_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and _54531_ (_09824_, _09823_, _09822_);
  and _54532_ (_09825_, _09824_, _34581_);
  or _54533_ (_09826_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or _54534_ (_09827_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and _54535_ (_09828_, _09827_, _09826_);
  and _54536_ (_09829_, _09828_, _34796_);
  or _54537_ (_09830_, _09829_, _09825_);
  and _54538_ (_09831_, _09830_, _34790_);
  or _54539_ (_09832_, _09831_, _09821_);
  and _54540_ (_09833_, _09832_, _34719_);
  or _54541_ (_09834_, _09833_, _09811_);
  and _54542_ (_09835_, _09834_, _34700_);
  or _54543_ (_09836_, _09835_, _09789_);
  and _54544_ (_09837_, _09836_, _34638_);
  and _54545_ (_09838_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and _54546_ (_09839_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or _54547_ (_09840_, _09839_, _09838_);
  and _54548_ (_09841_, _09840_, _34581_);
  and _54549_ (_09842_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and _54550_ (_09843_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or _54551_ (_09844_, _09843_, _09842_);
  and _54552_ (_09845_, _09844_, _34796_);
  or _54553_ (_09846_, _09845_, _09841_);
  or _54554_ (_09847_, _09846_, _34790_);
  and _54555_ (_09848_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and _54556_ (_09849_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or _54557_ (_09850_, _09849_, _09848_);
  and _54558_ (_09851_, _09850_, _34581_);
  and _54559_ (_09852_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and _54560_ (_09853_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or _54561_ (_09854_, _09853_, _09852_);
  and _54562_ (_09855_, _09854_, _34796_);
  or _54563_ (_09856_, _09855_, _09851_);
  or _54564_ (_09857_, _09856_, _34772_);
  and _54565_ (_09858_, _09857_, _34803_);
  and _54566_ (_09859_, _09858_, _09847_);
  or _54567_ (_09860_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or _54568_ (_09861_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and _54569_ (_09862_, _09861_, _09860_);
  and _54570_ (_09863_, _09862_, _34581_);
  or _54571_ (_09864_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or _54572_ (_09865_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and _54573_ (_09866_, _09865_, _09864_);
  and _54574_ (_09867_, _09866_, _34796_);
  or _54575_ (_09868_, _09867_, _09863_);
  or _54576_ (_09869_, _09868_, _34790_);
  or _54577_ (_09870_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or _54578_ (_09871_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and _54579_ (_09872_, _09871_, _09870_);
  and _54580_ (_09873_, _09872_, _34581_);
  or _54581_ (_09874_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or _54582_ (_09875_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and _54583_ (_09876_, _09875_, _09874_);
  and _54584_ (_09877_, _09876_, _34796_);
  or _54585_ (_09878_, _09877_, _09873_);
  or _54586_ (_09879_, _09878_, _34772_);
  and _54587_ (_09880_, _09879_, _34719_);
  and _54588_ (_09881_, _09880_, _09869_);
  or _54589_ (_09882_, _09881_, _09859_);
  and _54590_ (_09883_, _09882_, _34700_);
  and _54591_ (_09884_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and _54592_ (_09885_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or _54593_ (_09886_, _09885_, _09884_);
  and _54594_ (_09887_, _09886_, _34581_);
  and _54595_ (_09888_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and _54596_ (_09889_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or _54597_ (_09890_, _09889_, _09888_);
  and _54598_ (_09891_, _09890_, _34796_);
  or _54599_ (_09892_, _09891_, _09887_);
  or _54600_ (_09893_, _09892_, _34790_);
  and _54601_ (_09894_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and _54602_ (_09895_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or _54603_ (_09896_, _09895_, _09894_);
  and _54604_ (_09897_, _09896_, _34581_);
  and _54605_ (_09898_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and _54606_ (_09899_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or _54607_ (_09900_, _09899_, _09898_);
  and _54608_ (_09901_, _09900_, _34796_);
  or _54609_ (_09902_, _09901_, _09897_);
  or _54610_ (_09903_, _09902_, _34772_);
  and _54611_ (_09904_, _09903_, _34803_);
  and _54612_ (_09905_, _09904_, _09893_);
  or _54613_ (_09906_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or _54614_ (_09907_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and _54615_ (_09908_, _09907_, _34796_);
  and _54616_ (_09909_, _09908_, _09906_);
  or _54617_ (_09910_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or _54618_ (_09911_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and _54619_ (_09912_, _09911_, _34581_);
  and _54620_ (_09913_, _09912_, _09910_);
  or _54621_ (_09914_, _09913_, _09909_);
  or _54622_ (_09915_, _09914_, _34790_);
  or _54623_ (_09916_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or _54624_ (_09917_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and _54625_ (_09918_, _09917_, _34796_);
  and _54626_ (_09919_, _09918_, _09916_);
  or _54627_ (_09920_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or _54628_ (_09921_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and _54629_ (_09922_, _09921_, _34581_);
  and _54630_ (_09923_, _09922_, _09920_);
  or _54631_ (_09924_, _09923_, _09919_);
  or _54632_ (_09925_, _09924_, _34772_);
  and _54633_ (_09926_, _09925_, _34719_);
  and _54634_ (_09927_, _09926_, _09915_);
  or _54635_ (_09928_, _09927_, _09905_);
  and _54636_ (_09929_, _09928_, _34789_);
  or _54637_ (_09930_, _09929_, _09883_);
  and _54638_ (_09931_, _09930_, _34840_);
  or _54639_ (_09932_, _09931_, _09837_);
  or _54640_ (_09933_, _09932_, _34692_);
  and _54641_ (_09934_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and _54642_ (_09935_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or _54643_ (_09936_, _09935_, _09934_);
  and _54644_ (_09937_, _09936_, _34796_);
  and _54645_ (_09938_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and _54646_ (_09939_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or _54647_ (_09940_, _09939_, _09938_);
  and _54648_ (_09941_, _09940_, _34581_);
  or _54649_ (_09942_, _09941_, _09937_);
  or _54650_ (_09943_, _09942_, _34790_);
  and _54651_ (_09944_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and _54652_ (_09945_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or _54653_ (_09946_, _09945_, _09944_);
  and _54654_ (_09947_, _09946_, _34796_);
  and _54655_ (_09948_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and _54656_ (_09949_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or _54657_ (_09950_, _09949_, _09948_);
  and _54658_ (_09951_, _09950_, _34581_);
  or _54659_ (_09952_, _09951_, _09947_);
  or _54660_ (_09953_, _09952_, _34772_);
  and _54661_ (_09954_, _09953_, _34803_);
  and _54662_ (_09955_, _09954_, _09943_);
  or _54663_ (_09956_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or _54664_ (_09957_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and _54665_ (_09958_, _09957_, _34581_);
  and _54666_ (_09959_, _09958_, _09956_);
  or _54667_ (_09960_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or _54668_ (_09961_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and _54669_ (_09962_, _09961_, _34796_);
  and _54670_ (_09963_, _09962_, _09960_);
  or _54671_ (_09964_, _09963_, _09959_);
  or _54672_ (_09965_, _09964_, _34790_);
  or _54673_ (_09966_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or _54674_ (_09967_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and _54675_ (_09968_, _09967_, _34581_);
  and _54676_ (_09969_, _09968_, _09966_);
  or _54677_ (_09970_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or _54678_ (_09971_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and _54679_ (_09972_, _09971_, _34796_);
  and _54680_ (_09973_, _09972_, _09970_);
  or _54681_ (_09974_, _09973_, _09969_);
  or _54682_ (_09975_, _09974_, _34772_);
  and _54683_ (_09976_, _09975_, _34719_);
  and _54684_ (_09977_, _09976_, _09965_);
  or _54685_ (_09978_, _09977_, _09955_);
  and _54686_ (_09979_, _09978_, _34789_);
  and _54687_ (_09980_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and _54688_ (_09981_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or _54689_ (_09982_, _09981_, _34581_);
  or _54690_ (_09983_, _09982_, _09980_);
  and _54691_ (_09984_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and _54692_ (_09985_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or _54693_ (_09986_, _09985_, _34796_);
  or _54694_ (_09987_, _09986_, _09984_);
  and _54695_ (_09988_, _09987_, _09983_);
  or _54696_ (_09989_, _09988_, _34790_);
  and _54697_ (_09990_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and _54698_ (_09991_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or _54699_ (_09992_, _09991_, _34581_);
  or _54700_ (_09993_, _09992_, _09990_);
  and _54701_ (_09994_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and _54702_ (_09995_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or _54703_ (_09996_, _09995_, _34796_);
  or _54704_ (_09997_, _09996_, _09994_);
  and _54705_ (_09998_, _09997_, _09993_);
  or _54706_ (_09999_, _09998_, _34772_);
  and _54707_ (_10000_, _09999_, _34803_);
  and _54708_ (_10001_, _10000_, _09989_);
  or _54709_ (_10002_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or _54710_ (_10003_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and _54711_ (_10004_, _10003_, _10002_);
  or _54712_ (_10005_, _10004_, _34796_);
  or _54713_ (_10006_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or _54714_ (_10007_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and _54715_ (_10008_, _10007_, _10006_);
  or _54716_ (_10009_, _10008_, _34581_);
  and _54717_ (_10010_, _10009_, _10005_);
  or _54718_ (_10011_, _10010_, _34790_);
  or _54719_ (_10012_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or _54720_ (_10013_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and _54721_ (_10014_, _10013_, _10012_);
  or _54722_ (_10015_, _10014_, _34796_);
  or _54723_ (_10016_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or _54724_ (_10017_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and _54725_ (_10018_, _10017_, _10016_);
  or _54726_ (_10019_, _10018_, _34581_);
  and _54727_ (_10020_, _10019_, _10015_);
  or _54728_ (_10021_, _10020_, _34772_);
  and _54729_ (_10022_, _10021_, _34719_);
  and _54730_ (_10023_, _10022_, _10011_);
  or _54731_ (_10024_, _10023_, _10001_);
  and _54732_ (_10025_, _10024_, _34700_);
  or _54733_ (_10026_, _10025_, _09979_);
  and _54734_ (_10027_, _10026_, _34840_);
  and _54735_ (_10028_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and _54736_ (_10029_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or _54737_ (_10030_, _10029_, _10028_);
  and _54738_ (_10031_, _10030_, _34581_);
  and _54739_ (_10032_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and _54740_ (_10033_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or _54741_ (_10034_, _10033_, _10032_);
  and _54742_ (_10035_, _10034_, _34796_);
  or _54743_ (_10036_, _10035_, _10031_);
  and _54744_ (_10037_, _10036_, _34772_);
  and _54745_ (_10038_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and _54746_ (_10039_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or _54747_ (_10040_, _10039_, _10038_);
  and _54748_ (_10041_, _10040_, _34581_);
  and _54749_ (_10042_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and _54750_ (_10043_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or _54751_ (_10044_, _10043_, _10042_);
  and _54752_ (_10045_, _10044_, _34796_);
  or _54753_ (_10046_, _10045_, _10041_);
  and _54754_ (_10047_, _10046_, _34790_);
  or _54755_ (_10048_, _10047_, _10037_);
  and _54756_ (_10049_, _10048_, _34803_);
  or _54757_ (_10050_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or _54758_ (_10051_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and _54759_ (_10052_, _10051_, _10050_);
  and _54760_ (_10053_, _10052_, _34581_);
  or _54761_ (_10054_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or _54762_ (_10055_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and _54763_ (_10056_, _10055_, _10054_);
  and _54764_ (_10057_, _10056_, _34796_);
  or _54765_ (_10058_, _10057_, _10053_);
  and _54766_ (_10059_, _10058_, _34772_);
  or _54767_ (_10060_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or _54768_ (_10061_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and _54769_ (_10062_, _10061_, _10060_);
  and _54770_ (_10063_, _10062_, _34581_);
  or _54771_ (_10064_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or _54772_ (_10065_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and _54773_ (_10066_, _10065_, _10064_);
  and _54774_ (_10067_, _10066_, _34796_);
  or _54775_ (_10068_, _10067_, _10063_);
  and _54776_ (_10069_, _10068_, _34790_);
  or _54777_ (_10070_, _10069_, _10059_);
  and _54778_ (_10071_, _10070_, _34719_);
  or _54779_ (_10072_, _10071_, _10049_);
  and _54780_ (_10073_, _10072_, _34700_);
  and _54781_ (_10074_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  and _54782_ (_10075_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or _54783_ (_10076_, _10075_, _10074_);
  and _54784_ (_10077_, _10076_, _34581_);
  and _54785_ (_10078_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  and _54786_ (_10079_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or _54787_ (_10080_, _10079_, _10078_);
  and _54788_ (_10081_, _10080_, _34796_);
  or _54789_ (_10082_, _10081_, _10077_);
  and _54790_ (_10083_, _10082_, _34772_);
  and _54791_ (_10084_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  and _54792_ (_10085_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or _54793_ (_10086_, _10085_, _10084_);
  and _54794_ (_10087_, _10086_, _34581_);
  and _54795_ (_10088_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  and _54796_ (_10089_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or _54797_ (_10090_, _10089_, _10088_);
  and _54798_ (_10091_, _10090_, _34796_);
  or _54799_ (_10092_, _10091_, _10087_);
  and _54800_ (_10093_, _10092_, _34790_);
  or _54801_ (_10094_, _10093_, _10083_);
  and _54802_ (_10095_, _10094_, _34803_);
  or _54803_ (_10096_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or _54804_ (_10097_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  and _54805_ (_10098_, _10097_, _10096_);
  and _54806_ (_10099_, _10098_, _34581_);
  or _54807_ (_10100_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or _54808_ (_10101_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  and _54809_ (_10102_, _10101_, _10100_);
  and _54810_ (_10103_, _10102_, _34796_);
  or _54811_ (_10104_, _10103_, _10099_);
  and _54812_ (_10105_, _10104_, _34772_);
  or _54813_ (_10106_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or _54814_ (_10107_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  and _54815_ (_10108_, _10107_, _10106_);
  and _54816_ (_10109_, _10108_, _34581_);
  or _54817_ (_10110_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or _54818_ (_10111_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  and _54819_ (_10112_, _10111_, _10110_);
  and _54820_ (_10113_, _10112_, _34796_);
  or _54821_ (_10114_, _10113_, _10109_);
  and _54822_ (_10115_, _10114_, _34790_);
  or _54823_ (_10116_, _10115_, _10105_);
  and _54824_ (_10117_, _10116_, _34719_);
  or _54825_ (_10118_, _10117_, _10095_);
  and _54826_ (_10119_, _10118_, _34789_);
  or _54827_ (_10120_, _10119_, _10073_);
  and _54828_ (_10121_, _10120_, _34638_);
  or _54829_ (_10122_, _10121_, _10027_);
  or _54830_ (_10123_, _10122_, _34985_);
  and _54831_ (_10124_, _10123_, _09933_);
  or _54832_ (_10125_, _10124_, _35178_);
  and _54833_ (_10126_, _10125_, _09743_);
  or _54834_ (_10127_, _10126_, _34788_);
  or _54835_ (_10128_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and _54836_ (_10129_, _10128_, _38997_);
  and _54837_ (_38984_[5], _10129_, _10127_);
  and _54838_ (_10130_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and _54839_ (_10131_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or _54840_ (_10132_, _10131_, _10130_);
  and _54841_ (_10133_, _10132_, _34581_);
  and _54842_ (_10134_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and _54843_ (_10135_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or _54844_ (_10136_, _10135_, _10134_);
  and _54845_ (_10137_, _10136_, _34796_);
  or _54846_ (_10138_, _10137_, _10133_);
  or _54847_ (_10139_, _10138_, _34790_);
  and _54848_ (_10140_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and _54849_ (_10141_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or _54850_ (_10142_, _10141_, _10140_);
  and _54851_ (_10143_, _10142_, _34581_);
  and _54852_ (_10144_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and _54853_ (_10145_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or _54854_ (_10146_, _10145_, _10144_);
  and _54855_ (_10147_, _10146_, _34796_);
  or _54856_ (_10148_, _10147_, _10143_);
  or _54857_ (_10149_, _10148_, _34772_);
  and _54858_ (_10150_, _10149_, _34803_);
  and _54859_ (_10151_, _10150_, _10139_);
  or _54860_ (_10152_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or _54861_ (_10153_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and _54862_ (_10154_, _10153_, _10152_);
  and _54863_ (_10155_, _10154_, _34581_);
  or _54864_ (_10156_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or _54865_ (_10157_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and _54866_ (_10158_, _10157_, _10156_);
  and _54867_ (_10159_, _10158_, _34796_);
  or _54868_ (_10160_, _10159_, _10155_);
  or _54869_ (_10161_, _10160_, _34790_);
  or _54870_ (_10162_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or _54871_ (_10163_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  and _54872_ (_10164_, _10163_, _10162_);
  and _54873_ (_10165_, _10164_, _34581_);
  or _54874_ (_10166_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or _54875_ (_10167_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and _54876_ (_10168_, _10167_, _10166_);
  and _54877_ (_10169_, _10168_, _34796_);
  or _54878_ (_10170_, _10169_, _10165_);
  or _54879_ (_10171_, _10170_, _34772_);
  and _54880_ (_10172_, _10171_, _34719_);
  and _54881_ (_10173_, _10172_, _10161_);
  or _54882_ (_10174_, _10173_, _10151_);
  and _54883_ (_10175_, _10174_, _34700_);
  and _54884_ (_10176_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and _54885_ (_10177_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or _54886_ (_10178_, _10177_, _10176_);
  and _54887_ (_10179_, _10178_, _34581_);
  and _54888_ (_10180_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and _54889_ (_10181_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or _54890_ (_10182_, _10181_, _10180_);
  and _54891_ (_10183_, _10182_, _34796_);
  or _54892_ (_10184_, _10183_, _10179_);
  or _54893_ (_10185_, _10184_, _34790_);
  and _54894_ (_10186_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and _54895_ (_10187_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or _54896_ (_10188_, _10187_, _10186_);
  and _54897_ (_10189_, _10188_, _34581_);
  and _54898_ (_10190_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and _54899_ (_10191_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or _54900_ (_10192_, _10191_, _10190_);
  and _54901_ (_10193_, _10192_, _34796_);
  or _54902_ (_10194_, _10193_, _10189_);
  or _54903_ (_10195_, _10194_, _34772_);
  and _54904_ (_10196_, _10195_, _34803_);
  and _54905_ (_10197_, _10196_, _10185_);
  or _54906_ (_10198_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or _54907_ (_10199_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and _54908_ (_10200_, _10199_, _34796_);
  and _54909_ (_10201_, _10200_, _10198_);
  or _54910_ (_10202_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or _54911_ (_10203_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and _54912_ (_10204_, _10203_, _34581_);
  and _54913_ (_10205_, _10204_, _10202_);
  or _54914_ (_10206_, _10205_, _10201_);
  or _54915_ (_10207_, _10206_, _34790_);
  or _54916_ (_10208_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or _54917_ (_10209_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and _54918_ (_10210_, _10209_, _34796_);
  and _54919_ (_10211_, _10210_, _10208_);
  or _54920_ (_10212_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or _54921_ (_10213_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and _54922_ (_10214_, _10213_, _34581_);
  and _54923_ (_10215_, _10214_, _10212_);
  or _54924_ (_10216_, _10215_, _10211_);
  or _54925_ (_10217_, _10216_, _34772_);
  and _54926_ (_10218_, _10217_, _34719_);
  and _54927_ (_10219_, _10218_, _10207_);
  or _54928_ (_10220_, _10219_, _10197_);
  and _54929_ (_10221_, _10220_, _34789_);
  or _54930_ (_10222_, _10221_, _10175_);
  and _54931_ (_10223_, _10222_, _34840_);
  and _54932_ (_10224_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and _54933_ (_10225_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or _54934_ (_10226_, _10225_, _10224_);
  and _54935_ (_10227_, _10226_, _34581_);
  and _54936_ (_10228_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and _54937_ (_10229_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or _54938_ (_10230_, _10229_, _10228_);
  and _54939_ (_10231_, _10230_, _34796_);
  or _54940_ (_10232_, _10231_, _10227_);
  and _54941_ (_10233_, _10232_, _34772_);
  and _54942_ (_10234_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and _54943_ (_10235_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _54944_ (_10236_, _10235_, _10234_);
  and _54945_ (_10237_, _10236_, _34581_);
  and _54946_ (_10238_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and _54947_ (_10239_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _54948_ (_10240_, _10239_, _10238_);
  and _54949_ (_10241_, _10240_, _34796_);
  or _54950_ (_10242_, _10241_, _10237_);
  and _54951_ (_10243_, _10242_, _34790_);
  or _54952_ (_10244_, _10243_, _10233_);
  and _54953_ (_10245_, _10244_, _34803_);
  or _54954_ (_10246_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or _54955_ (_10247_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and _54956_ (_10248_, _10247_, _34796_);
  and _54957_ (_10249_, _10248_, _10246_);
  or _54958_ (_10250_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _54959_ (_10251_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and _54960_ (_10252_, _10251_, _34581_);
  and _54961_ (_10253_, _10252_, _10250_);
  or _54962_ (_10254_, _10253_, _10249_);
  and _54963_ (_10255_, _10254_, _34772_);
  or _54964_ (_10256_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or _54965_ (_10257_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and _54966_ (_10258_, _10257_, _34796_);
  and _54967_ (_10259_, _10258_, _10256_);
  or _54968_ (_10260_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or _54969_ (_10261_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and _54970_ (_10262_, _10261_, _34581_);
  and _54971_ (_10263_, _10262_, _10260_);
  or _54972_ (_10264_, _10263_, _10259_);
  and _54973_ (_10265_, _10264_, _34790_);
  or _54974_ (_10266_, _10265_, _10255_);
  and _54975_ (_10267_, _10266_, _34719_);
  or _54976_ (_10268_, _10267_, _10245_);
  and _54977_ (_10269_, _10268_, _34789_);
  and _54978_ (_10270_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  and _54979_ (_10271_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or _54980_ (_10272_, _10271_, _10270_);
  and _54981_ (_10273_, _10272_, _34581_);
  and _54982_ (_10274_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and _54983_ (_10275_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or _54984_ (_10276_, _10275_, _10274_);
  and _54985_ (_10277_, _10276_, _34796_);
  or _54986_ (_10278_, _10277_, _10273_);
  and _54987_ (_10279_, _10278_, _34772_);
  and _54988_ (_10280_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  and _54989_ (_10281_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or _54990_ (_10282_, _10281_, _10280_);
  and _54991_ (_10283_, _10282_, _34581_);
  and _54992_ (_10284_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  and _54993_ (_10285_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or _54994_ (_10286_, _10285_, _10284_);
  and _54995_ (_10287_, _10286_, _34796_);
  or _54996_ (_10288_, _10287_, _10283_);
  and _54997_ (_10289_, _10288_, _34790_);
  or _54998_ (_10290_, _10289_, _10279_);
  and _54999_ (_10291_, _10290_, _34803_);
  or _55000_ (_10292_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or _55001_ (_10293_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  and _55002_ (_10294_, _10293_, _10292_);
  and _55003_ (_10295_, _10294_, _34581_);
  or _55004_ (_10296_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or _55005_ (_10297_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and _55006_ (_10298_, _10297_, _10296_);
  and _55007_ (_10299_, _10298_, _34796_);
  or _55008_ (_10300_, _10299_, _10295_);
  and _55009_ (_10301_, _10300_, _34772_);
  or _55010_ (_10302_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or _55011_ (_10303_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  and _55012_ (_10304_, _10303_, _10302_);
  and _55013_ (_10305_, _10304_, _34581_);
  or _55014_ (_10306_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or _55015_ (_10307_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and _55016_ (_10308_, _10307_, _10306_);
  and _55017_ (_10309_, _10308_, _34796_);
  or _55018_ (_10310_, _10309_, _10305_);
  and _55019_ (_10311_, _10310_, _34790_);
  or _55020_ (_10312_, _10311_, _10301_);
  and _55021_ (_10313_, _10312_, _34719_);
  or _55022_ (_10314_, _10313_, _10291_);
  and _55023_ (_10315_, _10314_, _34700_);
  or _55024_ (_10316_, _10315_, _10269_);
  and _55025_ (_10317_, _10316_, _34638_);
  or _55026_ (_10318_, _10317_, _10223_);
  or _55027_ (_10319_, _10318_, _34692_);
  and _55028_ (_10320_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  and _55029_ (_10321_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or _55030_ (_10322_, _10321_, _10320_);
  and _55031_ (_10323_, _10322_, _34581_);
  and _55032_ (_10324_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and _55033_ (_10325_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or _55034_ (_10326_, _10325_, _10324_);
  and _55035_ (_10327_, _10326_, _34796_);
  or _55036_ (_10328_, _10327_, _10323_);
  or _55037_ (_10329_, _10328_, _34790_);
  and _55038_ (_10330_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and _55039_ (_10331_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or _55040_ (_10332_, _10331_, _10330_);
  and _55041_ (_10333_, _10332_, _34581_);
  and _55042_ (_10334_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  and _55043_ (_10335_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or _55044_ (_10336_, _10335_, _10334_);
  and _55045_ (_10337_, _10336_, _34796_);
  or _55046_ (_10338_, _10337_, _10333_);
  or _55047_ (_10339_, _10338_, _34772_);
  and _55048_ (_10340_, _10339_, _34803_);
  and _55049_ (_10341_, _10340_, _10329_);
  or _55050_ (_10342_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or _55051_ (_10343_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and _55052_ (_10344_, _10343_, _34796_);
  and _55053_ (_10345_, _10344_, _10342_);
  or _55054_ (_10346_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or _55055_ (_10347_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and _55056_ (_10348_, _10347_, _34581_);
  and _55057_ (_10349_, _10348_, _10346_);
  or _55058_ (_10350_, _10349_, _10345_);
  or _55059_ (_10351_, _10350_, _34790_);
  or _55060_ (_10352_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or _55061_ (_10353_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and _55062_ (_10354_, _10353_, _34796_);
  and _55063_ (_10355_, _10354_, _10352_);
  or _55064_ (_10356_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or _55065_ (_10357_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and _55066_ (_10358_, _10357_, _34581_);
  and _55067_ (_10359_, _10358_, _10356_);
  or _55068_ (_10360_, _10359_, _10355_);
  or _55069_ (_10361_, _10360_, _34772_);
  and _55070_ (_10362_, _10361_, _34719_);
  and _55071_ (_10363_, _10362_, _10351_);
  or _55072_ (_10364_, _10363_, _10341_);
  and _55073_ (_10365_, _10364_, _34789_);
  and _55074_ (_10366_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and _55075_ (_10367_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or _55076_ (_10368_, _10367_, _10366_);
  and _55077_ (_10369_, _10368_, _34581_);
  and _55078_ (_10370_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and _55079_ (_10371_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or _55080_ (_10372_, _10371_, _10370_);
  and _55081_ (_10373_, _10372_, _34796_);
  or _55082_ (_10374_, _10373_, _10369_);
  or _55083_ (_10375_, _10374_, _34790_);
  and _55084_ (_10376_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and _55085_ (_10377_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or _55086_ (_10378_, _10377_, _10376_);
  and _55087_ (_10379_, _10378_, _34581_);
  and _55088_ (_10380_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and _55089_ (_10381_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or _55090_ (_10382_, _10381_, _10380_);
  and _55091_ (_10383_, _10382_, _34796_);
  or _55092_ (_10384_, _10383_, _10379_);
  or _55093_ (_10385_, _10384_, _34772_);
  and _55094_ (_10386_, _10385_, _34803_);
  and _55095_ (_10387_, _10386_, _10375_);
  or _55096_ (_10388_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or _55097_ (_10389_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and _55098_ (_10390_, _10389_, _10388_);
  and _55099_ (_10391_, _10390_, _34581_);
  or _55100_ (_10392_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or _55101_ (_10393_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and _55102_ (_10394_, _10393_, _10392_);
  and _55103_ (_10395_, _10394_, _34796_);
  or _55104_ (_10396_, _10395_, _10391_);
  or _55105_ (_10397_, _10396_, _34790_);
  or _55106_ (_10398_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or _55107_ (_10399_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and _55108_ (_10400_, _10399_, _10398_);
  and _55109_ (_10401_, _10400_, _34581_);
  or _55110_ (_10402_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or _55111_ (_10403_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and _55112_ (_10404_, _10403_, _10402_);
  and _55113_ (_10405_, _10404_, _34796_);
  or _55114_ (_10406_, _10405_, _10401_);
  or _55115_ (_10407_, _10406_, _34772_);
  and _55116_ (_10408_, _10407_, _34719_);
  and _55117_ (_10409_, _10408_, _10397_);
  or _55118_ (_10410_, _10409_, _10387_);
  and _55119_ (_10411_, _10410_, _34700_);
  or _55120_ (_10412_, _10411_, _10365_);
  and _55121_ (_10413_, _10412_, _34840_);
  or _55122_ (_10414_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or _55123_ (_10415_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and _55124_ (_10416_, _10415_, _10414_);
  and _55125_ (_10417_, _10416_, _34581_);
  or _55126_ (_10418_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or _55127_ (_10419_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  and _55128_ (_10420_, _10419_, _10418_);
  and _55129_ (_10421_, _10420_, _34796_);
  or _55130_ (_10422_, _10421_, _10417_);
  and _55131_ (_10423_, _10422_, _34790_);
  or _55132_ (_10424_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or _55133_ (_10425_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and _55134_ (_10426_, _10425_, _10424_);
  and _55135_ (_10427_, _10426_, _34581_);
  or _55136_ (_10428_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or _55137_ (_10429_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and _55138_ (_10430_, _10429_, _10428_);
  and _55139_ (_10431_, _10430_, _34796_);
  or _55140_ (_10432_, _10431_, _10427_);
  and _55141_ (_10433_, _10432_, _34772_);
  or _55142_ (_10434_, _10433_, _10423_);
  and _55143_ (_10435_, _10434_, _34719_);
  and _55144_ (_10436_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and _55145_ (_10437_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or _55146_ (_10438_, _10437_, _10436_);
  and _55147_ (_10439_, _10438_, _34581_);
  and _55148_ (_10440_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and _55149_ (_10441_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or _55150_ (_10442_, _10441_, _10440_);
  and _55151_ (_10443_, _10442_, _34796_);
  or _55152_ (_10444_, _10443_, _10439_);
  and _55153_ (_10445_, _10444_, _34790_);
  and _55154_ (_10446_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and _55155_ (_10447_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or _55156_ (_10448_, _10447_, _10446_);
  and _55157_ (_10449_, _10448_, _34581_);
  and _55158_ (_10450_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  and _55159_ (_10451_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or _55160_ (_10452_, _10451_, _10450_);
  and _55161_ (_10453_, _10452_, _34796_);
  or _55162_ (_10454_, _10453_, _10449_);
  and _55163_ (_10455_, _10454_, _34772_);
  or _55164_ (_10456_, _10455_, _10445_);
  and _55165_ (_10457_, _10456_, _34803_);
  or _55166_ (_10458_, _10457_, _10435_);
  and _55167_ (_10459_, _10458_, _34700_);
  or _55168_ (_10460_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or _55169_ (_10461_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and _55170_ (_10462_, _10461_, _34796_);
  and _55171_ (_10463_, _10462_, _10460_);
  or _55172_ (_10464_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or _55173_ (_10465_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and _55174_ (_10466_, _10465_, _34581_);
  and _55175_ (_10467_, _10466_, _10464_);
  or _55176_ (_10468_, _10467_, _10463_);
  and _55177_ (_10469_, _10468_, _34790_);
  or _55178_ (_10470_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or _55179_ (_10471_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and _55180_ (_10472_, _10471_, _34796_);
  and _55181_ (_10473_, _10472_, _10470_);
  or _55182_ (_10474_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or _55183_ (_10475_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and _55184_ (_10476_, _10475_, _34581_);
  and _55185_ (_10477_, _10476_, _10474_);
  or _55186_ (_10478_, _10477_, _10473_);
  and _55187_ (_10479_, _10478_, _34772_);
  or _55188_ (_10480_, _10479_, _10469_);
  and _55189_ (_10481_, _10480_, _34719_);
  and _55190_ (_10482_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and _55191_ (_10483_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or _55192_ (_10484_, _10483_, _10482_);
  and _55193_ (_10485_, _10484_, _34581_);
  and _55194_ (_10486_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and _55195_ (_10487_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or _55196_ (_10488_, _10487_, _10486_);
  and _55197_ (_10489_, _10488_, _34796_);
  or _55198_ (_10490_, _10489_, _10485_);
  and _55199_ (_10491_, _10490_, _34790_);
  and _55200_ (_10492_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and _55201_ (_10493_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or _55202_ (_10494_, _10493_, _10492_);
  and _55203_ (_10495_, _10494_, _34581_);
  and _55204_ (_10496_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and _55205_ (_10497_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or _55206_ (_10498_, _10497_, _10496_);
  and _55207_ (_10499_, _10498_, _34796_);
  or _55208_ (_10500_, _10499_, _10495_);
  and _55209_ (_10501_, _10500_, _34772_);
  or _55210_ (_10502_, _10501_, _10491_);
  and _55211_ (_10503_, _10502_, _34803_);
  or _55212_ (_10504_, _10503_, _10481_);
  and _55213_ (_10505_, _10504_, _34789_);
  or _55214_ (_10506_, _10505_, _10459_);
  and _55215_ (_10507_, _10506_, _34638_);
  or _55216_ (_10508_, _10507_, _10413_);
  or _55217_ (_10509_, _10508_, _34985_);
  and _55218_ (_10510_, _10509_, _10319_);
  or _55219_ (_10511_, _10510_, _34346_);
  and _55220_ (_10512_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and _55221_ (_10513_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or _55222_ (_10514_, _10513_, _10512_);
  and _55223_ (_10515_, _10514_, _34581_);
  and _55224_ (_10516_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and _55225_ (_10517_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or _55226_ (_10518_, _10517_, _10516_);
  and _55227_ (_10519_, _10518_, _34796_);
  or _55228_ (_10520_, _10519_, _10515_);
  or _55229_ (_10521_, _10520_, _34790_);
  and _55230_ (_10522_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and _55231_ (_10523_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or _55232_ (_10524_, _10523_, _10522_);
  and _55233_ (_10525_, _10524_, _34581_);
  and _55234_ (_10526_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and _55235_ (_10527_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or _55236_ (_10528_, _10527_, _10526_);
  and _55237_ (_10529_, _10528_, _34796_);
  or _55238_ (_10530_, _10529_, _10525_);
  or _55239_ (_10531_, _10530_, _34772_);
  and _55240_ (_10532_, _10531_, _34803_);
  and _55241_ (_10533_, _10532_, _10521_);
  or _55242_ (_10534_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or _55243_ (_10535_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and _55244_ (_10536_, _10535_, _10534_);
  and _55245_ (_10537_, _10536_, _34581_);
  or _55246_ (_10538_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or _55247_ (_10539_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and _55248_ (_10540_, _10539_, _10538_);
  and _55249_ (_10541_, _10540_, _34796_);
  or _55250_ (_10542_, _10541_, _10537_);
  or _55251_ (_10543_, _10542_, _34790_);
  or _55252_ (_10544_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or _55253_ (_10545_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and _55254_ (_10546_, _10545_, _10544_);
  and _55255_ (_10547_, _10546_, _34581_);
  or _55256_ (_10548_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or _55257_ (_10549_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and _55258_ (_10550_, _10549_, _10548_);
  and _55259_ (_10551_, _10550_, _34796_);
  or _55260_ (_10552_, _10551_, _10547_);
  or _55261_ (_10553_, _10552_, _34772_);
  and _55262_ (_10554_, _10553_, _34719_);
  and _55263_ (_10555_, _10554_, _10543_);
  or _55264_ (_10556_, _10555_, _10533_);
  and _55265_ (_10557_, _10556_, _34700_);
  and _55266_ (_10558_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and _55267_ (_10559_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or _55268_ (_10560_, _10559_, _10558_);
  and _55269_ (_10561_, _10560_, _34581_);
  and _55270_ (_10562_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and _55271_ (_10563_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or _55272_ (_10564_, _10563_, _10562_);
  and _55273_ (_10565_, _10564_, _34796_);
  or _55274_ (_10566_, _10565_, _10561_);
  or _55275_ (_10567_, _10566_, _34790_);
  and _55276_ (_10568_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and _55277_ (_10569_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or _55278_ (_10570_, _10569_, _10568_);
  and _55279_ (_10571_, _10570_, _34581_);
  and _55280_ (_10572_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and _55281_ (_10573_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or _55282_ (_10574_, _10573_, _10572_);
  and _55283_ (_10575_, _10574_, _34796_);
  or _55284_ (_10576_, _10575_, _10571_);
  or _55285_ (_10577_, _10576_, _34772_);
  and _55286_ (_10578_, _10577_, _34803_);
  and _55287_ (_10579_, _10578_, _10567_);
  or _55288_ (_10580_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or _55289_ (_10581_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and _55290_ (_10582_, _10581_, _34796_);
  and _55291_ (_10583_, _10582_, _10580_);
  or _55292_ (_10584_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or _55293_ (_10585_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and _55294_ (_10586_, _10585_, _34581_);
  and _55295_ (_10587_, _10586_, _10584_);
  or _55296_ (_10588_, _10587_, _10583_);
  or _55297_ (_10589_, _10588_, _34790_);
  or _55298_ (_10590_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or _55299_ (_10591_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and _55300_ (_10592_, _10591_, _34796_);
  and _55301_ (_10593_, _10592_, _10590_);
  or _55302_ (_10594_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or _55303_ (_10595_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and _55304_ (_10596_, _10595_, _34581_);
  and _55305_ (_10597_, _10596_, _10594_);
  or _55306_ (_10598_, _10597_, _10593_);
  or _55307_ (_10599_, _10598_, _34772_);
  and _55308_ (_10600_, _10599_, _34719_);
  and _55309_ (_10601_, _10600_, _10589_);
  or _55310_ (_10602_, _10601_, _10579_);
  and _55311_ (_10603_, _10602_, _34789_);
  or _55312_ (_10604_, _10603_, _10557_);
  and _55313_ (_10605_, _10604_, _34840_);
  and _55314_ (_10606_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and _55315_ (_10607_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or _55316_ (_10608_, _10607_, _10606_);
  and _55317_ (_10609_, _10608_, _34581_);
  and _55318_ (_10610_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and _55319_ (_10611_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or _55320_ (_10612_, _10611_, _10610_);
  and _55321_ (_10613_, _10612_, _34796_);
  or _55322_ (_10614_, _10613_, _10609_);
  and _55323_ (_10615_, _10614_, _34772_);
  and _55324_ (_10616_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and _55325_ (_10617_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or _55326_ (_10618_, _10617_, _10616_);
  and _55327_ (_10619_, _10618_, _34581_);
  and _55328_ (_10620_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and _55329_ (_10621_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or _55330_ (_10622_, _10621_, _10620_);
  and _55331_ (_10623_, _10622_, _34796_);
  or _55332_ (_10624_, _10623_, _10619_);
  and _55333_ (_10625_, _10624_, _34790_);
  or _55334_ (_10626_, _10625_, _10615_);
  and _55335_ (_10627_, _10626_, _34803_);
  or _55336_ (_10628_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or _55337_ (_10629_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and _55338_ (_10630_, _10629_, _34796_);
  and _55339_ (_10631_, _10630_, _10628_);
  or _55340_ (_10632_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or _55341_ (_10633_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and _55342_ (_10634_, _10633_, _34581_);
  and _55343_ (_10635_, _10634_, _10632_);
  or _55344_ (_10636_, _10635_, _10631_);
  and _55345_ (_10637_, _10636_, _34772_);
  or _55346_ (_10638_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or _55347_ (_10639_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and _55348_ (_10640_, _10639_, _34796_);
  and _55349_ (_10641_, _10640_, _10638_);
  or _55350_ (_10642_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or _55351_ (_10643_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and _55352_ (_10644_, _10643_, _34581_);
  and _55353_ (_10645_, _10644_, _10642_);
  or _55354_ (_10646_, _10645_, _10641_);
  and _55355_ (_10647_, _10646_, _34790_);
  or _55356_ (_10648_, _10647_, _10637_);
  and _55357_ (_10649_, _10648_, _34719_);
  or _55358_ (_10650_, _10649_, _10627_);
  and _55359_ (_10651_, _10650_, _34789_);
  and _55360_ (_10652_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and _55361_ (_10653_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or _55362_ (_10654_, _10653_, _10652_);
  and _55363_ (_10655_, _10654_, _34581_);
  and _55364_ (_10656_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and _55365_ (_10657_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or _55366_ (_10658_, _10657_, _10656_);
  and _55367_ (_10659_, _10658_, _34796_);
  or _55368_ (_10660_, _10659_, _10655_);
  and _55369_ (_10661_, _10660_, _34772_);
  and _55370_ (_10662_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and _55371_ (_10663_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or _55372_ (_10664_, _10663_, _10662_);
  and _55373_ (_10665_, _10664_, _34581_);
  and _55374_ (_10666_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and _55375_ (_10667_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or _55376_ (_10668_, _10667_, _10666_);
  and _55377_ (_10669_, _10668_, _34796_);
  or _55378_ (_10670_, _10669_, _10665_);
  and _55379_ (_10671_, _10670_, _34790_);
  or _55380_ (_10672_, _10671_, _10661_);
  and _55381_ (_10673_, _10672_, _34803_);
  or _55382_ (_10674_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or _55383_ (_10675_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and _55384_ (_10676_, _10675_, _10674_);
  and _55385_ (_10677_, _10676_, _34581_);
  or _55386_ (_10678_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or _55387_ (_10679_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and _55388_ (_10680_, _10679_, _10678_);
  and _55389_ (_10681_, _10680_, _34796_);
  or _55390_ (_10682_, _10681_, _10677_);
  and _55391_ (_10683_, _10682_, _34772_);
  or _55392_ (_10684_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or _55393_ (_10685_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and _55394_ (_10686_, _10685_, _10684_);
  and _55395_ (_10687_, _10686_, _34581_);
  or _55396_ (_10688_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or _55397_ (_10689_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and _55398_ (_10690_, _10689_, _10688_);
  and _55399_ (_10691_, _10690_, _34796_);
  or _55400_ (_10692_, _10691_, _10687_);
  and _55401_ (_10693_, _10692_, _34790_);
  or _55402_ (_10694_, _10693_, _10683_);
  and _55403_ (_10695_, _10694_, _34719_);
  or _55404_ (_10696_, _10695_, _10673_);
  and _55405_ (_10697_, _10696_, _34700_);
  or _55406_ (_10698_, _10697_, _10651_);
  and _55407_ (_10699_, _10698_, _34638_);
  or _55408_ (_10700_, _10699_, _10605_);
  or _55409_ (_10701_, _10700_, _34692_);
  and _55410_ (_10702_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and _55411_ (_10703_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or _55412_ (_10704_, _10703_, _10702_);
  and _55413_ (_10705_, _10704_, _34581_);
  and _55414_ (_10706_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and _55415_ (_10707_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or _55416_ (_10708_, _10707_, _10706_);
  and _55417_ (_10709_, _10708_, _34796_);
  or _55418_ (_10710_, _10709_, _10705_);
  or _55419_ (_10711_, _10710_, _34790_);
  and _55420_ (_10712_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and _55421_ (_10713_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or _55422_ (_10714_, _10713_, _10712_);
  and _55423_ (_10715_, _10714_, _34581_);
  and _55424_ (_10716_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and _55425_ (_10717_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or _55426_ (_10718_, _10717_, _10716_);
  and _55427_ (_10719_, _10718_, _34796_);
  or _55428_ (_10720_, _10719_, _10715_);
  or _55429_ (_10721_, _10720_, _34772_);
  and _55430_ (_10722_, _10721_, _34803_);
  and _55431_ (_10723_, _10722_, _10711_);
  or _55432_ (_10724_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or _55433_ (_10725_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and _55434_ (_10726_, _10725_, _34796_);
  and _55435_ (_10727_, _10726_, _10724_);
  or _55436_ (_10728_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or _55437_ (_10729_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and _55438_ (_10730_, _10729_, _34581_);
  and _55439_ (_10731_, _10730_, _10728_);
  or _55440_ (_10732_, _10731_, _10727_);
  or _55441_ (_10733_, _10732_, _34790_);
  or _55442_ (_10734_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or _55443_ (_10735_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and _55444_ (_10736_, _10735_, _34796_);
  and _55445_ (_10737_, _10736_, _10734_);
  or _55446_ (_10738_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or _55447_ (_10739_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and _55448_ (_10740_, _10739_, _34581_);
  and _55449_ (_10741_, _10740_, _10738_);
  or _55450_ (_10742_, _10741_, _10737_);
  or _55451_ (_10743_, _10742_, _34772_);
  and _55452_ (_10744_, _10743_, _34719_);
  and _55453_ (_10745_, _10744_, _10733_);
  or _55454_ (_10746_, _10745_, _10723_);
  and _55455_ (_10747_, _10746_, _34789_);
  and _55456_ (_10748_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and _55457_ (_10749_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or _55458_ (_10750_, _10749_, _10748_);
  and _55459_ (_10751_, _10750_, _34581_);
  and _55460_ (_10752_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and _55461_ (_10753_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or _55462_ (_10754_, _10753_, _10752_);
  and _55463_ (_10755_, _10754_, _34796_);
  or _55464_ (_10756_, _10755_, _10751_);
  or _55465_ (_10757_, _10756_, _34790_);
  and _55466_ (_10758_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and _55467_ (_10759_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or _55468_ (_10760_, _10759_, _10758_);
  and _55469_ (_10761_, _10760_, _34581_);
  and _55470_ (_10762_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and _55471_ (_10763_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or _55472_ (_10764_, _10763_, _10762_);
  and _55473_ (_10765_, _10764_, _34796_);
  or _55474_ (_10766_, _10765_, _10761_);
  or _55475_ (_10767_, _10766_, _34772_);
  and _55476_ (_10768_, _10767_, _34803_);
  and _55477_ (_10769_, _10768_, _10757_);
  or _55478_ (_10770_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or _55479_ (_10771_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and _55480_ (_10772_, _10771_, _10770_);
  and _55481_ (_10773_, _10772_, _34581_);
  or _55482_ (_10774_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or _55483_ (_10775_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and _55484_ (_10776_, _10775_, _10774_);
  and _55485_ (_10777_, _10776_, _34796_);
  or _55486_ (_10778_, _10777_, _10773_);
  or _55487_ (_10779_, _10778_, _34790_);
  or _55488_ (_10780_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or _55489_ (_10781_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and _55490_ (_10782_, _10781_, _10780_);
  and _55491_ (_10783_, _10782_, _34581_);
  or _55492_ (_10784_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or _55493_ (_10785_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and _55494_ (_10786_, _10785_, _10784_);
  and _55495_ (_10787_, _10786_, _34796_);
  or _55496_ (_10788_, _10787_, _10783_);
  or _55497_ (_10789_, _10788_, _34772_);
  and _55498_ (_10790_, _10789_, _34719_);
  and _55499_ (_10791_, _10790_, _10779_);
  or _55500_ (_10792_, _10791_, _10769_);
  and _55501_ (_10793_, _10792_, _34700_);
  or _55502_ (_10794_, _10793_, _10747_);
  and _55503_ (_10795_, _10794_, _34840_);
  or _55504_ (_10796_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or _55505_ (_10797_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and _55506_ (_10798_, _10797_, _10796_);
  and _55507_ (_10799_, _10798_, _34581_);
  or _55508_ (_10800_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or _55509_ (_10801_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and _55510_ (_10802_, _10801_, _10800_);
  and _55511_ (_10803_, _10802_, _34796_);
  or _55512_ (_10804_, _10803_, _10799_);
  and _55513_ (_10805_, _10804_, _34790_);
  or _55514_ (_10806_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or _55515_ (_10807_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and _55516_ (_10808_, _10807_, _10806_);
  and _55517_ (_10809_, _10808_, _34581_);
  or _55518_ (_10810_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or _55519_ (_10811_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and _55520_ (_10812_, _10811_, _10810_);
  and _55521_ (_10813_, _10812_, _34796_);
  or _55522_ (_10814_, _10813_, _10809_);
  and _55523_ (_10815_, _10814_, _34772_);
  or _55524_ (_10816_, _10815_, _10805_);
  and _55525_ (_10817_, _10816_, _34719_);
  and _55526_ (_10818_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and _55527_ (_10819_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or _55528_ (_10820_, _10819_, _10818_);
  and _55529_ (_10821_, _10820_, _34581_);
  and _55530_ (_10822_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and _55531_ (_10823_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or _55532_ (_10824_, _10823_, _10822_);
  and _55533_ (_10825_, _10824_, _34796_);
  or _55534_ (_10826_, _10825_, _10821_);
  and _55535_ (_10827_, _10826_, _34790_);
  and _55536_ (_10828_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and _55537_ (_10829_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or _55538_ (_10830_, _10829_, _10828_);
  and _55539_ (_10831_, _10830_, _34581_);
  and _55540_ (_10832_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and _55541_ (_10833_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or _55542_ (_10834_, _10833_, _10832_);
  and _55543_ (_10835_, _10834_, _34796_);
  or _55544_ (_10836_, _10835_, _10831_);
  and _55545_ (_10837_, _10836_, _34772_);
  or _55546_ (_10838_, _10837_, _10827_);
  and _55547_ (_10839_, _10838_, _34803_);
  or _55548_ (_10840_, _10839_, _10817_);
  and _55549_ (_10841_, _10840_, _34700_);
  or _55550_ (_10842_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or _55551_ (_10843_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and _55552_ (_10844_, _10843_, _34796_);
  and _55553_ (_10845_, _10844_, _10842_);
  or _55554_ (_10846_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or _55555_ (_10847_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and _55556_ (_10848_, _10847_, _34581_);
  and _55557_ (_10849_, _10848_, _10846_);
  or _55558_ (_10850_, _10849_, _10845_);
  and _55559_ (_10851_, _10850_, _34790_);
  or _55560_ (_10852_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or _55561_ (_10853_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and _55562_ (_10854_, _10853_, _34796_);
  and _55563_ (_10855_, _10854_, _10852_);
  or _55564_ (_10856_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or _55565_ (_10857_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and _55566_ (_10858_, _10857_, _34581_);
  and _55567_ (_10859_, _10858_, _10856_);
  or _55568_ (_10860_, _10859_, _10855_);
  and _55569_ (_10861_, _10860_, _34772_);
  or _55570_ (_10862_, _10861_, _10851_);
  and _55571_ (_10863_, _10862_, _34719_);
  and _55572_ (_10864_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and _55573_ (_10865_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or _55574_ (_10866_, _10865_, _10864_);
  and _55575_ (_10867_, _10866_, _34581_);
  and _55576_ (_10868_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and _55577_ (_10869_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or _55578_ (_10870_, _10869_, _10868_);
  and _55579_ (_10871_, _10870_, _34796_);
  or _55580_ (_10872_, _10871_, _10867_);
  and _55581_ (_10873_, _10872_, _34790_);
  and _55582_ (_10874_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and _55583_ (_10875_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or _55584_ (_10876_, _10875_, _10874_);
  and _55585_ (_10877_, _10876_, _34581_);
  and _55586_ (_10878_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and _55587_ (_10879_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or _55588_ (_10880_, _10879_, _10878_);
  and _55589_ (_10881_, _10880_, _34796_);
  or _55590_ (_10882_, _10881_, _10877_);
  and _55591_ (_10883_, _10882_, _34772_);
  or _55592_ (_10884_, _10883_, _10873_);
  and _55593_ (_10885_, _10884_, _34803_);
  or _55594_ (_10886_, _10885_, _10863_);
  and _55595_ (_10887_, _10886_, _34789_);
  or _55596_ (_10888_, _10887_, _10841_);
  and _55597_ (_10889_, _10888_, _34638_);
  or _55598_ (_10890_, _10889_, _10795_);
  or _55599_ (_10891_, _10890_, _34985_);
  and _55600_ (_10892_, _10891_, _10701_);
  or _55601_ (_10893_, _10892_, _35178_);
  and _55602_ (_10894_, _10893_, _10511_);
  or _55603_ (_10895_, _10894_, _34788_);
  or _55604_ (_10896_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and _55605_ (_10897_, _10896_, _38997_);
  and _55606_ (_38984_[6], _10897_, _10895_);
  nor _55607_ (_10898_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _55608_ (_39040_, _10898_, rst);
  and _55609_ (_10899_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _55610_ (_10900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor _55611_ (_10901_, _10898_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and _55612_ (_10902_, _10901_, _10900_);
  not _55613_ (_10903_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _55614_ (_10904_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _10903_);
  or _55615_ (_10905_, _10904_, _10902_);
  nor _55616_ (_10906_, _10905_, _10899_);
  or _55617_ (_10907_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _55618_ (_10908_, _10907_, _38997_);
  nor _55619_ (_39041_, _10908_, _10906_);
  nor _55620_ (_10909_, _10906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _55621_ (_10910_, _10909_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _55622_ (_10911_, _10909_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _55623_ (_10912_, _10911_, _38997_);
  and _55624_ (_39042_, _10912_, _10910_);
  not _55625_ (_10913_, rxd_i);
  and _55626_ (_10914_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _10913_);
  nor _55627_ (_10915_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _55628_ (_10916_, _10915_);
  and _55629_ (_10917_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and _55630_ (_10918_, _10917_, _10916_);
  and _55631_ (_10919_, _10918_, _10914_);
  not _55632_ (_10920_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _55633_ (_10921_, _10920_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _55634_ (_10922_, _10921_, _10915_);
  or _55635_ (_10923_, _10922_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or _55636_ (_10924_, _10923_, _10919_);
  and _55637_ (_10925_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _38997_);
  and _55638_ (_39043_, _10925_, _10924_);
  and _55639_ (_10926_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _55640_ (_10927_, _10926_, _10916_);
  nor _55641_ (_10928_, _10915_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _55642_ (_10929_, _10928_, _10920_);
  nor _55643_ (_10930_, _10929_, _10927_);
  not _55644_ (_10931_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _55645_ (_10932_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _10931_);
  not _55646_ (_10933_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _55647_ (_10934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _10933_);
  and _55648_ (_10935_, _10934_, _10932_);
  not _55649_ (_10936_, _10935_);
  or _55650_ (_10937_, _10936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and _55651_ (_10938_, _10935_, _10927_);
  and _55652_ (_10939_, _10927_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _55653_ (_10940_, _10939_, _10938_);
  and _55654_ (_10941_, _10940_, _10937_);
  or _55655_ (_10942_, _10941_, _10930_);
  and _55656_ (_10943_, _10915_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _55657_ (_10944_, _10943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  not _55658_ (_10945_, _10944_);
  or _55659_ (_10946_, _10945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand _55660_ (_10947_, _10946_, _10942_);
  nand _55661_ (_39044_, _10947_, _10925_);
  not _55662_ (_10948_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not _55663_ (_10949_, _10927_);
  nor _55664_ (_10950_, _10920_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _55665_ (_10951_, _10950_);
  not _55666_ (_10952_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _55667_ (_10953_, _10915_, _10952_);
  and _55668_ (_10954_, _10953_, _10951_);
  and _55669_ (_10955_, _10954_, _10949_);
  nor _55670_ (_10956_, _10955_, _10948_);
  and _55671_ (_10957_, _10955_, rxd_i);
  or _55672_ (_10958_, _10957_, rst);
  or _55673_ (_39045_, _10958_, _10956_);
  nor _55674_ (_10959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _55675_ (_10960_, _10959_, _10932_);
  and _55676_ (_10961_, _10960_, _10939_);
  nand _55677_ (_10962_, _10961_, _10913_);
  or _55678_ (_10963_, _10961_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _55679_ (_10964_, _10963_, _38997_);
  and _55680_ (_39046_[1], _10964_, _10962_);
  and _55681_ (_10965_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _55682_ (_10966_, _10965_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _55683_ (_10967_, _10966_, _10931_);
  and _55684_ (_10968_, _10967_, _10939_);
  and _55685_ (_10969_, _10918_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _55686_ (_10970_, _10969_, _10939_);
  nor _55687_ (_10971_, _10966_, _10949_);
  or _55688_ (_10972_, _10971_, _10970_);
  and _55689_ (_10973_, _10972_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _55690_ (_10974_, _10973_, _10968_);
  and _55691_ (_39047_[3], _10974_, _38997_);
  and _55692_ (_10975_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _38997_);
  nand _55693_ (_10976_, _10975_, _10952_);
  nand _55694_ (_10977_, _10925_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand _55695_ (_39048_[7], _10977_, _10976_);
  and _55696_ (_10978_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _10952_);
  not _55697_ (_10979_, _10918_);
  not _55698_ (_10980_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand _55699_ (_10981_, _10922_, _10980_);
  and _55700_ (_10982_, _10981_, _10979_);
  nand _55701_ (_10983_, _10982_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand _55702_ (_10984_, _10983_, _10949_);
  or _55703_ (_10985_, _10935_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor _55704_ (_10986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _55705_ (_10987_, _10986_, _10938_);
  and _55706_ (_10988_, _10987_, _10985_);
  and _55707_ (_10989_, _10988_, _10984_);
  or _55708_ (_10990_, _10989_, _10944_);
  nand _55709_ (_10991_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _55710_ (_10992_, _10991_, _10927_);
  or _55711_ (_10993_, _10992_, _10936_);
  and _55712_ (_10994_, _10993_, _10945_);
  or _55713_ (_10995_, _10994_, rxd_i);
  and _55714_ (_10996_, _10995_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _55715_ (_10997_, _10996_, _10990_);
  or _55716_ (_10998_, _10997_, _10978_);
  and _55717_ (_39049_[11], _10998_, _38997_);
  and _55718_ (_10999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _55719_ (_11000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _55720_ (_11001_, _10901_, _11000_);
  or _55721_ (_11002_, _11001_, _10904_);
  nor _55722_ (_11003_, _11002_, _10999_);
  or _55723_ (_11004_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _55724_ (_11005_, _11004_, _38997_);
  nor _55725_ (_39050_, _11005_, _11003_);
  nor _55726_ (_11006_, _11003_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _55727_ (_11007_, _11006_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _55728_ (_11008_, _11006_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _55729_ (_11009_, _11008_, _38997_);
  and _55730_ (_39051_, _11009_, _11007_);
  not _55731_ (_11010_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and _55732_ (_11011_, _34233_, _33632_);
  and _55733_ (_11012_, _34254_, _33662_);
  and _55734_ (_11013_, _11012_, _11011_);
  and _55735_ (_11014_, _11013_, _38997_);
  nand _55736_ (_11015_, _11014_, _11010_);
  and _55737_ (_11016_, _10943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  not _55738_ (_11017_, _11016_);
  nor _55739_ (_11018_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not _55740_ (_11019_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _55741_ (_11020_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _55742_ (_11021_, _11020_, _11019_);
  and _55743_ (_11022_, _11021_, _11018_);
  not _55744_ (_11023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _55745_ (_11024_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _55746_ (_11025_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _55747_ (_11026_, _11025_, _11024_);
  and _55748_ (_11027_, _11026_, _11023_);
  and _55749_ (_11028_, _11027_, _11022_);
  or _55750_ (_11029_, _11028_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  not _55751_ (_11030_, _11028_);
  or _55752_ (_11031_, _11030_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and _55753_ (_11032_, _11031_, _11029_);
  or _55754_ (_11033_, _11032_, _11017_);
  nor _55755_ (_11034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _55756_ (_11035_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _55757_ (_11036_, _11035_, _11034_);
  and _55758_ (_11037_, _10916_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _55759_ (_11038_, _11037_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _55760_ (_11039_, _11038_, _11036_);
  not _55761_ (_11040_, _11039_);
  or _55762_ (_11041_, _11040_, _11029_);
  and _55763_ (_11042_, _11036_, _11037_);
  not _55764_ (_11043_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or _55765_ (_11044_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _11043_);
  or _55766_ (_11045_, _11044_, _11042_);
  or _55767_ (_11046_, _11045_, _11016_);
  and _55768_ (_11047_, _11046_, _11041_);
  nand _55769_ (_11048_, _11047_, _11033_);
  nor _55770_ (_11049_, _11013_, rst);
  nand _55771_ (_11050_, _11049_, _11048_);
  and _55772_ (_39052_, _11050_, _11015_);
  nor _55773_ (_11051_, _11030_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand _55774_ (_11052_, _11042_, _11051_);
  and _55775_ (_11053_, _11028_, _11016_);
  or _55776_ (_11054_, _11043_, rst);
  nor _55777_ (_11055_, _11054_, _11053_);
  and _55778_ (_11056_, _11055_, _11052_);
  or _55779_ (_39053_, _11056_, _11014_);
  or _55780_ (_11057_, _11040_, _11051_);
  or _55781_ (_11058_, _11042_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _55782_ (_11059_, _10943_, _11043_);
  and _55783_ (_11060_, _11059_, _11058_);
  and _55784_ (_11061_, _11060_, _11057_);
  or _55785_ (_11062_, _11061_, _11053_);
  and _55786_ (_39054_, _11062_, _11049_);
  and _55787_ (_11063_, _11038_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _55788_ (_11064_, _11063_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _55789_ (_11065_, _11064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or _55790_ (_11066_, _11065_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand _55791_ (_11067_, _11065_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _55792_ (_11068_, _11067_, _11066_);
  and _55793_ (_39055_[3], _11068_, _11049_);
  nor _55794_ (_11069_, _11039_, _11016_);
  and _55795_ (_11070_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _55796_ (_11071_, _11070_, _11049_);
  and _55797_ (_11072_, _11014_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _55798_ (_39056_[10], _11072_, _11071_);
  not _55799_ (_11073_, _33644_);
  nor _55800_ (_11074_, _33571_, _33558_);
  and _55801_ (_11075_, _11074_, _11073_);
  and _55802_ (_11076_, _11075_, _33663_);
  and _55803_ (_11077_, _11076_, _33633_);
  nand _55804_ (_11078_, _11077_, _34221_);
  or _55805_ (_11079_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _55806_ (_11080_, _11079_, _38997_);
  and _55807_ (_39057_[7], _11080_, _11078_);
  and _55808_ (_11081_, _33630_, _33591_);
  nor _55809_ (_11082_, _33657_, _33604_);
  and _55810_ (_11083_, _33661_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _55811_ (_11084_, _11083_, _34706_);
  and _55812_ (_11085_, _11084_, _11082_);
  and _55813_ (_11086_, _11085_, _11081_);
  and _55814_ (_11087_, _11086_, _11075_);
  or _55815_ (_11088_, _11087_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  not _55816_ (_11089_, _33662_);
  nor _55817_ (_11090_, _11089_, _33657_);
  and _55818_ (_11091_, _11090_, _34229_);
  and _55819_ (_11092_, _11091_, _11011_);
  not _55820_ (_11093_, _11092_);
  and _55821_ (_11094_, _11093_, _11088_);
  nand _55822_ (_11095_, _11087_, _35722_);
  and _55823_ (_11096_, _11095_, _11094_);
  nor _55824_ (_11097_, _11093_, _34221_);
  or _55825_ (_11098_, _11097_, _11096_);
  and _55826_ (_39058_[7], _11098_, _38997_);
  nor _55827_ (_11099_, _10944_, _10938_);
  not _55828_ (_11100_, _11099_);
  nor _55829_ (_11101_, _10982_, _10927_);
  nor _55830_ (_11102_, _11101_, _11100_);
  nor _55831_ (_11103_, _11102_, _10952_);
  or _55832_ (_11104_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _55833_ (_11105_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _10952_);
  or _55834_ (_11106_, _11105_, _11099_);
  and _55835_ (_11107_, _11106_, _38997_);
  and _55836_ (_39049_[0], _11107_, _11104_);
  or _55837_ (_11108_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _55838_ (_11109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _10952_);
  or _55839_ (_11110_, _11109_, _11099_);
  and _55840_ (_11111_, _11110_, _38997_);
  and _55841_ (_39049_[1], _11111_, _11108_);
  or _55842_ (_11112_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _55843_ (_11113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _10952_);
  or _55844_ (_11114_, _11113_, _11099_);
  and _55845_ (_11115_, _11114_, _38997_);
  and _55846_ (_39049_[2], _11115_, _11112_);
  or _55847_ (_11116_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _55848_ (_11117_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _10952_);
  or _55849_ (_11118_, _11117_, _11099_);
  and _55850_ (_11119_, _11118_, _38997_);
  and _55851_ (_39049_[3], _11119_, _11116_);
  or _55852_ (_11120_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _55853_ (_11121_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _10952_);
  or _55854_ (_11122_, _11121_, _11099_);
  and _55855_ (_11123_, _11122_, _38997_);
  and _55856_ (_39049_[4], _11123_, _11120_);
  or _55857_ (_11124_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _55858_ (_11125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _10952_);
  or _55859_ (_11126_, _11125_, _11099_);
  and _55860_ (_11127_, _11126_, _38997_);
  and _55861_ (_39049_[5], _11127_, _11124_);
  or _55862_ (_11128_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _55863_ (_11129_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _10952_);
  or _55864_ (_11130_, _11129_, _11099_);
  and _55865_ (_11131_, _11130_, _38997_);
  and _55866_ (_39049_[6], _11131_, _11128_);
  or _55867_ (_11132_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _55868_ (_11133_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _10952_);
  or _55869_ (_11134_, _11133_, _11099_);
  and _55870_ (_11135_, _11134_, _38997_);
  and _55871_ (_39049_[7], _11135_, _11132_);
  nor _55872_ (_11136_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and _55873_ (_11137_, _11136_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _55874_ (_11138_, _10936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or _55875_ (_11139_, _10935_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _55876_ (_11140_, _11139_, _10927_);
  and _55877_ (_11141_, _11140_, _11138_);
  or _55878_ (_11142_, _10918_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _55879_ (_11143_, _11142_, _10981_);
  and _55880_ (_11144_, _11143_, _10949_);
  or _55881_ (_11145_, _11144_, _11141_);
  or _55882_ (_11146_, _11145_, _10944_);
  or _55883_ (_11147_, _10945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _55884_ (_11148_, _11147_, _10925_);
  and _55885_ (_11149_, _11148_, _11146_);
  or _55886_ (_39049_[8], _11149_, _11137_);
  and _55887_ (_11150_, _10935_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _55888_ (_11151_, _11150_, _10982_);
  or _55889_ (_11152_, _11151_, _11102_);
  and _55890_ (_11153_, _11152_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _55891_ (_11154_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _10952_);
  nand _55892_ (_11155_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _55893_ (_11156_, _11155_, _11099_);
  or _55894_ (_11157_, _11156_, _11154_);
  or _55895_ (_11158_, _11157_, _11153_);
  and _55896_ (_39049_[9], _11158_, _38997_);
  not _55897_ (_11159_, _11103_);
  and _55898_ (_11160_, _11159_, _10975_);
  or _55899_ (_11161_, _11151_, _11100_);
  and _55900_ (_11162_, _10925_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _55901_ (_11163_, _11162_, _11161_);
  or _55902_ (_39049_[10], _11163_, _11160_);
  or _55903_ (_11164_, _10968_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand _55904_ (_11165_, _10968_, _10913_);
  and _55905_ (_11166_, _11165_, _38997_);
  and _55906_ (_39046_[0], _11166_, _11164_);
  or _55907_ (_11167_, _10970_, _10933_);
  or _55908_ (_11168_, _10939_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _55909_ (_11169_, _11168_, _38997_);
  and _55910_ (_39047_[0], _11169_, _11167_);
  and _55911_ (_11170_, _10970_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _55912_ (_11171_, _10959_, _10965_);
  and _55913_ (_11172_, _11171_, _10939_);
  or _55914_ (_11173_, _11172_, _11170_);
  and _55915_ (_39047_[1], _11173_, _38997_);
  and _55916_ (_11174_, _10972_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _55917_ (_11175_, _10965_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _55918_ (_11176_, _11175_, _10971_);
  or _55919_ (_11177_, _11176_, _11174_);
  and _55920_ (_39047_[2], _11177_, _38997_);
  and _55921_ (_11178_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _10952_);
  and _55922_ (_11179_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _55923_ (_11180_, _11179_, _11178_);
  and _55924_ (_39048_[0], _11180_, _38997_);
  and _55925_ (_11181_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _10952_);
  and _55926_ (_11182_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _55927_ (_11183_, _11182_, _11181_);
  and _55928_ (_39048_[1], _11183_, _38997_);
  and _55929_ (_11184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _10952_);
  and _55930_ (_11185_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _55931_ (_11186_, _11185_, _11184_);
  and _55932_ (_39048_[2], _11186_, _38997_);
  and _55933_ (_11187_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _10952_);
  and _55934_ (_11188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _55935_ (_11189_, _11188_, _11187_);
  and _55936_ (_39048_[3], _11189_, _38997_);
  and _55937_ (_11190_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _10952_);
  and _55938_ (_11191_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _55939_ (_11192_, _11191_, _11190_);
  and _55940_ (_39048_[4], _11192_, _38997_);
  and _55941_ (_11193_, _10925_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _55942_ (_39048_[5], _11193_, _11137_);
  and _55943_ (_11194_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _55944_ (_11195_, _11194_, _11154_);
  and _55945_ (_39048_[6], _11195_, _38997_);
  nor _55946_ (_11196_, _11038_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _55947_ (_11197_, _11196_, _11063_);
  and _55948_ (_39055_[0], _11197_, _11049_);
  nor _55949_ (_11198_, _11063_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _55950_ (_11199_, _11198_, _11064_);
  and _55951_ (_39055_[1], _11199_, _11049_);
  nor _55952_ (_11200_, _11064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _55953_ (_11201_, _11200_, _11065_);
  and _55954_ (_39055_[2], _11201_, _11049_);
  or _55955_ (_11202_, _11039_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _55956_ (_11203_, _11040_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _55957_ (_11204_, _11203_, _11202_);
  and _55958_ (_11205_, _11204_, _11017_);
  and _55959_ (_11206_, _11028_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _55960_ (_11207_, _11206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _55961_ (_11208_, _11207_, _11016_);
  or _55962_ (_11209_, _11208_, _11205_);
  and _55963_ (_11210_, _11209_, _11049_);
  nor _55964_ (_11211_, _10916_, _34148_);
  and _55965_ (_11212_, _11211_, _11014_);
  or _55966_ (_39056_[0], _11212_, _11210_);
  not _55967_ (_11213_, _11069_);
  and _55968_ (_11214_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _55969_ (_11215_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _55970_ (_11216_, _11215_, _11214_);
  and _55971_ (_11217_, _11216_, _11049_);
  or _55972_ (_11218_, _10916_, _34122_);
  nand _55973_ (_11219_, _10916_, _34148_);
  and _55974_ (_11220_, _11219_, _11014_);
  and _55975_ (_11221_, _11220_, _11218_);
  or _55976_ (_39056_[1], _11221_, _11217_);
  nor _55977_ (_11222_, _11069_, _11023_);
  and _55978_ (_11223_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or _55979_ (_11224_, _11223_, _11222_);
  and _55980_ (_11225_, _11224_, _11049_);
  or _55981_ (_11226_, _10916_, _34089_);
  or _55982_ (_11227_, _10915_, _34122_);
  and _55983_ (_11228_, _11227_, _11014_);
  and _55984_ (_11229_, _11228_, _11226_);
  or _55985_ (_39056_[2], _11229_, _11225_);
  nor _55986_ (_11230_, _11069_, _11019_);
  and _55987_ (_11231_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or _55988_ (_11232_, _11231_, _11230_);
  and _55989_ (_11233_, _11232_, _11049_);
  or _55990_ (_11234_, _10915_, _34089_);
  nand _55991_ (_11235_, _10915_, _34052_);
  and _55992_ (_11236_, _11235_, _11014_);
  and _55993_ (_11237_, _11236_, _11234_);
  or _55994_ (_39056_[3], _11237_, _11233_);
  and _55995_ (_11238_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _55996_ (_11239_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  or _55997_ (_11240_, _11239_, _11238_);
  and _55998_ (_11241_, _11240_, _11049_);
  nand _55999_ (_11242_, _10916_, _34052_);
  nand _56000_ (_11243_, _10915_, _34017_);
  and _56001_ (_11244_, _11243_, _11014_);
  and _56002_ (_11245_, _11244_, _11242_);
  or _56003_ (_39056_[4], _11245_, _11241_);
  and _56004_ (_11246_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _56005_ (_11247_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or _56006_ (_11248_, _11247_, _11246_);
  and _56007_ (_11249_, _11248_, _11049_);
  or _56008_ (_11250_, _10916_, _33978_);
  nand _56009_ (_11251_, _10916_, _34017_);
  and _56010_ (_11252_, _11251_, _11014_);
  and _56011_ (_11253_, _11252_, _11250_);
  or _56012_ (_39056_[5], _11253_, _11249_);
  and _56013_ (_11254_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _56014_ (_11255_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or _56015_ (_11256_, _11255_, _11254_);
  and _56016_ (_11257_, _11256_, _11049_);
  or _56017_ (_11258_, _10915_, _33978_);
  or _56018_ (_11259_, _10916_, _33942_);
  and _56019_ (_11260_, _11259_, _11014_);
  and _56020_ (_11261_, _11260_, _11258_);
  or _56021_ (_39056_[6], _11261_, _11257_);
  and _56022_ (_11262_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _56023_ (_11263_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or _56024_ (_11264_, _11263_, _11262_);
  and _56025_ (_11265_, _11264_, _11049_);
  nand _56026_ (_11266_, _10915_, _34221_);
  or _56027_ (_11267_, _10915_, _33942_);
  and _56028_ (_11268_, _11267_, _11014_);
  and _56029_ (_11269_, _11268_, _11266_);
  or _56030_ (_39056_[7], _11269_, _11265_);
  or _56031_ (_11270_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  or _56032_ (_11271_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  and _56033_ (_11272_, _11271_, _38997_);
  and _56034_ (_11273_, _11272_, _11270_);
  or _56035_ (_11274_, _11273_, _11014_);
  and _56036_ (_11275_, _11013_, _10916_);
  nand _56037_ (_11276_, _11275_, _34221_);
  and _56038_ (_39056_[8], _11276_, _11274_);
  and _56039_ (_11277_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _56040_ (_11278_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _56041_ (_11279_, _11278_, _11277_);
  and _56042_ (_11280_, _11279_, _11049_);
  not _56043_ (_11281_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _56044_ (_11282_, _11281_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _56045_ (_11283_, _11282_, _10916_);
  and _56046_ (_11284_, _11283_, _11014_);
  or _56047_ (_39056_[9], _11284_, _11280_);
  nand _56048_ (_11285_, _11077_, _34148_);
  or _56049_ (_11286_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _56050_ (_11287_, _11286_, _38997_);
  and _56051_ (_39057_[0], _11287_, _11285_);
  not _56052_ (_11288_, _11077_);
  or _56053_ (_11289_, _11288_, _34122_);
  or _56054_ (_11290_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _56055_ (_11291_, _11290_, _38997_);
  and _56056_ (_39057_[1], _11291_, _11289_);
  or _56057_ (_11292_, _11288_, _34089_);
  or _56058_ (_11293_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _56059_ (_11294_, _11293_, _38997_);
  and _56060_ (_39057_[2], _11294_, _11292_);
  nand _56061_ (_11295_, _11077_, _34052_);
  or _56062_ (_11296_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _56063_ (_11297_, _11296_, _38997_);
  and _56064_ (_39057_[3], _11297_, _11295_);
  nand _56065_ (_11298_, _11077_, _34017_);
  or _56066_ (_11299_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _56067_ (_11300_, _11299_, _38997_);
  and _56068_ (_39057_[4], _11300_, _11298_);
  or _56069_ (_11301_, _11288_, _33978_);
  or _56070_ (_11302_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _56071_ (_11303_, _11302_, _38997_);
  and _56072_ (_39057_[5], _11303_, _11301_);
  or _56073_ (_11304_, _11288_, _33942_);
  or _56074_ (_11305_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _56075_ (_11306_, _11305_, _38997_);
  and _56076_ (_39057_[6], _11306_, _11304_);
  not _56077_ (_11307_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _56078_ (_11308_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _11307_);
  or _56079_ (_11309_, _11308_, _10915_);
  nor _56080_ (_11310_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _56081_ (_11311_, _11310_, _11309_);
  or _56082_ (_11312_, _11311_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _56083_ (_11313_, _11312_, _11086_);
  not _56084_ (_11314_, _34229_);
  nor _56085_ (_11315_, _35722_, _11314_);
  nand _56086_ (_11316_, _11314_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand _56087_ (_11317_, _11316_, _11086_);
  or _56088_ (_11318_, _11317_, _11315_);
  and _56089_ (_11319_, _11318_, _11313_);
  or _56090_ (_11320_, _11319_, _11092_);
  nand _56091_ (_11321_, _11092_, _34148_);
  and _56092_ (_11322_, _11321_, _38997_);
  and _56093_ (_39058_[0], _11322_, _11320_);
  or _56094_ (_11323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _56095_ (_11324_, _11323_, _11086_);
  not _56096_ (_11325_, _34253_);
  nor _56097_ (_11326_, _35722_, _11325_);
  nand _56098_ (_11327_, _11325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _56099_ (_11328_, _11327_, _11086_);
  or _56100_ (_11329_, _11328_, _11326_);
  and _56101_ (_11330_, _11329_, _11324_);
  or _56102_ (_11331_, _11330_, _11092_);
  or _56103_ (_11332_, _11093_, _34122_);
  and _56104_ (_11333_, _11332_, _38997_);
  and _56105_ (_39058_[1], _11333_, _11331_);
  not _56106_ (_11334_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not _56107_ (_11335_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and _56108_ (_11336_, _10928_, _11335_);
  nor _56109_ (_11337_, _11336_, _11334_);
  and _56110_ (_11338_, _11336_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _56111_ (_11339_, _11338_, _11337_);
  or _56112_ (_11340_, _11339_, _11086_);
  not _56113_ (_11341_, _33571_);
  and _56114_ (_11342_, _11341_, _33558_);
  and _56115_ (_11343_, _11342_, _33644_);
  not _56116_ (_11344_, _11343_);
  nor _56117_ (_11345_, _11344_, _35722_);
  or _56118_ (_11346_, _11343_, _11334_);
  nand _56119_ (_11347_, _11346_, _11086_);
  or _56120_ (_11348_, _11347_, _11345_);
  and _56121_ (_11349_, _11348_, _11340_);
  or _56122_ (_11350_, _11349_, _11092_);
  or _56123_ (_11351_, _11093_, _34089_);
  and _56124_ (_11352_, _11351_, _38997_);
  and _56125_ (_39058_[2], _11352_, _11350_);
  nand _56126_ (_11353_, _11086_, _33644_);
  and _56127_ (_11354_, _11353_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _56128_ (_11355_, _11354_, _11092_);
  and _56129_ (_11356_, _11074_, _33644_);
  and _56130_ (_11357_, _11356_, _35723_);
  or _56131_ (_11358_, _11074_, _11073_);
  not _56132_ (_11359_, _11358_);
  and _56133_ (_11360_, _11359_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _56134_ (_11361_, _11360_, _11357_);
  and _56135_ (_11362_, _11361_, _11086_);
  or _56136_ (_11363_, _11362_, _11355_);
  nand _56137_ (_11364_, _11092_, _34052_);
  and _56138_ (_11365_, _11364_, _38997_);
  and _56139_ (_39058_[3], _11365_, _11363_);
  and _56140_ (_11366_, _11083_, _34251_);
  and _56141_ (_11367_, _11366_, _34227_);
  and _56142_ (_11368_, _11367_, _34706_);
  nand _56143_ (_11369_, _11368_, _11081_);
  and _56144_ (_11370_, _34228_, _11073_);
  nor _56145_ (_11371_, _34228_, _11073_);
  nor _56146_ (_11372_, _11371_, _11370_);
  or _56147_ (_11373_, _11372_, _11369_);
  and _56148_ (_11374_, _11373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _56149_ (_11375_, _11374_, _11092_);
  and _56150_ (_11376_, _11370_, _35723_);
  and _56151_ (_11377_, _11371_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _56152_ (_11378_, _11377_, _11376_);
  and _56153_ (_11379_, _11378_, _11086_);
  or _56154_ (_11380_, _11379_, _11375_);
  nand _56155_ (_11381_, _11092_, _34017_);
  and _56156_ (_11382_, _11381_, _38997_);
  and _56157_ (_39058_[4], _11382_, _11380_);
  and _56158_ (_11383_, _11073_, _33572_);
  and _56159_ (_11384_, _11086_, _11383_);
  or _56160_ (_11385_, _11384_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _56161_ (_11386_, _11385_, _11093_);
  nand _56162_ (_11387_, _11384_, _35722_);
  and _56163_ (_11388_, _11387_, _11386_);
  and _56164_ (_11389_, _11092_, _33978_);
  or _56165_ (_11390_, _11389_, _11388_);
  and _56166_ (_39058_[5], _11390_, _38997_);
  nor _56167_ (_11391_, _33644_, _33571_);
  and _56168_ (_11392_, _11391_, _33558_);
  not _56169_ (_11393_, _11392_);
  or _56170_ (_11394_, _11369_, _11393_);
  and _56171_ (_11395_, _11394_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _56172_ (_11396_, _11395_, _11092_);
  nor _56173_ (_11397_, _11394_, _35722_);
  or _56174_ (_11398_, _11397_, _11396_);
  or _56175_ (_11399_, _11093_, _33942_);
  and _56176_ (_11400_, _11399_, _38997_);
  and _56177_ (_39058_[6], _11400_, _11398_);
  and _56178_ (_39019_, t0_i, _38997_);
  and _56179_ (_39020_, t1_i, _38997_);
  and _56180_ (_11401_, _11090_, _11356_);
  and _56181_ (_11402_, _11401_, _33633_);
  nand _56182_ (_11403_, _11402_, _34221_);
  not _56183_ (_11404_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _56184_ (_11405_, _11404_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  not _56185_ (_11406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _56186_ (_11407_, _11406_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _56187_ (_11408_, t1_i);
  and _56188_ (_11409_, _11408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _56189_ (_11410_, _11409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or _56190_ (_11411_, _11410_, _11407_);
  and _56191_ (_11412_, _11411_, _11405_);
  and _56192_ (_11413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _56193_ (_11414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _56194_ (_11415_, _11414_, _11413_);
  and _56195_ (_11416_, _11415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _56196_ (_11417_, _11416_, _11412_);
  and _56197_ (_11418_, _11417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _56198_ (_11419_, _11418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  not _56199_ (_11420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _56200_ (_11421_, _11420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _56201_ (_11422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _56202_ (_11423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _11422_);
  nor _56203_ (_11424_, _11423_, _11421_);
  and _56204_ (_11425_, _11090_, _11383_);
  and _56205_ (_11426_, _11425_, _33633_);
  nor _56206_ (_11427_, _11426_, _11424_);
  and _56207_ (_11428_, _11427_, _11419_);
  or _56208_ (_11429_, _11428_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _56209_ (_11430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _56210_ (_11431_, _11430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _56211_ (_11432_, _11431_, _11417_);
  nand _56212_ (_11433_, _11432_, _11427_);
  and _56213_ (_11434_, _11433_, _11429_);
  and _56214_ (_11435_, _11419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _56215_ (_11436_, _11435_, _11421_);
  nand _56216_ (_11437_, _11436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _56217_ (_11438_, _11437_, _11426_);
  or _56218_ (_11439_, _11438_, _11434_);
  or _56219_ (_11440_, _11439_, _11402_);
  and _56220_ (_11441_, _11440_, _38997_);
  and _56221_ (_39021_[7], _11441_, _11403_);
  not _56222_ (_11442_, _11402_);
  and _56223_ (_11443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _56224_ (_11444_, _11443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _56225_ (_11445_, _11444_, _11417_);
  and _56226_ (_11446_, _11445_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _56227_ (_11447_, _11446_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _56228_ (_11448_, _11447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _56229_ (_11449_, _11448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _56230_ (_11450_, _11449_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _56231_ (_11451_, _11450_, _11431_);
  not _56232_ (_11452_, _11423_);
  nor _56233_ (_11453_, _11431_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _56234_ (_11454_, _11453_, _11452_);
  nor _56235_ (_11455_, _11454_, _11451_);
  and _56236_ (_11456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _56237_ (_11457_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _56238_ (_11458_, _11450_);
  and _56239_ (_11459_, _11458_, _11457_);
  or _56240_ (_11460_, _11459_, _11456_);
  or _56241_ (_11461_, _11460_, _11455_);
  nor _56242_ (_11462_, _11449_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _56243_ (_11463_, _11462_, _11426_);
  and _56244_ (_11464_, _11463_, _11461_);
  not _56245_ (_11465_, _11426_);
  nor _56246_ (_11466_, _11465_, _34221_);
  or _56247_ (_11467_, _11466_, _11464_);
  and _56248_ (_11468_, _11467_, _11442_);
  and _56249_ (_11469_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _56250_ (_11470_, _11469_, _11468_);
  and _56251_ (_39022_[7], _11470_, _38997_);
  not _56252_ (_11471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _56253_ (_11472_, _11412_, _11471_);
  or _56254_ (_11473_, _11472_, _11451_);
  and _56255_ (_11474_, _11473_, _11423_);
  or _56256_ (_11475_, _11472_, _11450_);
  and _56257_ (_11476_, _11475_, _11457_);
  and _56258_ (_11477_, _11432_, _11421_);
  nand _56259_ (_11478_, _11412_, _11420_);
  and _56260_ (_11479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and _56261_ (_11480_, _11479_, _11478_);
  or _56262_ (_11481_, _11480_, _11477_);
  or _56263_ (_11482_, _11481_, _11476_);
  or _56264_ (_11483_, _11482_, _11474_);
  nor _56265_ (_11484_, _11402_, rst);
  and _56266_ (_11485_, _11484_, _11465_);
  and _56267_ (_39023_, _11485_, _11483_);
  and _56268_ (_11486_, _11090_, _11370_);
  and _56269_ (_11487_, _11486_, _33633_);
  nor _56270_ (_11488_, _11487_, rst);
  not _56271_ (_11489_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not _56272_ (_11490_, t0_i);
  and _56273_ (_11491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _11490_);
  nor _56274_ (_11492_, _11491_, _11489_);
  not _56275_ (_11493_, _11492_);
  not _56276_ (_11494_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _56277_ (_11495_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor _56278_ (_11496_, _11495_, _11494_);
  and _56279_ (_11497_, _11496_, _11493_);
  not _56280_ (_11498_, _11497_);
  and _56281_ (_11499_, _11498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _56282_ (_11500_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _56283_ (_11501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _56284_ (_11502_, _11501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _56285_ (_11503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _56286_ (_11504_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _56287_ (_11505_, _11504_, _11503_);
  and _56288_ (_11506_, _11505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _56289_ (_11507_, _11506_, _11497_);
  and _56290_ (_11508_, _11507_, _11502_);
  and _56291_ (_11509_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _56292_ (_11510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _56293_ (_11511_, _11510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _56294_ (_11512_, _11511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _56295_ (_11513_, _11512_, _11509_);
  and _56296_ (_11514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _56297_ (_11515_, _11514_, _11513_);
  or _56298_ (_11516_, _11515_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _56299_ (_11517_, _11516_, _11508_);
  nor _56300_ (_11518_, _11517_, _11500_);
  and _56301_ (_11519_, _11513_, _11507_);
  nand _56302_ (_11520_, _11519_, _11514_);
  and _56303_ (_11521_, _11520_, _11500_);
  nor _56304_ (_11522_, _11521_, _11518_);
  nor _56305_ (_11523_, _11522_, _11499_);
  and _56306_ (_11524_, _11090_, _11343_);
  and _56307_ (_11525_, _11524_, _33633_);
  nor _56308_ (_11526_, _11525_, _11523_);
  and _56309_ (_39024_, _11526_, _11488_);
  and _56310_ (_11527_, _11500_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _56311_ (_11528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _56312_ (_11529_, _11528_, _11507_);
  or _56313_ (_11530_, _11529_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _56314_ (_11531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _56315_ (_11532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _11531_);
  and _56316_ (_11533_, _11532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor _56317_ (_11534_, _11508_, _11500_);
  or _56318_ (_11535_, _11534_, _11533_);
  or _56319_ (_11536_, _11535_, _11487_);
  and _56320_ (_11537_, _11536_, _11530_);
  or _56321_ (_11538_, _11537_, _11527_);
  not _56322_ (_11539_, _11525_);
  not _56323_ (_11540_, _11487_);
  or _56324_ (_11541_, _11540_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _56325_ (_11542_, _11541_, _11539_);
  and _56326_ (_11543_, _11542_, _11538_);
  nor _56327_ (_11544_, _11539_, _34221_);
  or _56328_ (_11545_, _11544_, _11543_);
  and _56329_ (_39025_[7], _11545_, _38997_);
  nand _56330_ (_11546_, _11487_, _34221_);
  and _56331_ (_11547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _11531_);
  or _56332_ (_11548_, _11532_, _11547_);
  not _56333_ (_11549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _56334_ (_11550_, _11506_, _11502_);
  and _56335_ (_11551_, _11497_, _11531_);
  and _56336_ (_11552_, _11551_, _11550_);
  and _56337_ (_11553_, _11552_, _11513_);
  and _56338_ (_11554_, _11553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _56339_ (_11555_, _11554_, _11549_);
  and _56340_ (_11556_, _11554_, _11549_);
  or _56341_ (_11557_, _11556_, _11555_);
  and _56342_ (_11558_, _11557_, _11548_);
  and _56343_ (_11559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _56344_ (_11560_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _56345_ (_11561_, _11560_, _11512_);
  and _56346_ (_11562_, _11561_, _11509_);
  and _56347_ (_11563_, _11562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _56348_ (_11564_, _11563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _56349_ (_11565_, _11560_, _11515_);
  and _56350_ (_11566_, _11565_, _11564_);
  and _56351_ (_11567_, _11566_, _11559_);
  and _56352_ (_11568_, _11519_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _56353_ (_11569_, _11568_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _56354_ (_11570_, _11569_, _11521_);
  or _56355_ (_11571_, _11570_, _11567_);
  or _56356_ (_11572_, _11571_, _11558_);
  or _56357_ (_11573_, _11572_, _11487_);
  and _56358_ (_11574_, _11573_, _11539_);
  and _56359_ (_11575_, _11574_, _11546_);
  and _56360_ (_11576_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _56361_ (_11577_, _11576_, _11575_);
  and _56362_ (_39026_[7], _11577_, _38997_);
  or _56363_ (_11578_, _11560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and _56364_ (_11579_, _11559_, _38997_);
  and _56365_ (_11580_, _11579_, _11578_);
  not _56366_ (_11581_, _11560_);
  or _56367_ (_11582_, _11581_, _11515_);
  nand _56368_ (_11583_, _11582_, _11580_);
  nor _56369_ (_11584_, _11583_, _11487_);
  and _56370_ (_39027_, _11584_, _11539_);
  and _56371_ (_11585_, _34254_, _33633_);
  and _56372_ (_11586_, _11585_, _33662_);
  or _56373_ (_11587_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _56374_ (_11588_, _11587_, _38997_);
  nand _56375_ (_11589_, _11586_, _34221_);
  and _56376_ (_39028_[7], _11589_, _11588_);
  and _56377_ (_11590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _56378_ (_11591_, _11590_, _11426_);
  not _56379_ (_11592_, _11591_);
  and _56380_ (_11593_, _11592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _56381_ (_11594_, _11431_, _11416_);
  and _56382_ (_11595_, _11594_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _56383_ (_11596_, _11595_, _11421_);
  not _56384_ (_11597_, _11590_);
  and _56385_ (_11598_, _11412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _56386_ (_11599_, _11412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _56387_ (_11600_, _11599_, _11598_);
  and _56388_ (_11601_, _11600_, _11597_);
  nor _56389_ (_11602_, _11601_, _11596_);
  nor _56390_ (_11603_, _11602_, _11426_);
  or _56391_ (_11604_, _11603_, _11402_);
  or _56392_ (_11605_, _11604_, _11593_);
  nand _56393_ (_11606_, _11402_, _34148_);
  and _56394_ (_11607_, _11606_, _38997_);
  and _56395_ (_39021_[0], _11607_, _11605_);
  or _56396_ (_11608_, _11442_, _34122_);
  and _56397_ (_11609_, _11598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _56398_ (_11610_, _11598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _56399_ (_11611_, _11610_, _11609_);
  and _56400_ (_11612_, _11611_, _11591_);
  and _56401_ (_11613_, _11592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand _56402_ (_11614_, _11477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _56403_ (_11615_, _11614_, _11426_);
  or _56404_ (_11616_, _11615_, _11613_);
  or _56405_ (_11617_, _11616_, _11612_);
  or _56406_ (_11618_, _11617_, _11402_);
  and _56407_ (_11619_, _11618_, _38997_);
  and _56408_ (_39021_[1], _11619_, _11608_);
  or _56409_ (_11620_, _11442_, _34089_);
  and _56410_ (_11621_, _11598_, _11413_);
  nor _56411_ (_11622_, _11609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _56412_ (_11623_, _11622_, _11621_);
  and _56413_ (_11624_, _11623_, _11591_);
  and _56414_ (_11625_, _11592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nand _56415_ (_11626_, _11436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _56416_ (_11627_, _11626_, _11426_);
  or _56417_ (_11628_, _11627_, _11625_);
  or _56418_ (_11629_, _11628_, _11624_);
  or _56419_ (_11630_, _11629_, _11402_);
  and _56420_ (_11631_, _11630_, _38997_);
  and _56421_ (_39021_[2], _11631_, _11620_);
  nand _56422_ (_11632_, _11402_, _34052_);
  and _56423_ (_11633_, _11415_, _11412_);
  nor _56424_ (_11634_, _11621_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _56425_ (_11635_, _11634_, _11633_);
  and _56426_ (_11636_, _11635_, _11591_);
  and _56427_ (_11637_, _11592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand _56428_ (_11638_, _11477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _56429_ (_11639_, _11638_, _11426_);
  or _56430_ (_11640_, _11639_, _11637_);
  or _56431_ (_11641_, _11640_, _11636_);
  or _56432_ (_11642_, _11641_, _11402_);
  and _56433_ (_11643_, _11642_, _38997_);
  and _56434_ (_39021_[3], _11643_, _11632_);
  nand _56435_ (_11644_, _11402_, _34017_);
  and _56436_ (_11645_, _11592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _56437_ (_11646_, _11436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _56438_ (_11647_, _11633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _56439_ (_11648_, _11647_, _11417_);
  and _56440_ (_11649_, _11648_, _11597_);
  nor _56441_ (_11650_, _11649_, _11646_);
  nor _56442_ (_11651_, _11650_, _11426_);
  or _56443_ (_11652_, _11651_, _11645_);
  or _56444_ (_11653_, _11652_, _11402_);
  and _56445_ (_11654_, _11653_, _38997_);
  and _56446_ (_39021_[4], _11654_, _11644_);
  or _56447_ (_11655_, _11442_, _33978_);
  not _56448_ (_11656_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _56449_ (_11657_, _11427_, _11656_);
  and _56450_ (_11658_, _11436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not _56451_ (_11659_, _11424_);
  nor _56452_ (_11660_, _11417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _56453_ (_11661_, _11660_, _11418_);
  and _56454_ (_11662_, _11661_, _11659_);
  nor _56455_ (_11663_, _11662_, _11658_);
  nor _56456_ (_11664_, _11663_, _11426_);
  or _56457_ (_11665_, _11664_, _11657_);
  or _56458_ (_11666_, _11665_, _11402_);
  and _56459_ (_11667_, _11666_, _38997_);
  and _56460_ (_39021_[5], _11667_, _11655_);
  or _56461_ (_11668_, _11442_, _33942_);
  not _56462_ (_11669_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _56463_ (_11670_, _11427_, _11669_);
  and _56464_ (_11671_, _11421_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _56465_ (_11672_, _11671_, _11412_);
  and _56466_ (_11673_, _11672_, _11594_);
  or _56467_ (_11674_, _11418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand _56468_ (_11675_, _11674_, _11659_);
  nor _56469_ (_11676_, _11675_, _11419_);
  nor _56470_ (_11677_, _11676_, _11673_);
  nor _56471_ (_11678_, _11677_, _11426_);
  or _56472_ (_11679_, _11678_, _11670_);
  or _56473_ (_11680_, _11679_, _11402_);
  and _56474_ (_11681_, _11680_, _38997_);
  and _56475_ (_39021_[6], _11681_, _11668_);
  not _56476_ (_11682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _56477_ (_11683_, _11417_, _11422_);
  nor _56478_ (_11684_, _11431_, _11420_);
  not _56479_ (_11685_, _11684_);
  and _56480_ (_11686_, _11685_, _11683_);
  and _56481_ (_11687_, _11686_, _11682_);
  nor _56482_ (_11688_, _11686_, _11682_);
  or _56483_ (_11689_, _11688_, _11687_);
  or _56484_ (_11690_, _11689_, _11426_);
  nand _56485_ (_11691_, _11426_, _34148_);
  and _56486_ (_11692_, _11691_, _11690_);
  or _56487_ (_11693_, _11692_, _11402_);
  nand _56488_ (_11694_, _11402_, _11682_);
  and _56489_ (_11695_, _11694_, _38997_);
  and _56490_ (_39022_[0], _11695_, _11693_);
  or _56491_ (_11696_, _11465_, _34122_);
  not _56492_ (_11697_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _56493_ (_11698_, _11432_, _11452_);
  not _56494_ (_11699_, _11698_);
  nor _56495_ (_11700_, _11683_, _11423_);
  nor _56496_ (_11701_, _11700_, _11682_);
  and _56497_ (_11702_, _11701_, _11699_);
  nor _56498_ (_11703_, _11702_, _11697_);
  and _56499_ (_11704_, _11702_, _11697_);
  or _56500_ (_11705_, _11704_, _11703_);
  or _56501_ (_11706_, _11705_, _11426_);
  and _56502_ (_11707_, _11706_, _11442_);
  and _56503_ (_11708_, _11707_, _11696_);
  and _56504_ (_11709_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _56505_ (_11710_, _11709_, _11708_);
  and _56506_ (_39022_[1], _11710_, _38997_);
  or _56507_ (_11711_, _11465_, _34089_);
  and _56508_ (_11712_, _11445_, _11422_);
  and _56509_ (_11713_, _11685_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _56510_ (_11714_, _11713_, _11712_);
  or _56511_ (_11715_, _11684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _56512_ (_11716_, _11715_);
  and _56513_ (_11717_, _11443_, _11417_);
  and _56514_ (_11718_, _11717_, _11716_);
  or _56515_ (_11719_, _11718_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _56516_ (_11720_, _11719_, _11714_);
  or _56517_ (_11721_, _11720_, _11426_);
  and _56518_ (_11722_, _11721_, _11442_);
  and _56519_ (_11723_, _11722_, _11711_);
  and _56520_ (_11724_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _56521_ (_11725_, _11724_, _11723_);
  and _56522_ (_39022_[2], _11725_, _38997_);
  nand _56523_ (_11726_, _11426_, _34052_);
  or _56524_ (_11727_, _11712_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _56525_ (_11728_, _11712_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _56526_ (_11729_, _11728_, _11727_);
  or _56527_ (_11730_, _11729_, _11423_);
  and _56528_ (_11731_, _11443_, _11594_);
  and _56529_ (_11732_, _11731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _56530_ (_11733_, _11732_, _11412_);
  nor _56531_ (_11734_, _11733_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _56532_ (_11735_, _11733_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _56533_ (_11736_, _11735_, _11734_);
  or _56534_ (_11737_, _11736_, _11452_);
  and _56535_ (_11738_, _11737_, _11730_);
  or _56536_ (_11739_, _11738_, _11426_);
  and _56537_ (_11740_, _11739_, _11442_);
  and _56538_ (_11741_, _11740_, _11726_);
  and _56539_ (_11742_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _56540_ (_11743_, _11742_, _11741_);
  and _56541_ (_39022_[3], _11743_, _38997_);
  nand _56542_ (_11744_, _11426_, _34017_);
  or _56543_ (_11745_, _11735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _56544_ (_11746_, _11447_, _11431_);
  and _56545_ (_11747_, _11746_, _11423_);
  and _56546_ (_11748_, _11747_, _11745_);
  and _56547_ (_11749_, _11443_, _11416_);
  and _56548_ (_11750_, _11749_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _56549_ (_11751_, _11750_, _11412_);
  and _56550_ (_11752_, _11751_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _56551_ (_11753_, _11752_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _56552_ (_11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  not _56553_ (_11755_, _11447_);
  and _56554_ (_11756_, _11755_, _11457_);
  or _56555_ (_11757_, _11756_, _11754_);
  and _56556_ (_11758_, _11757_, _11753_);
  or _56557_ (_11759_, _11758_, _11748_);
  or _56558_ (_11760_, _11759_, _11426_);
  and _56559_ (_11761_, _11760_, _11442_);
  and _56560_ (_11762_, _11761_, _11744_);
  and _56561_ (_11763_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _56562_ (_11764_, _11763_, _11762_);
  and _56563_ (_39022_[4], _11764_, _38997_);
  or _56564_ (_11765_, _11465_, _33978_);
  not _56565_ (_11766_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _56566_ (_11767_, _11716_, _11447_);
  nor _56567_ (_11768_, _11767_, _11766_);
  and _56568_ (_11769_, _11767_, _11766_);
  or _56569_ (_11770_, _11769_, _11768_);
  or _56570_ (_11771_, _11770_, _11426_);
  and _56571_ (_11772_, _11771_, _11442_);
  and _56572_ (_11773_, _11772_, _11765_);
  and _56573_ (_11774_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _56574_ (_11775_, _11774_, _11773_);
  and _56575_ (_39022_[5], _11775_, _38997_);
  or _56576_ (_11776_, _11465_, _33942_);
  not _56577_ (_11777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _56578_ (_11778_, _11716_, _11448_);
  nor _56579_ (_11779_, _11778_, _11777_);
  and _56580_ (_11780_, _11778_, _11777_);
  or _56581_ (_11781_, _11780_, _11779_);
  or _56582_ (_11782_, _11781_, _11426_);
  and _56583_ (_11783_, _11782_, _11442_);
  and _56584_ (_11784_, _11783_, _11776_);
  and _56585_ (_11785_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _56586_ (_11786_, _11785_, _11784_);
  and _56587_ (_39022_[6], _11786_, _38997_);
  nor _56588_ (_11787_, _11498_, _11487_);
  or _56589_ (_11788_, _11787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _56590_ (_11789_, _11532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _56591_ (_11790_, _11789_, _11550_);
  and _56592_ (_11791_, _11497_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand _56593_ (_11792_, _11791_, _11790_);
  or _56594_ (_11793_, _11792_, _11487_);
  and _56595_ (_11794_, _11793_, _11788_);
  or _56596_ (_11795_, _11794_, _11525_);
  nand _56597_ (_11796_, _11525_, _34148_);
  and _56598_ (_11797_, _11796_, _38997_);
  and _56599_ (_39025_[0], _11797_, _11795_);
  or _56600_ (_11798_, _11539_, _34122_);
  and _56601_ (_11799_, _11487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _56602_ (_11800_, _11799_, _11525_);
  and _56603_ (_11801_, _11800_, _38997_);
  nor _56604_ (_11802_, _11791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _56605_ (_11803_, _11791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _56606_ (_11804_, _11803_, _11802_);
  and _56607_ (_11805_, _11532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _56608_ (_11806_, _11805_, _11508_);
  or _56609_ (_11807_, _11806_, _11804_);
  and _56610_ (_11808_, _11807_, _11488_);
  or _56611_ (_11809_, _11808_, _11801_);
  and _56612_ (_39025_[1], _11809_, _11798_);
  or _56613_ (_11810_, _11539_, _34089_);
  nor _56614_ (_11811_, _11803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _56615_ (_11812_, _11791_, _11503_);
  nor _56616_ (_11813_, _11812_, _11811_);
  and _56617_ (_11814_, _11532_, _11508_);
  and _56618_ (_11815_, _11814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _56619_ (_11816_, _11815_, _11813_);
  nor _56620_ (_11817_, _11816_, _11487_);
  and _56621_ (_11818_, _11487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _56622_ (_11819_, _11818_, _11817_);
  or _56623_ (_11820_, _11819_, _11525_);
  and _56624_ (_11821_, _11820_, _38997_);
  and _56625_ (_39025_[2], _11821_, _11810_);
  and _56626_ (_11822_, _11505_, _11497_);
  nor _56627_ (_11823_, _11812_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _56628_ (_11824_, _11823_, _11822_);
  and _56629_ (_11825_, _11814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _56630_ (_11826_, _11825_, _11824_);
  nor _56631_ (_11827_, _11826_, _11487_);
  and _56632_ (_11828_, _11487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _56633_ (_11829_, _11828_, _11827_);
  and _56634_ (_11830_, _11829_, _11539_);
  nor _56635_ (_11831_, _11539_, _34052_);
  or _56636_ (_11832_, _11831_, _11830_);
  and _56637_ (_39025_[3], _11832_, _38997_);
  nor _56638_ (_11833_, _11822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _56639_ (_11834_, _11833_, _11507_);
  and _56640_ (_11835_, _11814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _56641_ (_11836_, _11835_, _11834_);
  nor _56642_ (_11837_, _11836_, _11487_);
  and _56643_ (_11838_, _11487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _56644_ (_11839_, _11838_, _11837_);
  and _56645_ (_11840_, _11839_, _11539_);
  nor _56646_ (_11841_, _11539_, _34017_);
  or _56647_ (_11842_, _11841_, _11840_);
  and _56648_ (_39025_[4], _11842_, _38997_);
  or _56649_ (_11843_, _11539_, _33978_);
  nand _56650_ (_11844_, _11814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not _56651_ (_11845_, _11500_);
  nand _56652_ (_11846_, _11507_, _11845_);
  or _56653_ (_11847_, _11846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _56654_ (_11848_, _11847_, _11844_);
  nor _56655_ (_11849_, _11848_, _11487_);
  not _56656_ (_11850_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _56657_ (_11851_, _11846_, _11850_);
  or _56658_ (_11852_, _11851_, _11487_);
  and _56659_ (_11853_, _11852_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _56660_ (_11854_, _11853_, _11849_);
  or _56661_ (_11855_, _11854_, _11525_);
  and _56662_ (_11856_, _11855_, _38997_);
  and _56663_ (_39025_[5], _11856_, _11843_);
  and _56664_ (_11857_, _11852_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _56665_ (_11858_, _11532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _56666_ (_11859_, _11858_, _11497_);
  and _56667_ (_11860_, _11859_, _11550_);
  nor _56668_ (_11861_, _11851_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor _56669_ (_11862_, _11861_, _11860_);
  nor _56670_ (_11863_, _11862_, _11487_);
  or _56671_ (_11864_, _11863_, _11857_);
  and _56672_ (_11865_, _11864_, _11539_);
  and _56673_ (_11866_, _11525_, _33942_);
  or _56674_ (_11867_, _11866_, _11865_);
  and _56675_ (_39025_[6], _11867_, _38997_);
  or _56676_ (_11868_, _11552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _56677_ (_11869_, _11552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not _56678_ (_11870_, _11869_);
  and _56679_ (_11871_, _11870_, _11548_);
  and _56680_ (_11872_, _11871_, _11868_);
  and _56681_ (_11873_, _11560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _56682_ (_11874_, _11560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _56683_ (_11875_, _11874_, _11559_);
  nor _56684_ (_11876_, _11875_, _11873_);
  and _56685_ (_11877_, _11507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _56686_ (_11878_, _11507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _56687_ (_11879_, _11878_, _11500_);
  nor _56688_ (_11880_, _11879_, _11877_);
  or _56689_ (_11881_, _11880_, _11876_);
  nor _56690_ (_11882_, _11881_, _11872_);
  nand _56691_ (_11883_, _11882_, _11540_);
  nand _56692_ (_11884_, _11487_, _34148_);
  and _56693_ (_11885_, _11884_, _11539_);
  and _56694_ (_11886_, _11885_, _11883_);
  and _56695_ (_11887_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _56696_ (_11888_, _11887_, _11886_);
  and _56697_ (_39026_[0], _11888_, _38997_);
  or _56698_ (_11889_, _11540_, _34122_);
  or _56699_ (_11890_, _11869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _56700_ (_11891_, _11550_, _11497_);
  and _56701_ (_11892_, _11891_, _11510_);
  not _56702_ (_11893_, _11892_);
  or _56703_ (_11894_, _11893_, _11532_);
  and _56704_ (_11895_, _11894_, _11548_);
  and _56705_ (_11896_, _11895_, _11890_);
  and _56706_ (_11897_, _11560_, _11510_);
  or _56707_ (_11898_, _11873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _56708_ (_11899_, _11898_, _11559_);
  nor _56709_ (_11900_, _11899_, _11897_);
  and _56710_ (_11901_, _11877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _56711_ (_11902_, _11877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _56712_ (_11903_, _11902_, _11500_);
  nor _56713_ (_11904_, _11903_, _11901_);
  or _56714_ (_11905_, _11904_, _11900_);
  or _56715_ (_11906_, _11905_, _11896_);
  or _56716_ (_11907_, _11906_, _11487_);
  and _56717_ (_11908_, _11907_, _11539_);
  and _56718_ (_11909_, _11908_, _11889_);
  and _56719_ (_11910_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _56720_ (_11911_, _11910_, _11909_);
  and _56721_ (_39026_[1], _11911_, _38997_);
  or _56722_ (_11912_, _11540_, _34089_);
  or _56723_ (_11913_, _11892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _56724_ (_11914_, _11891_, _11511_);
  not _56725_ (_11915_, _11914_);
  and _56726_ (_11916_, _11915_, _11547_);
  and _56727_ (_11917_, _11916_, _11913_);
  and _56728_ (_11918_, _11510_, _11497_);
  and _56729_ (_11919_, _11918_, _11506_);
  or _56730_ (_11920_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _56731_ (_11921_, _11511_, _11507_);
  nor _56732_ (_11922_, _11921_, _11845_);
  and _56733_ (_11923_, _11922_, _11920_);
  and _56734_ (_11924_, _11897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _56735_ (_11925_, _11924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _56736_ (_11926_, _11560_, _11511_);
  nand _56737_ (_11927_, _11926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _56738_ (_11928_, _11927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _56739_ (_11929_, _11928_, _11925_);
  or _56740_ (_11930_, _11929_, _11923_);
  or _56741_ (_11931_, _11930_, _11917_);
  or _56742_ (_11932_, _11931_, _11487_);
  and _56743_ (_11933_, _11932_, _11539_);
  and _56744_ (_11934_, _11933_, _11912_);
  and _56745_ (_11935_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _56746_ (_11936_, _11935_, _11934_);
  and _56747_ (_39026_[2], _11936_, _38997_);
  nand _56748_ (_11937_, _11487_, _34052_);
  not _56749_ (_11938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _56750_ (_11939_, _11914_, _11531_);
  nor _56751_ (_11940_, _11939_, _11938_);
  and _56752_ (_11941_, _11939_, _11938_);
  or _56753_ (_11942_, _11941_, _11940_);
  and _56754_ (_11943_, _11942_, _11548_);
  or _56755_ (_11944_, _11926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _56756_ (_11945_, _11561_);
  and _56757_ (_11946_, _11945_, _11559_);
  and _56758_ (_11947_, _11946_, _11944_);
  or _56759_ (_11948_, _11921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _56760_ (_11949_, _11512_, _11507_);
  nor _56761_ (_11950_, _11949_, _11845_);
  and _56762_ (_11951_, _11950_, _11948_);
  or _56763_ (_11952_, _11951_, _11947_);
  or _56764_ (_11953_, _11952_, _11943_);
  or _56765_ (_11954_, _11953_, _11487_);
  and _56766_ (_11955_, _11954_, _11539_);
  and _56767_ (_11956_, _11955_, _11937_);
  and _56768_ (_11957_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _56769_ (_11958_, _11957_, _11956_);
  and _56770_ (_39026_[3], _11958_, _38997_);
  nand _56771_ (_11959_, _11487_, _34017_);
  or _56772_ (_11960_, _11949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _56773_ (_11961_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _56774_ (_11962_, _11961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _56775_ (_11963_, _11962_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _56776_ (_11964_, _11963_, _11845_);
  and _56777_ (_11965_, _11964_, _11960_);
  and _56778_ (_11966_, _11512_, _11497_);
  and _56779_ (_11967_, _11966_, _11550_);
  or _56780_ (_11968_, _11967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _56781_ (_11969_, _11967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not _56782_ (_11970_, _11969_);
  and _56783_ (_11971_, _11970_, _11547_);
  and _56784_ (_11972_, _11971_, _11968_);
  and _56785_ (_11973_, _11561_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _56786_ (_11974_, _11973_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _56787_ (_11975_, _11561_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _56788_ (_11976_, _11975_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _56789_ (_11977_, _11976_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _56790_ (_11978_, _11977_, _11974_);
  or _56791_ (_11979_, _11978_, _11972_);
  or _56792_ (_11980_, _11979_, _11965_);
  or _56793_ (_11981_, _11980_, _11487_);
  and _56794_ (_11982_, _11981_, _11539_);
  and _56795_ (_11983_, _11982_, _11959_);
  and _56796_ (_11984_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _56797_ (_11985_, _11984_, _11983_);
  and _56798_ (_39026_[4], _11985_, _38997_);
  or _56799_ (_11986_, _11540_, _33978_);
  not _56800_ (_11987_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _56801_ (_11988_, _11963_, _11987_);
  nor _56802_ (_11989_, _11963_, _11987_);
  or _56803_ (_11990_, _11989_, _11988_);
  and _56804_ (_11991_, _11990_, _11500_);
  not _56805_ (_11992_, _11562_);
  and _56806_ (_11993_, _11992_, _11559_);
  or _56807_ (_11994_, _11973_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _56808_ (_11995_, _11994_, _11993_);
  and _56809_ (_11996_, _11969_, _11531_);
  nand _56810_ (_11997_, _11996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _56811_ (_11998_, _11996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _56812_ (_11999_, _11998_, _11997_);
  and _56813_ (_12000_, _11999_, _11548_);
  or _56814_ (_12001_, _12000_, _11995_);
  or _56815_ (_12002_, _12001_, _11991_);
  or _56816_ (_12003_, _12002_, _11487_);
  and _56817_ (_12004_, _12003_, _11539_);
  and _56818_ (_12005_, _12004_, _11986_);
  and _56819_ (_12006_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _56820_ (_12007_, _12006_, _12005_);
  and _56821_ (_39026_[5], _12007_, _38997_);
  or _56822_ (_12008_, _11540_, _33942_);
  or _56823_ (_12009_, _11553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _56824_ (_12010_, _12009_, _11548_);
  nor _56825_ (_12011_, _12010_, _11554_);
  or _56826_ (_12012_, _11562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _56827_ (_12013_, _11563_);
  and _56828_ (_12014_, _12013_, _11559_);
  and _56829_ (_12015_, _12014_, _12012_);
  or _56830_ (_12016_, _11519_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _56831_ (_12017_, _11568_, _11845_);
  and _56832_ (_12018_, _12017_, _12016_);
  or _56833_ (_12019_, _12018_, _12015_);
  or _56834_ (_12020_, _12019_, _12011_);
  or _56835_ (_12021_, _12020_, _11487_);
  and _56836_ (_12022_, _12021_, _11539_);
  and _56837_ (_12023_, _12022_, _12008_);
  and _56838_ (_12024_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _56839_ (_12025_, _12024_, _12023_);
  and _56840_ (_39026_[6], _12025_, _38997_);
  nand _56841_ (_12026_, _11586_, _34148_);
  or _56842_ (_12027_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _56843_ (_12028_, _12027_, _38997_);
  and _56844_ (_39028_[0], _12028_, _12026_);
  or _56845_ (_12029_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _56846_ (_12030_, _12029_, _38997_);
  not _56847_ (_12031_, _11586_);
  or _56848_ (_12032_, _12031_, _34122_);
  and _56849_ (_39028_[1], _12032_, _12030_);
  or _56850_ (_12033_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _56851_ (_12034_, _12033_, _38997_);
  or _56852_ (_12035_, _12031_, _34089_);
  and _56853_ (_39028_[2], _12035_, _12034_);
  or _56854_ (_12036_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _56855_ (_12037_, _12036_, _38997_);
  nand _56856_ (_12038_, _11586_, _34052_);
  and _56857_ (_39028_[3], _12038_, _12037_);
  or _56858_ (_12039_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _56859_ (_12040_, _12039_, _38997_);
  nand _56860_ (_12041_, _11586_, _34017_);
  and _56861_ (_39028_[4], _12041_, _12040_);
  or _56862_ (_12042_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _56863_ (_12043_, _12042_, _38997_);
  or _56864_ (_12044_, _12031_, _33978_);
  and _56865_ (_39028_[5], _12044_, _12043_);
  or _56866_ (_12045_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _56867_ (_12046_, _12045_, _38997_);
  or _56868_ (_12047_, _12031_, _33942_);
  and _56869_ (_39028_[6], _12047_, _12046_);
  and _56870_ (_12048_, _33630_, _34232_);
  and _56871_ (_12049_, _12048_, _11085_);
  and _56872_ (_12050_, _12049_, _11075_);
  or _56873_ (_12051_, _12050_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nor _56874_ (_12052_, _33604_, _33591_);
  and _56875_ (_12053_, _12052_, _33632_);
  and _56876_ (_12054_, _12053_, _11076_);
  not _56877_ (_12055_, _12054_);
  and _56878_ (_12056_, _12055_, _12051_);
  nand _56879_ (_12057_, _12050_, _35722_);
  and _56880_ (_12058_, _12057_, _12056_);
  nor _56881_ (_12059_, _12055_, _34221_);
  or _56882_ (_12060_, _12059_, _12058_);
  and _56883_ (_39011_[7], _12060_, _38997_);
  and _56884_ (_12061_, _34251_, _33604_);
  and _56885_ (_12062_, _12061_, _11084_);
  and _56886_ (_12063_, _12062_, _12048_);
  and _56887_ (_12064_, _12063_, _11075_);
  or _56888_ (_12065_, _12064_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _56889_ (_12066_, _33604_, _34232_);
  and _56890_ (_12067_, _12066_, _33632_);
  and _56891_ (_12068_, _12067_, _11091_);
  not _56892_ (_12069_, _12068_);
  and _56893_ (_12070_, _12069_, _12065_);
  nand _56894_ (_12071_, _12064_, _35722_);
  and _56895_ (_12072_, _12071_, _12070_);
  nor _56896_ (_12073_, _12069_, _34221_);
  or _56897_ (_12074_, _12073_, _12072_);
  and _56898_ (_39010_[7], _12074_, _38997_);
  and _56899_ (_12075_, _12062_, _11081_);
  nand _56900_ (_12076_, _12075_, _33558_);
  and _56901_ (_12077_, _12076_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _56902_ (_12078_, _11091_, _33633_);
  or _56903_ (_12079_, _12078_, _12077_);
  nor _56904_ (_12080_, _11393_, _35722_);
  nand _56905_ (_12081_, _33558_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _56906_ (_12082_, _12081_, _11391_);
  or _56907_ (_12083_, _12082_, _12080_);
  and _56908_ (_12084_, _12083_, _12075_);
  or _56909_ (_12085_, _12084_, _12079_);
  not _56910_ (_12086_, _12078_);
  or _56911_ (_12087_, _12086_, _33942_);
  and _56912_ (_12088_, _12087_, _38997_);
  and _56913_ (_39009_[3], _12088_, _12085_);
  nor _56914_ (_12089_, _10898_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not _56915_ (_12090_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _56916_ (_12091_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _56917_ (_12092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _56918_ (_12093_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _12092_);
  and _56919_ (_12094_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _56920_ (_12095_, _12094_, _12093_);
  nor _56921_ (_12096_, _12095_, _12091_);
  or _56922_ (_12097_, _12096_, _12090_);
  and _56923_ (_12098_, _12092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _56924_ (_12099_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _56925_ (_12100_, _12099_, _12098_);
  nor _56926_ (_12101_, _12100_, _12091_);
  and _56927_ (_12102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _12092_);
  and _56928_ (_12103_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _56929_ (_12104_, _12103_, _12102_);
  nand _56930_ (_12105_, _12104_, _12101_);
  or _56931_ (_12106_, _12105_, _12097_);
  and _56932_ (_12107_, _12106_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _56933_ (_12108_, _12107_, _12089_);
  and _56934_ (_12109_, _11366_, _33633_);
  and _56935_ (_12110_, _12109_, _11075_);
  or _56936_ (_12111_, _12110_, _12108_);
  and _56937_ (_12112_, _12111_, _12086_);
  nand _56938_ (_12113_, _12110_, _35722_);
  and _56939_ (_12114_, _12113_, _12112_);
  nor _56940_ (_12115_, _12086_, _34221_);
  or _56941_ (_12116_, _12115_, _12114_);
  and _56942_ (_39008_, _12116_, _38997_);
  not _56943_ (_12117_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and _56944_ (_12118_, _12117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _56945_ (_12119_, _12104_, _12091_);
  not _56946_ (_12120_, _12119_);
  or _56947_ (_12121_, _12120_, _12101_);
  or _56948_ (_12122_, _12121_, _12097_);
  and _56949_ (_12123_, _12122_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _56950_ (_12124_, _12123_, _12118_);
  and _56951_ (_12125_, _12109_, _11383_);
  or _56952_ (_12126_, _12125_, _12124_);
  and _56953_ (_12127_, _12126_, _12086_);
  nand _56954_ (_12128_, _12125_, _35722_);
  and _56955_ (_12129_, _12128_, _12127_);
  and _56956_ (_12130_, _12078_, _33978_);
  or _56957_ (_12131_, _12130_, _12129_);
  and _56958_ (_39007_, _12131_, _38997_);
  not _56959_ (_12132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _56960_ (_12133_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _12132_);
  nand _56961_ (_12134_, _12096_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _56962_ (_12135_, _12119_, _12101_);
  or _56963_ (_12136_, _12135_, _12134_);
  and _56964_ (_12137_, _12136_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _56965_ (_12138_, _12137_, _12133_);
  and _56966_ (_12139_, _11585_, _11083_);
  or _56967_ (_12140_, _12139_, _12138_);
  and _56968_ (_12141_, _12140_, _12086_);
  nand _56969_ (_12142_, _12139_, _35722_);
  and _56970_ (_12143_, _12142_, _12141_);
  and _56971_ (_12144_, _12078_, _34122_);
  or _56972_ (_12145_, _12144_, _12143_);
  and _56973_ (_39006_, _12145_, _38997_);
  nand _56974_ (_12146_, _12109_, _11356_);
  nor _56975_ (_12147_, _12146_, _35722_);
  and _56976_ (_12148_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _56977_ (_12149_, _12134_, _12121_);
  and _56978_ (_12150_, _12149_, _12148_);
  and _56979_ (_12151_, _12150_, _12146_);
  or _56980_ (_12152_, _12151_, _12078_);
  or _56981_ (_12153_, _12152_, _12147_);
  nand _56982_ (_12154_, _12078_, _34052_);
  and _56983_ (_12155_, _12154_, _38997_);
  and _56984_ (_39005_, _12155_, _12153_);
  nand _56985_ (_12156_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _56986_ (_12157_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _12092_);
  and _56987_ (_12158_, _12157_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _56988_ (_12159_, _12158_, _12156_);
  or _56989_ (_12160_, _12159_, _12091_);
  and _56990_ (_12161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _56991_ (_12162_, _12161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _56992_ (_12163_, _12162_);
  and _56993_ (_12164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _56994_ (_12165_, _12164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _56995_ (_12166_, _12165_);
  and _56996_ (_12167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _56997_ (_12168_, _12167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _56998_ (_12169_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _56999_ (_12170_, _12169_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _57000_ (_12171_, _12170_, _12168_);
  and _57001_ (_12172_, _12171_, _12166_);
  and _57002_ (_12173_, _12172_, _12163_);
  not _57003_ (_12174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _57004_ (_12175_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _57005_ (_12176_, _12175_, _12174_);
  nand _57006_ (_12177_, _12176_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not _57007_ (_12178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _57008_ (_12179_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _57009_ (_12180_, _12179_, _12178_);
  and _57010_ (_12181_, _12180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _57011_ (_12182_, _12181_);
  and _57012_ (_12183_, _12182_, _12177_);
  nand _57013_ (_12184_, _12183_, _12173_);
  and _57014_ (_12185_, _12184_, _12160_);
  and _57015_ (_12186_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _57016_ (_12187_, _12186_, _12092_);
  and _57017_ (_12188_, _12187_, _12185_);
  not _57018_ (_12189_, _12188_);
  not _57019_ (_12190_, _12187_);
  and _57020_ (_12191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _12091_);
  not _57021_ (_12192_, _12191_);
  not _57022_ (_12193_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _57023_ (_12194_, _12164_, _12193_);
  not _57024_ (_12195_, _12194_);
  not _57025_ (_12196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _57026_ (_12197_, _12167_, _12196_);
  not _57027_ (_12198_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _57028_ (_12199_, _12169_, _12198_);
  nor _57029_ (_12200_, _12199_, _12197_);
  and _57030_ (_12201_, _12200_, _12195_);
  nor _57031_ (_12202_, _12201_, _12192_);
  not _57032_ (_12203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _57033_ (_12204_, _12176_, _12203_);
  not _57034_ (_12205_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _57035_ (_12206_, _12180_, _12205_);
  nor _57036_ (_12207_, _12206_, _12204_);
  not _57037_ (_12208_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _57038_ (_12209_, _12161_, _12208_);
  not _57039_ (_12210_, _12209_);
  and _57040_ (_12211_, _12210_, _12207_);
  nor _57041_ (_12212_, _12211_, _12192_);
  nor _57042_ (_12213_, _12212_, _12202_);
  or _57043_ (_12214_, _12213_, _12190_);
  and _57044_ (_12215_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _38997_);
  and _57045_ (_12216_, _12215_, _12214_);
  and _57046_ (_39004_[1], _12216_, _12189_);
  nor _57047_ (_12217_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _57048_ (_12218_, _12217_);
  not _57049_ (_12219_, _12185_);
  and _57050_ (_12220_, _12213_, _12219_);
  nor _57051_ (_12221_, _12220_, _12218_);
  nand _57052_ (_12222_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _38997_);
  nor _57053_ (_39003_[1], _12222_, _12221_);
  and _57054_ (_12223_, _12183_, _12163_);
  nand _57055_ (_12224_, _12223_, _12185_);
  or _57056_ (_12225_, _12212_, _12185_);
  and _57057_ (_12226_, _12225_, _12187_);
  and _57058_ (_12227_, _12226_, _12224_);
  or _57059_ (_12228_, _12227_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or _57060_ (_12229_, _12189_, _12172_);
  nor _57061_ (_12230_, _12190_, _12185_);
  nand _57062_ (_12231_, _12230_, _12202_);
  and _57063_ (_12232_, _12231_, _38997_);
  and _57064_ (_12233_, _12232_, _12229_);
  and _57065_ (_39002_[2], _12233_, _12228_);
  and _57066_ (_12234_, _12224_, _12217_);
  or _57067_ (_12235_, _12234_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _57068_ (_12236_, _12217_, _12185_);
  not _57069_ (_12237_, _12236_);
  or _57070_ (_12238_, _12237_, _12172_);
  or _57071_ (_12239_, _12212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand _57072_ (_12240_, _12217_, _12202_);
  and _57073_ (_12241_, _12240_, _12239_);
  or _57074_ (_12242_, _12241_, _12185_);
  and _57075_ (_12243_, _12242_, _38997_);
  and _57076_ (_12244_, _12243_, _12238_);
  and _57077_ (_39001_[2], _12244_, _12235_);
  nand _57078_ (_12245_, _12220_, _12091_);
  nor _57079_ (_12246_, _12092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand _57080_ (_12247_, _12246_, _12186_);
  and _57081_ (_12248_, _12247_, _38997_);
  and _57082_ (_39000_, _12248_, _12245_);
  and _57083_ (_12249_, _12220_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _57084_ (_12250_, _12092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _57085_ (_12251_, _12250_, _12246_);
  nor _57086_ (_12252_, _12251_, _12219_);
  or _57087_ (_12253_, _12252_, _12186_);
  or _57088_ (_12254_, _12253_, _12249_);
  not _57089_ (_12255_, _12186_);
  or _57090_ (_12256_, _12251_, _12255_);
  and _57091_ (_12257_, _12256_, _38997_);
  and _57092_ (_38999_[1], _12257_, _12254_);
  and _57093_ (_12258_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _38997_);
  and _57094_ (_38998_[7], _12258_, _12186_);
  and _57095_ (_38995_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _38997_);
  nor _57096_ (_12259_, _12220_, _12186_);
  and _57097_ (_12260_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _57098_ (_12261_, _12260_, _12259_);
  and _57099_ (_38998_[0], _12261_, _38997_);
  and _57100_ (_12262_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _57101_ (_12263_, _12262_, _12259_);
  and _57102_ (_38998_[1], _12263_, _38997_);
  and _57103_ (_12264_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _38997_);
  and _57104_ (_38998_[2], _12264_, _12186_);
  not _57105_ (_12265_, _12199_);
  nor _57106_ (_12266_, _12206_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _57107_ (_12267_, _12266_, _12204_);
  or _57108_ (_12268_, _12267_, _12209_);
  and _57109_ (_12269_, _12268_, _12265_);
  or _57110_ (_12270_, _12269_, _12197_);
  nor _57111_ (_12271_, _12213_, _12185_);
  and _57112_ (_12272_, _12271_, _12195_);
  and _57113_ (_12273_, _12272_, _12270_);
  not _57114_ (_12274_, _12170_);
  or _57115_ (_12275_, _12181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _57116_ (_12276_, _12275_, _12177_);
  or _57117_ (_12277_, _12276_, _12162_);
  and _57118_ (_12278_, _12277_, _12274_);
  or _57119_ (_12279_, _12278_, _12168_);
  and _57120_ (_12280_, _12185_, _12166_);
  and _57121_ (_12281_, _12280_, _12279_);
  or _57122_ (_12282_, _12281_, _12186_);
  or _57123_ (_12283_, _12282_, _12273_);
  or _57124_ (_12284_, _12255_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _57125_ (_12285_, _12284_, _38997_);
  and _57126_ (_38998_[3], _12285_, _12283_);
  not _57127_ (_12286_, _12168_);
  or _57128_ (_12287_, _12170_, _12162_);
  and _57129_ (_12288_, _12183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _57130_ (_12289_, _12288_, _12287_);
  and _57131_ (_12290_, _12289_, _12286_);
  and _57132_ (_12291_, _12290_, _12280_);
  nor _57133_ (_12292_, _12197_, _12194_);
  or _57134_ (_12293_, _12209_, _12199_);
  and _57135_ (_12294_, _12207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _57136_ (_12295_, _12294_, _12293_);
  and _57137_ (_12296_, _12295_, _12292_);
  and _57138_ (_12297_, _12296_, _12271_);
  or _57139_ (_12298_, _12297_, _12186_);
  or _57140_ (_12299_, _12298_, _12291_);
  or _57141_ (_12300_, _12255_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _57142_ (_12301_, _12300_, _38997_);
  and _57143_ (_38998_[4], _12301_, _12299_);
  and _57144_ (_12302_, _12210_, _12191_);
  nand _57145_ (_12303_, _12302_, _12201_);
  or _57146_ (_12304_, _12303_, _12207_);
  nor _57147_ (_12305_, _12304_, _12185_);
  nand _57148_ (_12306_, _12173_, _12160_);
  nor _57149_ (_12307_, _12306_, _12183_);
  or _57150_ (_12308_, _12307_, _12186_);
  or _57151_ (_12309_, _12308_, _12305_);
  or _57152_ (_12310_, _12255_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _57153_ (_12311_, _12310_, _38997_);
  and _57154_ (_38998_[5], _12311_, _12309_);
  and _57155_ (_12312_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _38997_);
  and _57156_ (_38998_[6], _12312_, _12186_);
  and _57157_ (_12313_, _12186_, _12092_);
  or _57158_ (_12314_, _12313_, _12221_);
  or _57159_ (_12315_, _12314_, _12230_);
  and _57160_ (_38999_[0], _12315_, _38997_);
  not _57161_ (_12316_, _12259_);
  and _57162_ (_12317_, _12316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _57163_ (_12318_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _57164_ (_12319_, _12181_, _12092_);
  or _57165_ (_12320_, _12319_, _12318_);
  nor _57166_ (_12321_, _12177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _57167_ (_12322_, _12321_, _12162_);
  nand _57168_ (_12323_, _12322_, _12320_);
  or _57169_ (_12324_, _12163_, _12094_);
  and _57170_ (_12325_, _12324_, _12323_);
  or _57171_ (_12326_, _12325_, _12170_);
  or _57172_ (_12327_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _12092_);
  or _57173_ (_12328_, _12327_, _12274_);
  and _57174_ (_12329_, _12328_, _12286_);
  and _57175_ (_12330_, _12329_, _12326_);
  and _57176_ (_12331_, _12168_, _12094_);
  or _57177_ (_12332_, _12331_, _12165_);
  or _57178_ (_12333_, _12332_, _12330_);
  or _57179_ (_12334_, _12327_, _12166_);
  and _57180_ (_12335_, _12334_, _12185_);
  and _57181_ (_12336_, _12335_, _12333_);
  and _57182_ (_12337_, _12206_, _12092_);
  or _57183_ (_12338_, _12337_, _12318_);
  and _57184_ (_12339_, _12204_, _12092_);
  nor _57185_ (_12340_, _12339_, _12209_);
  nand _57186_ (_12341_, _12340_, _12338_);
  or _57187_ (_12342_, _12210_, _12094_);
  and _57188_ (_12343_, _12342_, _12341_);
  or _57189_ (_12344_, _12343_, _12199_);
  not _57190_ (_12345_, _12197_);
  or _57191_ (_12346_, _12327_, _12265_);
  and _57192_ (_12347_, _12346_, _12345_);
  and _57193_ (_12348_, _12347_, _12344_);
  and _57194_ (_12349_, _12197_, _12094_);
  or _57195_ (_12350_, _12349_, _12194_);
  or _57196_ (_12351_, _12350_, _12348_);
  and _57197_ (_12352_, _12327_, _12271_);
  or _57198_ (_12353_, _12352_, _12272_);
  and _57199_ (_12354_, _12353_, _12351_);
  or _57200_ (_12355_, _12354_, _12336_);
  and _57201_ (_12356_, _12355_, _12255_);
  or _57202_ (_12357_, _12356_, _12317_);
  and _57203_ (_39001_[0], _12357_, _38997_);
  and _57204_ (_12358_, _12316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or _57205_ (_12359_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _12092_);
  and _57206_ (_12360_, _12359_, _12166_);
  or _57207_ (_12361_, _12360_, _12172_);
  or _57208_ (_12362_, _12319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _57209_ (_12363_, _12362_, _12322_);
  nand _57210_ (_12364_, _12162_, _12103_);
  nand _57211_ (_12365_, _12364_, _12171_);
  or _57212_ (_12366_, _12365_, _12363_);
  and _57213_ (_12367_, _12366_, _12361_);
  and _57214_ (_12368_, _12165_, _12103_);
  or _57215_ (_12369_, _12368_, _12367_);
  and _57216_ (_12370_, _12369_, _12185_);
  and _57217_ (_12371_, _12194_, _12103_);
  and _57218_ (_12372_, _12359_, _12195_);
  or _57219_ (_12373_, _12372_, _12201_);
  and _57220_ (_12374_, _12209_, _12103_);
  not _57221_ (_12375_, _12200_);
  or _57222_ (_12376_, _12337_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _57223_ (_12377_, _12376_, _12340_);
  or _57224_ (_12378_, _12377_, _12375_);
  or _57225_ (_12379_, _12378_, _12374_);
  and _57226_ (_12380_, _12379_, _12373_);
  or _57227_ (_12381_, _12380_, _12371_);
  and _57228_ (_12382_, _12381_, _12271_);
  or _57229_ (_12383_, _12382_, _12370_);
  and _57230_ (_12384_, _12383_, _12255_);
  or _57231_ (_12385_, _12384_, _12358_);
  and _57232_ (_39001_[1], _12385_, _38997_);
  and _57233_ (_12386_, _12316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not _57234_ (_12387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _57235_ (_12388_, _12181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _57236_ (_12389_, _12388_, _12387_);
  nor _57237_ (_12390_, _12177_, _12092_);
  nor _57238_ (_12391_, _12390_, _12162_);
  nand _57239_ (_12392_, _12391_, _12389_);
  or _57240_ (_12393_, _12163_, _12093_);
  and _57241_ (_12394_, _12393_, _12392_);
  or _57242_ (_12395_, _12394_, _12170_);
  or _57243_ (_12396_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _57244_ (_12397_, _12396_, _12274_);
  and _57245_ (_12398_, _12397_, _12286_);
  and _57246_ (_12399_, _12398_, _12395_);
  and _57247_ (_12400_, _12168_, _12093_);
  or _57248_ (_12401_, _12400_, _12165_);
  or _57249_ (_12402_, _12401_, _12399_);
  or _57250_ (_12403_, _12396_, _12166_);
  and _57251_ (_12404_, _12403_, _12185_);
  and _57252_ (_12405_, _12404_, _12402_);
  and _57253_ (_12406_, _12206_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _57254_ (_12407_, _12406_, _12387_);
  and _57255_ (_12408_, _12204_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _57256_ (_12409_, _12408_, _12209_);
  nand _57257_ (_12410_, _12409_, _12407_);
  or _57258_ (_12411_, _12210_, _12093_);
  and _57259_ (_12412_, _12411_, _12410_);
  or _57260_ (_12413_, _12412_, _12199_);
  or _57261_ (_12414_, _12396_, _12265_);
  and _57262_ (_12415_, _12414_, _12345_);
  and _57263_ (_12416_, _12415_, _12413_);
  and _57264_ (_12417_, _12197_, _12093_);
  or _57265_ (_12418_, _12417_, _12194_);
  or _57266_ (_12419_, _12418_, _12416_);
  and _57267_ (_12420_, _12396_, _12271_);
  or _57268_ (_12421_, _12420_, _12272_);
  and _57269_ (_12422_, _12421_, _12419_);
  or _57270_ (_12423_, _12422_, _12405_);
  and _57271_ (_12424_, _12423_, _12255_);
  or _57272_ (_12425_, _12424_, _12386_);
  and _57273_ (_39002_[0], _12425_, _38997_);
  and _57274_ (_12426_, _12316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or _57275_ (_12427_, _12388_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _57276_ (_12428_, _12427_, _12391_);
  and _57277_ (_12429_, _12162_, _12102_);
  or _57278_ (_12430_, _12429_, _12428_);
  and _57279_ (_12431_, _12430_, _12171_);
  not _57280_ (_12432_, _12171_);
  or _57281_ (_12433_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _57282_ (_12434_, _12433_, _12432_);
  or _57283_ (_12435_, _12434_, _12165_);
  or _57284_ (_12436_, _12435_, _12431_);
  or _57285_ (_12437_, _12166_, _12102_);
  and _57286_ (_12438_, _12437_, _12185_);
  and _57287_ (_12439_, _12438_, _12436_);
  and _57288_ (_12440_, _12194_, _12102_);
  and _57289_ (_12441_, _12433_, _12195_);
  or _57290_ (_12442_, _12441_, _12201_);
  and _57291_ (_12443_, _12209_, _12102_);
  or _57292_ (_12444_, _12406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _57293_ (_12445_, _12444_, _12409_);
  or _57294_ (_12446_, _12445_, _12375_);
  or _57295_ (_12447_, _12446_, _12443_);
  and _57296_ (_12448_, _12447_, _12442_);
  or _57297_ (_12449_, _12448_, _12440_);
  and _57298_ (_12450_, _12449_, _12271_);
  or _57299_ (_12451_, _12450_, _12439_);
  and _57300_ (_12452_, _12451_, _12255_);
  or _57301_ (_12453_, _12452_, _12426_);
  and _57302_ (_39002_[1], _12453_, _38997_);
  or _57303_ (_12454_, _12218_, _12213_);
  and _57304_ (_12455_, _12454_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or _57305_ (_12456_, _12455_, _12236_);
  and _57306_ (_39003_[0], _12456_, _38997_);
  and _57307_ (_12457_, _12214_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or _57308_ (_12458_, _12457_, _12188_);
  and _57309_ (_39004_[0], _12458_, _38997_);
  and _57310_ (_12459_, _12075_, _34229_);
  or _57311_ (_12460_, _12459_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _57312_ (_12461_, _12460_, _12086_);
  nand _57313_ (_12462_, _12459_, _35722_);
  and _57314_ (_12463_, _12462_, _12461_);
  and _57315_ (_12464_, _12078_, _34149_);
  or _57316_ (_12465_, _12464_, _12463_);
  and _57317_ (_39009_[0], _12465_, _38997_);
  and _57318_ (_12466_, _12075_, _11343_);
  or _57319_ (_12467_, _12466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _57320_ (_12468_, _12467_, _12086_);
  nand _57321_ (_12469_, _12466_, _35722_);
  and _57322_ (_12470_, _12469_, _12468_);
  and _57323_ (_12471_, _12078_, _34089_);
  or _57324_ (_12472_, _12471_, _12470_);
  and _57325_ (_39009_[1], _12472_, _38997_);
  and _57326_ (_12473_, _12075_, _11370_);
  or _57327_ (_12474_, _12473_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _57328_ (_12475_, _12474_, _12086_);
  nand _57329_ (_12476_, _12473_, _35722_);
  and _57330_ (_12477_, _12476_, _12475_);
  nor _57331_ (_12478_, _12086_, _34017_);
  or _57332_ (_12479_, _12478_, _12477_);
  and _57333_ (_39009_[2], _12479_, _38997_);
  and _57334_ (_12480_, _11366_, _33604_);
  and _57335_ (_12481_, _12480_, _34706_);
  and _57336_ (_12482_, _12481_, _12048_);
  and _57337_ (_12483_, _12482_, _34229_);
  or _57338_ (_12484_, _12483_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _57339_ (_12485_, _12484_, _12069_);
  nand _57340_ (_12486_, _12483_, _35722_);
  and _57341_ (_12487_, _12486_, _12485_);
  and _57342_ (_12488_, _12068_, _34149_);
  or _57343_ (_12489_, _12488_, _12487_);
  and _57344_ (_39010_[0], _12489_, _38997_);
  not _57345_ (_12490_, _33572_);
  nand _57346_ (_12491_, _12482_, _33644_);
  or _57347_ (_12492_, _12491_, _12490_);
  nor _57348_ (_12493_, _12492_, _35722_);
  and _57349_ (_12494_, _12492_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _57350_ (_12495_, _12494_, _12068_);
  or _57351_ (_12496_, _12495_, _12493_);
  or _57352_ (_12497_, _12069_, _34122_);
  and _57353_ (_12498_, _12497_, _38997_);
  and _57354_ (_39010_[1], _12498_, _12496_);
  nand _57355_ (_12499_, _12482_, _11359_);
  and _57356_ (_12500_, _12499_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _57357_ (_12501_, _12500_, _12068_);
  and _57358_ (_12502_, _34252_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _57359_ (_12503_, _12502_, _11345_);
  and _57360_ (_12504_, _12503_, _12063_);
  or _57361_ (_12505_, _12504_, _12501_);
  or _57362_ (_12506_, _12069_, _34089_);
  and _57363_ (_12507_, _12506_, _38997_);
  and _57364_ (_39010_[2], _12507_, _12505_);
  and _57365_ (_12508_, _12491_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _57366_ (_12509_, _12508_, _12068_);
  and _57367_ (_12510_, _11359_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _57368_ (_12511_, _12510_, _11357_);
  and _57369_ (_12512_, _12511_, _12063_);
  or _57370_ (_12513_, _12512_, _12509_);
  nand _57371_ (_12514_, _12068_, _34052_);
  and _57372_ (_12515_, _12514_, _38997_);
  and _57373_ (_39010_[3], _12515_, _12513_);
  not _57374_ (_12516_, _12482_);
  or _57375_ (_12517_, _12516_, _11372_);
  and _57376_ (_12518_, _12517_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _57377_ (_12519_, _12518_, _12068_);
  and _57378_ (_12520_, _11371_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _57379_ (_12521_, _12520_, _11376_);
  and _57380_ (_12522_, _12521_, _12063_);
  or _57381_ (_12523_, _12522_, _12519_);
  nand _57382_ (_12524_, _12068_, _34017_);
  and _57383_ (_12525_, _12524_, _38997_);
  and _57384_ (_39010_[4], _12525_, _12523_);
  nand _57385_ (_12526_, _12482_, _11383_);
  nor _57386_ (_12527_, _12526_, _35722_);
  and _57387_ (_12528_, _12526_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _57388_ (_12529_, _12528_, _12068_);
  or _57389_ (_12530_, _12529_, _12527_);
  or _57390_ (_12531_, _12069_, _33978_);
  and _57391_ (_12532_, _12531_, _38997_);
  and _57392_ (_39010_[5], _12532_, _12530_);
  nand _57393_ (_12533_, _12482_, _11392_);
  and _57394_ (_12534_, _12533_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or _57395_ (_12535_, _12534_, _12068_);
  nor _57396_ (_12536_, _12533_, _35722_);
  or _57397_ (_12537_, _12536_, _12535_);
  or _57398_ (_12538_, _12069_, _33942_);
  and _57399_ (_12539_, _12538_, _38997_);
  and _57400_ (_39010_[6], _12539_, _12537_);
  and _57401_ (_12540_, _12048_, _11368_);
  and _57402_ (_12541_, _12540_, _34229_);
  or _57403_ (_12542_, _12541_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _57404_ (_12543_, _12542_, _12055_);
  nand _57405_ (_12544_, _12541_, _35722_);
  and _57406_ (_12545_, _12544_, _12543_);
  and _57407_ (_12546_, _12054_, _34149_);
  or _57408_ (_12547_, _12546_, _12545_);
  and _57409_ (_39011_[0], _12547_, _38997_);
  nand _57410_ (_12548_, _12540_, _33644_);
  or _57411_ (_12549_, _12548_, _12490_);
  nor _57412_ (_12550_, _12549_, _35722_);
  and _57413_ (_12551_, _12052_, _11076_);
  and _57414_ (_12552_, _12551_, _33632_);
  and _57415_ (_12553_, _12549_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _57416_ (_12554_, _12553_, _12552_);
  or _57417_ (_12555_, _12554_, _12550_);
  or _57418_ (_12556_, _12055_, _34122_);
  and _57419_ (_12557_, _12556_, _38997_);
  and _57420_ (_39011_[1], _12557_, _12555_);
  nand _57421_ (_12558_, _12049_, _11359_);
  and _57422_ (_12559_, _12558_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _57423_ (_12560_, _12559_, _12054_);
  and _57424_ (_12561_, _34252_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _57425_ (_12562_, _12561_, _11345_);
  and _57426_ (_12563_, _12562_, _12049_);
  or _57427_ (_12564_, _12563_, _12560_);
  or _57428_ (_12565_, _12055_, _34089_);
  and _57429_ (_12566_, _12565_, _38997_);
  and _57430_ (_39011_[2], _12566_, _12564_);
  and _57431_ (_12567_, _12540_, _11357_);
  not _57432_ (_12568_, _11074_);
  or _57433_ (_12569_, _12548_, _12568_);
  and _57434_ (_12570_, _12569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _57435_ (_12571_, _12570_, _12552_);
  or _57436_ (_12572_, _12571_, _12567_);
  nand _57437_ (_12573_, _12054_, _34052_);
  and _57438_ (_12574_, _12573_, _38997_);
  and _57439_ (_39011_[3], _12574_, _12572_);
  not _57440_ (_12575_, _12049_);
  or _57441_ (_12576_, _12575_, _11372_);
  and _57442_ (_12577_, _12576_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _57443_ (_12578_, _12577_, _12054_);
  and _57444_ (_12579_, _11371_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _57445_ (_12580_, _12579_, _11376_);
  and _57446_ (_12581_, _12580_, _12049_);
  or _57447_ (_12582_, _12581_, _12578_);
  nand _57448_ (_12583_, _12054_, _34017_);
  and _57449_ (_12584_, _12583_, _38997_);
  and _57450_ (_39011_[4], _12584_, _12582_);
  and _57451_ (_12585_, _12049_, _11383_);
  or _57452_ (_12586_, _12585_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _57453_ (_12587_, _12586_, _12055_);
  nand _57454_ (_12588_, _12585_, _35722_);
  and _57455_ (_12589_, _12588_, _12587_);
  and _57456_ (_12590_, _12054_, _33978_);
  or _57457_ (_12591_, _12590_, _12589_);
  and _57458_ (_39011_[5], _12591_, _38997_);
  nand _57459_ (_12592_, _12540_, _11392_);
  and _57460_ (_12593_, _12592_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _57461_ (_12594_, _12593_, _12054_);
  nor _57462_ (_12595_, _12592_, _35722_);
  or _57463_ (_12596_, _12595_, _12594_);
  or _57464_ (_12597_, _12055_, _33942_);
  and _57465_ (_12598_, _12597_, _38997_);
  and _57466_ (_39011_[6], _12598_, _12596_);
  and _57467_ (_39029_, t2_i, _38997_);
  nor _57468_ (_12599_, t2_i, rst);
  and _57469_ (_39030_, _12599_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand _57470_ (_12600_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _38997_);
  nor _57471_ (_39031_, _12600_, t2ex_i);
  and _57472_ (_39032_, t2ex_i, _38997_);
  and _57473_ (_12601_, _34231_, _33605_);
  and _57474_ (_12602_, _12601_, _11524_);
  nand _57475_ (_12603_, _12602_, _34221_);
  and _57476_ (_12604_, _12601_, _11401_);
  not _57477_ (_12605_, _12604_);
  and _57478_ (_12606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _57479_ (_12607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _57480_ (_12608_, _12607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _57481_ (_12609_, _12608_, _12606_);
  not _57482_ (_12610_, _12609_);
  and _57483_ (_12611_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _57484_ (_12612_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _57485_ (_12613_, _12612_, _12611_);
  or _57486_ (_12614_, _12613_, _12602_);
  and _57487_ (_12615_, _12614_, _12605_);
  and _57488_ (_12616_, _12615_, _12603_);
  and _57489_ (_12617_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _57490_ (_12618_, _12617_, _12616_);
  and _57491_ (_39033_[7], _12618_, _38997_);
  nand _57492_ (_12619_, _12604_, _34221_);
  nor _57493_ (_12620_, _12610_, _12602_);
  or _57494_ (_12621_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not _57495_ (_12622_, _12620_);
  or _57496_ (_12623_, _12622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _57497_ (_12624_, _12623_, _12621_);
  or _57498_ (_12625_, _12624_, _12604_);
  and _57499_ (_12626_, _12625_, _38997_);
  and _57500_ (_39034_[7], _12626_, _12619_);
  not _57501_ (_12627_, _12607_);
  or _57502_ (_12628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _57503_ (_12629_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _57504_ (_12630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _12629_);
  and _57505_ (_12631_, _12630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _57506_ (_12632_, _12631_, _12628_);
  and _57507_ (_12633_, _12601_, _11425_);
  and _57508_ (_12634_, _12601_, _11486_);
  nor _57509_ (_12635_, _12634_, _12633_);
  and _57510_ (_12636_, _12635_, _12632_);
  and _57511_ (_12637_, _12636_, _12627_);
  or _57512_ (_12638_, _12637_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _57513_ (_12639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _57514_ (_12640_, _12639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _57515_ (_12641_, _12640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _57516_ (_12642_, _12641_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _57517_ (_12643_, _12642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _57518_ (_12644_, _12643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _57519_ (_12645_, _12644_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _57520_ (_12646_, _12645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _57521_ (_12647_, _12646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _57522_ (_12648_, _12647_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _57523_ (_12649_, _12648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _57524_ (_12650_, _12649_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _57525_ (_12651_, _12650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _57526_ (_12652_, _12651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _57527_ (_12653_, _12652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not _57528_ (_12654_, _12653_);
  nand _57529_ (_12655_, _12654_, _12637_);
  and _57530_ (_12656_, _12655_, _38997_);
  and _57531_ (_39035_, _12656_, _12638_);
  not _57532_ (_12657_, _12634_);
  nor _57533_ (_12658_, _12657_, _34221_);
  not _57534_ (_12659_, _12608_);
  and _57535_ (_12660_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _57536_ (_12661_, _12660_, _12632_);
  and _57537_ (_12662_, _12661_, _12653_);
  nand _57538_ (_12663_, _12644_, _12632_);
  nor _57539_ (_12664_, _12663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  not _57540_ (_12665_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand _57541_ (_12666_, _12606_, _12665_);
  nor _57542_ (_12667_, _12666_, _12627_);
  and _57543_ (_12668_, _12663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _57544_ (_12669_, _12668_, _12667_);
  or _57545_ (_12670_, _12669_, _12664_);
  or _57546_ (_12671_, _12670_, _12662_);
  not _57547_ (_12672_, _12667_);
  or _57548_ (_12673_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _57549_ (_12674_, _12673_, _12635_);
  and _57550_ (_12675_, _12674_, _12671_);
  and _57551_ (_12676_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _57552_ (_12677_, _12676_, _12675_);
  or _57553_ (_12678_, _12677_, _12658_);
  and _57554_ (_39036_[7], _12678_, _38997_);
  nand _57555_ (_12679_, _12633_, _34221_);
  and _57556_ (_12680_, _12667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _57557_ (_12681_, _12652_, _12632_);
  or _57558_ (_12682_, _12681_, _12680_);
  and _57559_ (_12683_, _12682_, _12657_);
  or _57560_ (_12684_, _12683_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _57561_ (_12685_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _57562_ (_12686_, _12685_, _12632_);
  nand _57563_ (_12687_, _12686_, _12653_);
  and _57564_ (_12688_, _12687_, _12672_);
  or _57565_ (_12689_, _12680_, _12634_);
  or _57566_ (_12690_, _12689_, _12688_);
  and _57567_ (_12691_, _12690_, _12684_);
  or _57568_ (_12692_, _12691_, _12633_);
  and _57569_ (_12693_, _12692_, _38997_);
  and _57570_ (_39037_[7], _12693_, _12679_);
  not _57571_ (_12694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  nor _57572_ (_12695_, _12635_, _12694_);
  and _57573_ (_12696_, _12666_, _12607_);
  and _57574_ (_12697_, _12696_, _12653_);
  and _57575_ (_12698_, _12697_, _12636_);
  or _57576_ (_12699_, _12698_, _12695_);
  and _57577_ (_39038_, _12699_, _38997_);
  or _57578_ (_12700_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  nor _57579_ (_12701_, _33630_, _34232_);
  and _57580_ (_12702_, _12701_, _12062_);
  or _57581_ (_12703_, _12702_, _12700_);
  not _57582_ (_12704_, _11075_);
  nor _57583_ (_12705_, _12704_, _35722_);
  nand _57584_ (_12706_, _12704_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _57585_ (_12707_, _12706_, _12702_);
  or _57586_ (_12708_, _12707_, _12705_);
  and _57587_ (_12709_, _12708_, _12703_);
  and _57588_ (_12710_, _12601_, _11091_);
  or _57589_ (_12711_, _12710_, _12709_);
  nand _57590_ (_12712_, _12710_, _34221_);
  and _57591_ (_12713_, _12712_, _38997_);
  and _57592_ (_39039_[7], _12713_, _12711_);
  or _57593_ (_12714_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _57594_ (_12715_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _57595_ (_12716_, _12715_, _12714_);
  or _57596_ (_12717_, _12716_, _12602_);
  nand _57597_ (_12718_, _12602_, _34148_);
  and _57598_ (_12719_, _12718_, _12717_);
  or _57599_ (_12720_, _12719_, _12604_);
  or _57600_ (_12721_, _12605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _57601_ (_12722_, _12721_, _38997_);
  and _57602_ (_39033_[0], _12722_, _12720_);
  not _57603_ (_12723_, _12602_);
  or _57604_ (_12724_, _12723_, _34122_);
  and _57605_ (_12725_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _57606_ (_12726_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _57607_ (_12727_, _12726_, _12725_);
  or _57608_ (_12728_, _12727_, _12602_);
  and _57609_ (_12729_, _12728_, _12605_);
  and _57610_ (_12730_, _12729_, _12724_);
  and _57611_ (_12731_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _57612_ (_12732_, _12731_, _12730_);
  and _57613_ (_39033_[1], _12732_, _38997_);
  or _57614_ (_12733_, _12723_, _34089_);
  and _57615_ (_12734_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _57616_ (_12735_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _57617_ (_12736_, _12735_, _12734_);
  or _57618_ (_12737_, _12736_, _12602_);
  and _57619_ (_12738_, _12737_, _12605_);
  and _57620_ (_12739_, _12738_, _12733_);
  and _57621_ (_12740_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _57622_ (_12741_, _12740_, _12739_);
  and _57623_ (_39033_[2], _12741_, _38997_);
  nand _57624_ (_12742_, _12602_, _34052_);
  and _57625_ (_12743_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _57626_ (_12744_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _57627_ (_12745_, _12744_, _12743_);
  or _57628_ (_12746_, _12745_, _12602_);
  and _57629_ (_12747_, _12746_, _12605_);
  and _57630_ (_12748_, _12747_, _12742_);
  and _57631_ (_12749_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _57632_ (_12750_, _12749_, _12748_);
  and _57633_ (_39033_[3], _12750_, _38997_);
  nand _57634_ (_12751_, _12602_, _34017_);
  and _57635_ (_12752_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _57636_ (_12753_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _57637_ (_12754_, _12753_, _12752_);
  or _57638_ (_12755_, _12754_, _12602_);
  and _57639_ (_12756_, _12755_, _12605_);
  and _57640_ (_12757_, _12756_, _12751_);
  and _57641_ (_12758_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _57642_ (_12759_, _12758_, _12757_);
  and _57643_ (_39033_[4], _12759_, _38997_);
  or _57644_ (_12760_, _12723_, _33978_);
  and _57645_ (_12761_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _57646_ (_12762_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _57647_ (_12763_, _12762_, _12761_);
  or _57648_ (_12764_, _12763_, _12602_);
  and _57649_ (_12765_, _12764_, _12605_);
  and _57650_ (_12766_, _12765_, _12760_);
  and _57651_ (_12767_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _57652_ (_12768_, _12767_, _12766_);
  and _57653_ (_39033_[5], _12768_, _38997_);
  or _57654_ (_12769_, _12723_, _33942_);
  not _57655_ (_12770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor _57656_ (_12771_, _12609_, _12770_);
  and _57657_ (_12772_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _57658_ (_12773_, _12772_, _12771_);
  or _57659_ (_12774_, _12773_, _12602_);
  and _57660_ (_12775_, _12774_, _12605_);
  and _57661_ (_12776_, _12775_, _12769_);
  and _57662_ (_12777_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _57663_ (_12778_, _12777_, _12776_);
  and _57664_ (_39033_[6], _12778_, _38997_);
  and _57665_ (_12779_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _57666_ (_12780_, _12622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or _57667_ (_12781_, _12780_, _12779_);
  or _57668_ (_12782_, _12781_, _12604_);
  nand _57669_ (_12783_, _12604_, _34148_);
  and _57670_ (_12784_, _12783_, _38997_);
  and _57671_ (_39034_[0], _12784_, _12782_);
  or _57672_ (_12785_, _12605_, _34122_);
  and _57673_ (_12786_, _12622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _57674_ (_12787_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _57675_ (_12788_, _12787_, _12786_);
  or _57676_ (_12789_, _12788_, _12604_);
  and _57677_ (_12790_, _12789_, _38997_);
  and _57678_ (_39034_[1], _12790_, _12785_);
  or _57679_ (_12791_, _12605_, _34089_);
  and _57680_ (_12792_, _12622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _57681_ (_12793_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _57682_ (_12794_, _12793_, _12792_);
  or _57683_ (_12795_, _12794_, _12604_);
  and _57684_ (_12796_, _12795_, _38997_);
  and _57685_ (_39034_[2], _12796_, _12791_);
  nand _57686_ (_12797_, _12604_, _34052_);
  not _57687_ (_12798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor _57688_ (_12799_, _12620_, _12798_);
  and _57689_ (_12800_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _57690_ (_12801_, _12800_, _12799_);
  or _57691_ (_12802_, _12801_, _12604_);
  and _57692_ (_12803_, _12802_, _38997_);
  and _57693_ (_39034_[3], _12803_, _12797_);
  nand _57694_ (_12804_, _12604_, _34017_);
  not _57695_ (_12805_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor _57696_ (_12806_, _12620_, _12805_);
  and _57697_ (_12807_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _57698_ (_12808_, _12807_, _12806_);
  or _57699_ (_12809_, _12808_, _12604_);
  and _57700_ (_12810_, _12809_, _38997_);
  and _57701_ (_39034_[4], _12810_, _12804_);
  or _57702_ (_12811_, _12605_, _33978_);
  or _57703_ (_12812_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  not _57704_ (_12813_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nand _57705_ (_12814_, _12620_, _12813_);
  and _57706_ (_12815_, _12814_, _12812_);
  or _57707_ (_12816_, _12815_, _12604_);
  and _57708_ (_12817_, _12816_, _38997_);
  and _57709_ (_39034_[5], _12817_, _12811_);
  or _57710_ (_12818_, _12605_, _33942_);
  not _57711_ (_12819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor _57712_ (_12820_, _12620_, _12819_);
  and _57713_ (_12821_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _57714_ (_12822_, _12821_, _12820_);
  or _57715_ (_12823_, _12822_, _12604_);
  and _57716_ (_12824_, _12823_, _38997_);
  and _57717_ (_39034_[6], _12824_, _12818_);
  or _57718_ (_12825_, _12632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _57719_ (_12826_, _12632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  not _57720_ (_12827_, _12826_);
  and _57721_ (_12828_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _57722_ (_12829_, _12828_, _12653_);
  or _57723_ (_12830_, _12829_, _12827_);
  and _57724_ (_12831_, _12830_, _12825_);
  or _57725_ (_12832_, _12831_, _12667_);
  or _57726_ (_12833_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _57727_ (_12834_, _12833_, _12635_);
  and _57728_ (_12835_, _12834_, _12832_);
  and _57729_ (_12836_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _57730_ (_12837_, _12634_, _34149_);
  or _57731_ (_12838_, _12837_, _12836_);
  or _57732_ (_12839_, _12838_, _12835_);
  and _57733_ (_39036_[0], _12839_, _38997_);
  nor _57734_ (_12840_, _12827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _57735_ (_12841_, _12827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _57736_ (_12842_, _12841_, _12667_);
  or _57737_ (_12843_, _12842_, _12840_);
  and _57738_ (_12844_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _57739_ (_12845_, _12844_, _12632_);
  and _57740_ (_12846_, _12845_, _12653_);
  or _57741_ (_12847_, _12846_, _12843_);
  or _57742_ (_12848_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _57743_ (_12849_, _12848_, _12635_);
  and _57744_ (_12850_, _12849_, _12847_);
  and _57745_ (_12851_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _57746_ (_12852_, _12634_, _34122_);
  or _57747_ (_12853_, _12852_, _12851_);
  or _57748_ (_12854_, _12853_, _12850_);
  and _57749_ (_39036_[1], _12854_, _38997_);
  and _57750_ (_12855_, _12634_, _34089_);
  and _57751_ (_12856_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _57752_ (_12857_, _12653_, _12632_);
  and _57753_ (_12858_, _12857_, _12856_);
  nand _57754_ (_12859_, _12639_, _12632_);
  and _57755_ (_12860_, _12859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor _57756_ (_12861_, _12859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _57757_ (_12862_, _12861_, _12667_);
  or _57758_ (_12863_, _12862_, _12860_);
  or _57759_ (_12864_, _12863_, _12858_);
  or _57760_ (_12865_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _57761_ (_12866_, _12865_, _12635_);
  and _57762_ (_12867_, _12866_, _12864_);
  and _57763_ (_12868_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _57764_ (_12869_, _12868_, _12867_);
  or _57765_ (_12870_, _12869_, _12855_);
  and _57766_ (_39036_[2], _12870_, _38997_);
  nor _57767_ (_12871_, _12657_, _34052_);
  and _57768_ (_12872_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _57769_ (_12873_, _12872_, _12857_);
  nand _57770_ (_12874_, _12640_, _12632_);
  and _57771_ (_12875_, _12874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _57772_ (_12876_, _12874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _57773_ (_12877_, _12876_, _12667_);
  or _57774_ (_12878_, _12877_, _12875_);
  or _57775_ (_12879_, _12878_, _12873_);
  or _57776_ (_12880_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _57777_ (_12881_, _12880_, _12635_);
  and _57778_ (_12882_, _12881_, _12879_);
  and _57779_ (_12883_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _57780_ (_12884_, _12883_, _12882_);
  or _57781_ (_12885_, _12884_, _12871_);
  and _57782_ (_39036_[3], _12885_, _38997_);
  nor _57783_ (_12886_, _12657_, _34017_);
  and _57784_ (_12887_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _57785_ (_12888_, _12887_, _12857_);
  nand _57786_ (_12889_, _12641_, _12632_);
  and _57787_ (_12890_, _12889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor _57788_ (_12891_, _12889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _57789_ (_12892_, _12891_, _12667_);
  or _57790_ (_12893_, _12892_, _12890_);
  or _57791_ (_12894_, _12893_, _12888_);
  or _57792_ (_12895_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _57793_ (_12896_, _12895_, _12635_);
  and _57794_ (_12897_, _12896_, _12894_);
  and _57795_ (_12898_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _57796_ (_12899_, _12898_, _12897_);
  or _57797_ (_12900_, _12899_, _12886_);
  and _57798_ (_39036_[4], _12900_, _38997_);
  and _57799_ (_12901_, _12634_, _33978_);
  and _57800_ (_12902_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _57801_ (_12903_, _12902_, _12857_);
  nand _57802_ (_12904_, _12642_, _12632_);
  and _57803_ (_12905_, _12904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _57804_ (_12906_, _12904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _57805_ (_12907_, _12906_, _12667_);
  or _57806_ (_12908_, _12907_, _12905_);
  or _57807_ (_12909_, _12908_, _12903_);
  or _57808_ (_12910_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _57809_ (_12911_, _12910_, _12635_);
  and _57810_ (_12912_, _12911_, _12909_);
  and _57811_ (_12913_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _57812_ (_12914_, _12913_, _12912_);
  or _57813_ (_12915_, _12914_, _12901_);
  and _57814_ (_39036_[5], _12915_, _38997_);
  and _57815_ (_12916_, _12634_, _33942_);
  nor _57816_ (_12917_, _12608_, _12770_);
  and _57817_ (_12918_, _12917_, _12857_);
  and _57818_ (_12919_, _12643_, _12632_);
  or _57819_ (_12920_, _12919_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _57820_ (_12921_, _12920_, _12663_);
  or _57821_ (_12922_, _12921_, _12667_);
  or _57822_ (_12923_, _12922_, _12918_);
  nand _57823_ (_12924_, _12667_, _12770_);
  and _57824_ (_12925_, _12924_, _12635_);
  and _57825_ (_12926_, _12925_, _12923_);
  and _57826_ (_12927_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _57827_ (_12928_, _12927_, _12926_);
  or _57828_ (_12929_, _12928_, _12916_);
  and _57829_ (_39036_[6], _12929_, _38997_);
  and _57830_ (_12930_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _57831_ (_12931_, _12930_, _12857_);
  and _57832_ (_12932_, _12645_, _12632_);
  or _57833_ (_12933_, _12932_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _57834_ (_12934_, _12932_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _57835_ (_12935_, _12934_, _12933_);
  or _57836_ (_12936_, _12935_, _12667_);
  or _57837_ (_12937_, _12936_, _12931_);
  or _57838_ (_12938_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _57839_ (_12939_, _12938_, _12635_);
  and _57840_ (_12940_, _12939_, _12937_);
  and _57841_ (_12941_, _12634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _57842_ (_12942_, _12633_, _34149_);
  or _57843_ (_12943_, _12942_, _12941_);
  or _57844_ (_12944_, _12943_, _12940_);
  and _57845_ (_39037_[0], _12944_, _38997_);
  nor _57846_ (_12945_, _33657_, _33644_);
  and _57847_ (_12946_, _12945_, _33572_);
  and _57848_ (_12947_, _12601_, _12946_);
  and _57849_ (_12948_, _12947_, _33662_);
  not _57850_ (_12949_, _12948_);
  and _57851_ (_12950_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _57852_ (_12951_, _12950_, _12857_);
  and _57853_ (_12952_, _12646_, _12632_);
  or _57854_ (_12953_, _12952_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand _57855_ (_12954_, _12952_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _57856_ (_12955_, _12954_, _12953_);
  or _57857_ (_12956_, _12955_, _12667_);
  or _57858_ (_12957_, _12956_, _12951_);
  nor _57859_ (_12958_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _57860_ (_12959_, _12958_, _12634_);
  and _57861_ (_12960_, _12959_, _12957_);
  and _57862_ (_12961_, _12945_, _34228_);
  and _57863_ (_12962_, _12601_, _12961_);
  and _57864_ (_12963_, _12962_, _33662_);
  and _57865_ (_12964_, _12963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _57866_ (_12965_, _12964_, _12960_);
  and _57867_ (_12966_, _12965_, _12949_);
  and _57868_ (_12967_, _12948_, _34122_);
  or _57869_ (_12968_, _12967_, _12966_);
  and _57870_ (_39037_[1], _12968_, _38997_);
  and _57871_ (_12969_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _57872_ (_12970_, _12969_, _12857_);
  and _57873_ (_12971_, _12647_, _12632_);
  or _57874_ (_12972_, _12971_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand _57875_ (_12973_, _12971_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _57876_ (_12974_, _12973_, _12972_);
  or _57877_ (_12975_, _12974_, _12667_);
  or _57878_ (_12976_, _12975_, _12970_);
  nor _57879_ (_12977_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _57880_ (_12978_, _12977_, _12634_);
  and _57881_ (_12979_, _12978_, _12976_);
  and _57882_ (_12980_, _12963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _57883_ (_12981_, _12980_, _12979_);
  and _57884_ (_12982_, _12981_, _12949_);
  and _57885_ (_12983_, _12948_, _34089_);
  or _57886_ (_12984_, _12983_, _12982_);
  and _57887_ (_39037_[2], _12984_, _38997_);
  nor _57888_ (_12985_, _12608_, _12798_);
  and _57889_ (_12986_, _12985_, _12857_);
  nor _57890_ (_12987_, _12973_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _57891_ (_12988_, _12973_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _57892_ (_12989_, _12988_, _12667_);
  or _57893_ (_12990_, _12989_, _12987_);
  or _57894_ (_12991_, _12990_, _12986_);
  not _57895_ (_12992_, _12635_);
  and _57896_ (_12993_, _12667_, _12798_);
  nor _57897_ (_12994_, _12993_, _12992_);
  and _57898_ (_12995_, _12994_, _12991_);
  and _57899_ (_12996_, _12634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _57900_ (_12997_, _12996_, _12995_);
  nor _57901_ (_12998_, _12949_, _34052_);
  or _57902_ (_12999_, _12998_, _12997_);
  and _57903_ (_39037_[3], _12999_, _38997_);
  nor _57904_ (_13000_, _12608_, _12805_);
  and _57905_ (_13001_, _13000_, _12857_);
  nand _57906_ (_13002_, _12649_, _12632_);
  nor _57907_ (_13003_, _13002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _57908_ (_13004_, _13002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _57909_ (_13005_, _13004_, _12667_);
  or _57910_ (_13006_, _13005_, _13003_);
  or _57911_ (_13007_, _13006_, _13001_);
  nand _57912_ (_13008_, _12667_, _12805_);
  and _57913_ (_13009_, _13008_, _12635_);
  and _57914_ (_13010_, _13009_, _13007_);
  and _57915_ (_13011_, _12634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _57916_ (_13012_, _13011_, _13010_);
  nor _57917_ (_13013_, _12949_, _34017_);
  or _57918_ (_13014_, _13013_, _13012_);
  and _57919_ (_39037_[4], _13014_, _38997_);
  and _57920_ (_13015_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _57921_ (_13016_, _13015_, _12857_);
  and _57922_ (_13017_, _12650_, _12632_);
  nor _57923_ (_13018_, _13017_, _12813_);
  and _57924_ (_13019_, _13017_, _12813_);
  or _57925_ (_13020_, _13019_, _12667_);
  or _57926_ (_13021_, _13020_, _13018_);
  or _57927_ (_13022_, _13021_, _13016_);
  or _57928_ (_13023_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _57929_ (_13024_, _13023_, _12635_);
  and _57930_ (_13025_, _13024_, _13022_);
  and _57931_ (_13026_, _12634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _57932_ (_13027_, _13026_, _13025_);
  and _57933_ (_13028_, _12633_, _33978_);
  or _57934_ (_13029_, _13028_, _13027_);
  and _57935_ (_39037_[5], _13029_, _38997_);
  and _57936_ (_13030_, _12634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _57937_ (_13031_, _12608_, _12819_);
  and _57938_ (_13032_, _13031_, _12857_);
  and _57939_ (_13033_, _12651_, _12632_);
  nor _57940_ (_13034_, _13033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _57941_ (_13035_, _13034_, _12681_);
  or _57942_ (_13036_, _13035_, _12667_);
  or _57943_ (_13037_, _13036_, _13032_);
  and _57944_ (_13038_, _12667_, _12819_);
  nor _57945_ (_13039_, _13038_, _12992_);
  and _57946_ (_13040_, _13039_, _13037_);
  or _57947_ (_13041_, _13040_, _13030_);
  and _57948_ (_13042_, _12633_, _33942_);
  or _57949_ (_13043_, _13042_, _13041_);
  and _57950_ (_39037_[6], _13043_, _38997_);
  nand _57951_ (_13044_, _12701_, _12481_);
  or _57952_ (_13045_, _13044_, _11314_);
  nor _57953_ (_13046_, _13045_, _35722_);
  and _57954_ (_13047_, _13045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or _57955_ (_13048_, _13047_, _12710_);
  or _57956_ (_13049_, _13048_, _13046_);
  nand _57957_ (_13050_, _12710_, _34148_);
  and _57958_ (_13051_, _13050_, _38997_);
  and _57959_ (_39039_[0], _13051_, _13049_);
  not _57960_ (_13052_, _12710_);
  and _57961_ (_13053_, _12702_, _34253_);
  or _57962_ (_13054_, _13053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _57963_ (_13055_, _13054_, _13052_);
  nand _57964_ (_13056_, _13053_, _35722_);
  and _57965_ (_13057_, _13056_, _13055_);
  and _57966_ (_13058_, _12710_, _34122_);
  or _57967_ (_13059_, _13058_, _13057_);
  and _57968_ (_39039_[1], _13059_, _38997_);
  or _57969_ (_13060_, _13044_, _11358_);
  and _57970_ (_13061_, _13060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _57971_ (_13062_, _13061_, _12710_);
  and _57972_ (_13063_, _34252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _57973_ (_13064_, _13063_, _11345_);
  and _57974_ (_13065_, _13064_, _12702_);
  or _57975_ (_13066_, _13065_, _13062_);
  or _57976_ (_13067_, _13052_, _34089_);
  and _57977_ (_13068_, _13067_, _38997_);
  and _57978_ (_39039_[2], _13068_, _13066_);
  or _57979_ (_13069_, _13044_, _11073_);
  and _57980_ (_13070_, _13069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _57981_ (_13071_, _13070_, _12710_);
  and _57982_ (_13072_, _11359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _57983_ (_13073_, _13072_, _11357_);
  and _57984_ (_13074_, _13073_, _12702_);
  or _57985_ (_13075_, _13074_, _13071_);
  nand _57986_ (_13076_, _12710_, _34052_);
  and _57987_ (_13077_, _13076_, _38997_);
  and _57988_ (_39039_[3], _13077_, _13075_);
  or _57989_ (_13078_, _13044_, _11372_);
  and _57990_ (_13079_, _13078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _57991_ (_13080_, _13079_, _12710_);
  and _57992_ (_13081_, _11371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _57993_ (_13082_, _13081_, _11376_);
  and _57994_ (_13083_, _13082_, _12702_);
  or _57995_ (_13084_, _13083_, _13080_);
  nand _57996_ (_13085_, _12710_, _34017_);
  and _57997_ (_13086_, _13085_, _38997_);
  and _57998_ (_39039_[4], _13086_, _13084_);
  and _57999_ (_13087_, _12702_, _11383_);
  or _58000_ (_13088_, _13087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _58001_ (_13089_, _13088_, _13052_);
  nand _58002_ (_13090_, _13087_, _35722_);
  and _58003_ (_13091_, _13090_, _13089_);
  and _58004_ (_13092_, _12710_, _33978_);
  or _58005_ (_13093_, _13092_, _13091_);
  and _58006_ (_39039_[5], _13093_, _38997_);
  and _58007_ (_13094_, _12606_, _12694_);
  or _58008_ (_13095_, _13094_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _58009_ (_13096_, _13095_, _12702_);
  not _58010_ (_13097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _58011_ (_13098_, _11392_, _13097_);
  nand _58012_ (_13099_, _13098_, _12702_);
  or _58013_ (_13100_, _13099_, _12080_);
  and _58014_ (_13101_, _13100_, _13096_);
  or _58015_ (_13102_, _13101_, _12710_);
  or _58016_ (_13103_, _13052_, _33942_);
  and _58017_ (_13104_, _13103_, _38997_);
  and _58018_ (_39039_[6], _13104_, _13102_);
  and _58019_ (_13105_, _33657_, _33604_);
  and _58020_ (_13106_, _13105_, _34706_);
  and _58021_ (_13107_, _13106_, _11081_);
  and _58022_ (_13108_, _11075_, _13107_);
  nand _58023_ (_13109_, _13108_, _35722_);
  or _58024_ (_13110_, _13108_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _58025_ (_13111_, _13110_, _11083_);
  and _58026_ (_13112_, _13111_, _13109_);
  and _58027_ (_13113_, _34257_, _33633_);
  nand _58028_ (_13114_, _13113_, _34221_);
  or _58029_ (_13115_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _58030_ (_13116_, _13115_, _33662_);
  and _58031_ (_13117_, _13116_, _13114_);
  not _58032_ (_13118_, _33661_);
  and _58033_ (_13119_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _58034_ (_13120_, _13119_, rst);
  or _58035_ (_13121_, _13120_, _13117_);
  or _58036_ (_39012_[7], _13121_, _13112_);
  nor _58037_ (_13122_, _34251_, _33604_);
  and _58038_ (_13123_, _13122_, _34706_);
  and _58039_ (_13124_, _13123_, _11081_);
  and _58040_ (_13125_, _13124_, _11075_);
  nand _58041_ (_13126_, _13125_, _35722_);
  or _58042_ (_13127_, _13125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _58043_ (_13128_, _13127_, _11083_);
  and _58044_ (_13129_, _13128_, _13126_);
  and _58045_ (_13130_, _11011_, _34257_);
  nand _58046_ (_13131_, _13130_, _34221_);
  or _58047_ (_13132_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _58048_ (_13133_, _13132_, _33662_);
  and _58049_ (_13134_, _13133_, _13131_);
  and _58050_ (_13135_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _58051_ (_13136_, _13135_, rst);
  or _58052_ (_13137_, _13136_, _13134_);
  or _58053_ (_39013_[7], _13137_, _13129_);
  and _58054_ (_13138_, _12048_, _13106_);
  and _58055_ (_13139_, _13138_, _11075_);
  nand _58056_ (_13140_, _13139_, _35722_);
  or _58057_ (_13141_, _13139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _58058_ (_13142_, _13141_, _11083_);
  and _58059_ (_13143_, _13142_, _13140_);
  and _58060_ (_13144_, _12067_, _34257_);
  nand _58061_ (_13145_, _13144_, _34221_);
  or _58062_ (_13146_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _58063_ (_13147_, _13146_, _33662_);
  and _58064_ (_13148_, _13147_, _13145_);
  and _58065_ (_13149_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _58066_ (_13150_, _13149_, rst);
  or _58067_ (_13151_, _13150_, _13148_);
  or _58068_ (_39014_[7], _13151_, _13143_);
  and _58069_ (_13152_, _13123_, _12048_);
  and _58070_ (_13153_, _13152_, _11075_);
  nand _58071_ (_13154_, _13153_, _35722_);
  or _58072_ (_13155_, _13153_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _58073_ (_13156_, _13155_, _11083_);
  and _58074_ (_13157_, _13156_, _13154_);
  and _58075_ (_13158_, _12052_, _34257_);
  and _58076_ (_13159_, _13158_, _33632_);
  nand _58077_ (_13160_, _13159_, _34221_);
  or _58078_ (_13161_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _58079_ (_13162_, _13161_, _33662_);
  and _58080_ (_13163_, _13162_, _13160_);
  and _58081_ (_13164_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _58082_ (_13165_, _13164_, rst);
  or _58083_ (_13166_, _13165_, _13163_);
  or _58084_ (_39015_[7], _13166_, _13157_);
  nand _58085_ (_13167_, _13113_, _35722_);
  or _58086_ (_13168_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _58087_ (_13169_, _13168_, _11083_);
  and _58088_ (_13170_, _13169_, _13167_);
  nand _58089_ (_13171_, _13113_, _34148_);
  and _58090_ (_13172_, _13168_, _33662_);
  and _58091_ (_13173_, _13172_, _13171_);
  and _58092_ (_13174_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or _58093_ (_13175_, _13174_, rst);
  or _58094_ (_13176_, _13175_, _13173_);
  or _58095_ (_39012_[0], _13176_, _13170_);
  and _58096_ (_13177_, _34259_, _33633_);
  nand _58097_ (_13178_, _35722_, _13177_);
  or _58098_ (_13179_, _13177_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _58099_ (_13180_, _13179_, _11083_);
  and _58100_ (_13181_, _13180_, _13178_);
  not _58101_ (_13182_, _13113_);
  or _58102_ (_13183_, _13182_, _34122_);
  or _58103_ (_13184_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _58104_ (_13185_, _13184_, _33662_);
  and _58105_ (_13186_, _13185_, _13183_);
  and _58106_ (_13187_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _58107_ (_13188_, _13187_, rst);
  or _58108_ (_13189_, _13188_, _13186_);
  or _58109_ (_39012_[1], _13189_, _13181_);
  not _58110_ (_13190_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _58111_ (_13191_, _11359_, _13107_);
  nor _58112_ (_13192_, _13191_, _13190_);
  and _58113_ (_13193_, _34252_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _58114_ (_13194_, _13193_, _11345_);
  and _58115_ (_13195_, _13194_, _13107_);
  or _58116_ (_13196_, _13195_, _13192_);
  and _58117_ (_13197_, _13196_, _11083_);
  or _58118_ (_13198_, _13182_, _34089_);
  or _58119_ (_13199_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _58120_ (_13200_, _13199_, _33662_);
  and _58121_ (_13201_, _13200_, _13198_);
  nor _58122_ (_13202_, _33661_, _13190_);
  or _58123_ (_13203_, _13202_, rst);
  or _58124_ (_13204_, _13203_, _13201_);
  or _58125_ (_39012_[2], _13204_, _13197_);
  and _58126_ (_13205_, _11356_, _13107_);
  nand _58127_ (_13206_, _13205_, _35722_);
  or _58128_ (_13207_, _13205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _58129_ (_13208_, _13207_, _11083_);
  and _58130_ (_13209_, _13208_, _13206_);
  nand _58131_ (_13210_, _13113_, _34052_);
  or _58132_ (_13211_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _58133_ (_13212_, _13211_, _33662_);
  and _58134_ (_13213_, _13212_, _13210_);
  and _58135_ (_13214_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _58136_ (_13215_, _13214_, rst);
  or _58137_ (_13216_, _13215_, _13213_);
  or _58138_ (_39012_[3], _13216_, _13209_);
  not _58139_ (_13217_, _13107_);
  or _58140_ (_13218_, _11372_, _13217_);
  and _58141_ (_13219_, _13218_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _58142_ (_13220_, _11371_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _58143_ (_13221_, _13220_, _11376_);
  and _58144_ (_13222_, _13221_, _13107_);
  or _58145_ (_13223_, _13222_, _13219_);
  and _58146_ (_13224_, _13223_, _11083_);
  nand _58147_ (_13225_, _13113_, _34017_);
  or _58148_ (_13226_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _58149_ (_13227_, _13226_, _33662_);
  and _58150_ (_13228_, _13227_, _13225_);
  and _58151_ (_13229_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _58152_ (_13230_, _13229_, rst);
  or _58153_ (_13231_, _13230_, _13228_);
  or _58154_ (_39012_[4], _13231_, _13224_);
  and _58155_ (_13232_, _11383_, _13107_);
  nand _58156_ (_13233_, _13232_, _35722_);
  or _58157_ (_13234_, _13232_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _58158_ (_13235_, _13234_, _11083_);
  and _58159_ (_13236_, _13235_, _13233_);
  or _58160_ (_13237_, _13182_, _33978_);
  or _58161_ (_13238_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _58162_ (_13239_, _13238_, _33662_);
  and _58163_ (_13240_, _13239_, _13237_);
  and _58164_ (_13241_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _58165_ (_13242_, _13241_, rst);
  or _58166_ (_13243_, _13242_, _13240_);
  or _58167_ (_39012_[5], _13243_, _13236_);
  nand _58168_ (_13244_, _11392_, _13107_);
  or _58169_ (_13245_, _13244_, _35723_);
  not _58170_ (_13246_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nand _58171_ (_13247_, _13244_, _13246_);
  and _58172_ (_13248_, _13247_, _11083_);
  and _58173_ (_13249_, _13248_, _13245_);
  or _58174_ (_13250_, _13182_, _33942_);
  or _58175_ (_13251_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _58176_ (_13252_, _13251_, _33662_);
  and _58177_ (_13253_, _13252_, _13250_);
  nor _58178_ (_13254_, _33661_, _13246_);
  or _58179_ (_13255_, _13254_, rst);
  or _58180_ (_13256_, _13255_, _13253_);
  or _58181_ (_39012_[6], _13256_, _13249_);
  nand _58182_ (_13257_, _13130_, _35722_);
  or _58183_ (_13258_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _58184_ (_13259_, _13258_, _11083_);
  and _58185_ (_13260_, _13259_, _13257_);
  nand _58186_ (_13261_, _13130_, _34148_);
  and _58187_ (_13262_, _13258_, _33662_);
  and _58188_ (_13263_, _13262_, _13261_);
  and _58189_ (_13264_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or _58190_ (_13265_, _13264_, rst);
  or _58191_ (_13266_, _13265_, _13263_);
  or _58192_ (_39013_[0], _13266_, _13260_);
  and _58193_ (_13267_, _13124_, _34253_);
  nand _58194_ (_13268_, _13267_, _35722_);
  or _58195_ (_13269_, _13267_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _58196_ (_13270_, _13269_, _11083_);
  and _58197_ (_13271_, _13270_, _13268_);
  not _58198_ (_13272_, _13130_);
  or _58199_ (_13273_, _13272_, _34122_);
  or _58200_ (_13274_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _58201_ (_13275_, _13274_, _33662_);
  and _58202_ (_13276_, _13275_, _13273_);
  and _58203_ (_13277_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _58204_ (_13278_, _13277_, rst);
  or _58205_ (_13279_, _13278_, _13276_);
  or _58206_ (_39013_[1], _13279_, _13271_);
  and _58207_ (_13280_, _13124_, _11343_);
  nand _58208_ (_13281_, _13280_, _35722_);
  or _58209_ (_13282_, _13280_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _58210_ (_13283_, _13282_, _11083_);
  and _58211_ (_13284_, _13283_, _13281_);
  or _58212_ (_13285_, _13272_, _34089_);
  or _58213_ (_13286_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _58214_ (_13287_, _13286_, _33662_);
  and _58215_ (_13288_, _13287_, _13285_);
  and _58216_ (_13289_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _58217_ (_13290_, _13289_, rst);
  or _58218_ (_13291_, _13290_, _13288_);
  or _58219_ (_39013_[2], _13291_, _13284_);
  and _58220_ (_13292_, _13124_, _11356_);
  nand _58221_ (_13293_, _13292_, _35722_);
  or _58222_ (_13294_, _13292_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _58223_ (_13295_, _13294_, _11083_);
  and _58224_ (_13296_, _13295_, _13293_);
  nand _58225_ (_13297_, _13130_, _34052_);
  or _58226_ (_13298_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _58227_ (_13299_, _13298_, _33662_);
  and _58228_ (_13300_, _13299_, _13297_);
  and _58229_ (_13301_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _58230_ (_13302_, _13301_, rst);
  or _58231_ (_13303_, _13302_, _13300_);
  or _58232_ (_39013_[3], _13303_, _13296_);
  and _58233_ (_13304_, _13124_, _11370_);
  nand _58234_ (_13305_, _13304_, _35722_);
  or _58235_ (_13306_, _13304_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _58236_ (_13307_, _13306_, _11083_);
  and _58237_ (_13308_, _13307_, _13305_);
  nand _58238_ (_13309_, _13130_, _34017_);
  or _58239_ (_13310_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _58240_ (_13311_, _13310_, _33662_);
  and _58241_ (_13312_, _13311_, _13309_);
  and _58242_ (_13313_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _58243_ (_13314_, _13313_, rst);
  or _58244_ (_13315_, _13314_, _13312_);
  or _58245_ (_39013_[4], _13315_, _13308_);
  and _58246_ (_13316_, _13124_, _11383_);
  nand _58247_ (_13317_, _13316_, _35722_);
  or _58248_ (_13318_, _13316_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _58249_ (_13319_, _13318_, _11083_);
  and _58250_ (_13320_, _13319_, _13317_);
  or _58251_ (_13321_, _13272_, _33978_);
  or _58252_ (_13322_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _58253_ (_13323_, _13322_, _33662_);
  and _58254_ (_13324_, _13323_, _13321_);
  and _58255_ (_13325_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _58256_ (_13326_, _13325_, rst);
  or _58257_ (_13327_, _13326_, _13324_);
  or _58258_ (_39013_[5], _13327_, _13320_);
  nand _58259_ (_13328_, _13124_, _11392_);
  or _58260_ (_13329_, _13328_, _35723_);
  not _58261_ (_13330_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nand _58262_ (_13331_, _13328_, _13330_);
  and _58263_ (_13332_, _13331_, _11083_);
  and _58264_ (_13333_, _13332_, _13329_);
  or _58265_ (_13334_, _13272_, _33942_);
  or _58266_ (_13335_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _58267_ (_13336_, _13335_, _33662_);
  and _58268_ (_13337_, _13336_, _13334_);
  nor _58269_ (_13338_, _33661_, _13330_);
  or _58270_ (_13339_, _13338_, rst);
  or _58271_ (_13340_, _13339_, _13337_);
  or _58272_ (_39013_[6], _13340_, _13333_);
  and _58273_ (_13341_, _13138_, _34229_);
  nand _58274_ (_13342_, _13341_, _35722_);
  or _58275_ (_13343_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _58276_ (_13344_, _13343_, _11083_);
  and _58277_ (_13345_, _13344_, _13342_);
  nand _58278_ (_13346_, _13144_, _34148_);
  and _58279_ (_13347_, _13343_, _33662_);
  and _58280_ (_13348_, _13347_, _13346_);
  and _58281_ (_13349_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _58282_ (_13350_, _13349_, rst);
  or _58283_ (_13351_, _13350_, _13348_);
  or _58284_ (_39014_[0], _13351_, _13345_);
  and _58285_ (_13352_, _13138_, _34253_);
  nand _58286_ (_13353_, _13352_, _35722_);
  or _58287_ (_13354_, _13352_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _58288_ (_13355_, _13354_, _11083_);
  and _58289_ (_13356_, _13355_, _13353_);
  not _58290_ (_13357_, _13144_);
  or _58291_ (_13358_, _13357_, _34122_);
  or _58292_ (_13359_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _58293_ (_13360_, _13359_, _33662_);
  and _58294_ (_13361_, _13360_, _13358_);
  and _58295_ (_13362_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _58296_ (_13363_, _13362_, rst);
  or _58297_ (_13364_, _13363_, _13361_);
  or _58298_ (_39014_[1], _13364_, _13356_);
  and _58299_ (_13365_, _13138_, _11343_);
  nand _58300_ (_13366_, _13365_, _35722_);
  or _58301_ (_13367_, _13365_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _58302_ (_13368_, _13367_, _11083_);
  and _58303_ (_13369_, _13368_, _13366_);
  or _58304_ (_13370_, _13357_, _34089_);
  or _58305_ (_13371_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _58306_ (_13372_, _13371_, _33662_);
  and _58307_ (_13373_, _13372_, _13370_);
  and _58308_ (_13374_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _58309_ (_13375_, _13374_, rst);
  or _58310_ (_13376_, _13375_, _13373_);
  or _58311_ (_39014_[2], _13376_, _13369_);
  and _58312_ (_13377_, _13138_, _11356_);
  nand _58313_ (_13378_, _13377_, _35722_);
  or _58314_ (_13379_, _13377_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _58315_ (_13380_, _13379_, _11083_);
  and _58316_ (_13381_, _13380_, _13378_);
  nand _58317_ (_13382_, _13144_, _34052_);
  or _58318_ (_13383_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _58319_ (_13384_, _13383_, _33662_);
  and _58320_ (_13385_, _13384_, _13382_);
  and _58321_ (_13386_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _58322_ (_13387_, _13386_, rst);
  or _58323_ (_13388_, _13387_, _13385_);
  or _58324_ (_39014_[3], _13388_, _13381_);
  and _58325_ (_13389_, _13138_, _11370_);
  nand _58326_ (_13390_, _13389_, _35722_);
  or _58327_ (_13391_, _13389_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _58328_ (_13392_, _13391_, _11083_);
  and _58329_ (_13393_, _13392_, _13390_);
  nand _58330_ (_13394_, _13144_, _34017_);
  or _58331_ (_13395_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _58332_ (_13396_, _13395_, _33662_);
  and _58333_ (_13397_, _13396_, _13394_);
  and _58334_ (_13398_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _58335_ (_13399_, _13398_, rst);
  or _58336_ (_13400_, _13399_, _13397_);
  or _58337_ (_39014_[4], _13400_, _13393_);
  and _58338_ (_13401_, _13138_, _11383_);
  nand _58339_ (_13402_, _13401_, _35722_);
  or _58340_ (_13403_, _13401_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _58341_ (_13404_, _13403_, _11083_);
  and _58342_ (_13405_, _13404_, _13402_);
  or _58343_ (_13406_, _13357_, _33978_);
  or _58344_ (_13407_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _58345_ (_13408_, _13407_, _33662_);
  and _58346_ (_13409_, _13408_, _13406_);
  and _58347_ (_13410_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _58348_ (_13411_, _13410_, rst);
  or _58349_ (_13412_, _13411_, _13409_);
  or _58350_ (_39014_[5], _13412_, _13405_);
  nand _58351_ (_13413_, _13138_, _11392_);
  or _58352_ (_13414_, _13413_, _35723_);
  not _58353_ (_13415_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nand _58354_ (_13416_, _13413_, _13415_);
  and _58355_ (_13417_, _13416_, _11083_);
  and _58356_ (_13418_, _13417_, _13414_);
  or _58357_ (_13419_, _13357_, _33942_);
  or _58358_ (_13420_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _58359_ (_13421_, _13420_, _33662_);
  and _58360_ (_13422_, _13421_, _13419_);
  nor _58361_ (_13423_, _33661_, _13415_);
  or _58362_ (_13424_, _13423_, rst);
  or _58363_ (_13425_, _13424_, _13422_);
  or _58364_ (_39014_[6], _13425_, _13418_);
  and _58365_ (_13426_, _13152_, _34229_);
  nand _58366_ (_13427_, _13426_, _35722_);
  or _58367_ (_13428_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _58368_ (_13429_, _13428_, _11083_);
  and _58369_ (_13430_, _13429_, _13427_);
  nand _58370_ (_13431_, _13159_, _34148_);
  and _58371_ (_13432_, _13428_, _33662_);
  and _58372_ (_13433_, _13432_, _13431_);
  and _58373_ (_13434_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _58374_ (_13435_, _13434_, rst);
  or _58375_ (_13436_, _13435_, _13433_);
  or _58376_ (_39015_[0], _13436_, _13430_);
  and _58377_ (_13437_, _13152_, _34253_);
  nand _58378_ (_13438_, _13437_, _35722_);
  or _58379_ (_13439_, _13437_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _58380_ (_13440_, _13439_, _11083_);
  and _58381_ (_13441_, _13440_, _13438_);
  not _58382_ (_13442_, _13159_);
  or _58383_ (_13443_, _13442_, _34122_);
  or _58384_ (_13444_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _58385_ (_13445_, _13444_, _33662_);
  and _58386_ (_13446_, _13445_, _13443_);
  and _58387_ (_13447_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _58388_ (_13448_, _13447_, rst);
  or _58389_ (_13449_, _13448_, _13446_);
  or _58390_ (_39015_[1], _13449_, _13441_);
  and _58391_ (_13450_, _13152_, _11343_);
  nand _58392_ (_13451_, _13450_, _35722_);
  or _58393_ (_13452_, _13450_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _58394_ (_13453_, _13452_, _11083_);
  and _58395_ (_13454_, _13453_, _13451_);
  or _58396_ (_13455_, _13442_, _34089_);
  or _58397_ (_13456_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _58398_ (_13457_, _13456_, _33662_);
  and _58399_ (_13458_, _13457_, _13455_);
  and _58400_ (_13459_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _58401_ (_13460_, _13459_, rst);
  or _58402_ (_13461_, _13460_, _13458_);
  or _58403_ (_39015_[2], _13461_, _13454_);
  and _58404_ (_13462_, _13152_, _11356_);
  nand _58405_ (_13463_, _13462_, _35722_);
  or _58406_ (_13464_, _13462_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _58407_ (_13465_, _13464_, _11083_);
  and _58408_ (_13466_, _13465_, _13463_);
  nand _58409_ (_13467_, _13159_, _34052_);
  or _58410_ (_13468_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _58411_ (_13469_, _13468_, _33662_);
  and _58412_ (_13470_, _13469_, _13467_);
  and _58413_ (_13471_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _58414_ (_13472_, _13471_, rst);
  or _58415_ (_13473_, _13472_, _13470_);
  or _58416_ (_39015_[3], _13473_, _13466_);
  and _58417_ (_13474_, _13152_, _11370_);
  nand _58418_ (_13475_, _13474_, _35722_);
  or _58419_ (_13476_, _13474_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _58420_ (_13477_, _13476_, _11083_);
  and _58421_ (_13478_, _13477_, _13475_);
  nand _58422_ (_13479_, _13159_, _34017_);
  or _58423_ (_13480_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _58424_ (_13481_, _13480_, _33662_);
  and _58425_ (_13482_, _13481_, _13479_);
  and _58426_ (_13483_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _58427_ (_13484_, _13483_, rst);
  or _58428_ (_13485_, _13484_, _13482_);
  or _58429_ (_39015_[4], _13485_, _13478_);
  and _58430_ (_13486_, _13152_, _11383_);
  nand _58431_ (_13487_, _13486_, _35722_);
  or _58432_ (_13488_, _13486_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _58433_ (_13489_, _13488_, _11083_);
  and _58434_ (_13490_, _13489_, _13487_);
  or _58435_ (_13491_, _13442_, _33978_);
  or _58436_ (_13492_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _58437_ (_13493_, _13492_, _33662_);
  and _58438_ (_13494_, _13493_, _13491_);
  and _58439_ (_13495_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _58440_ (_13496_, _13495_, rst);
  or _58441_ (_13497_, _13496_, _13494_);
  or _58442_ (_39015_[5], _13497_, _13490_);
  nand _58443_ (_13498_, _13152_, _11392_);
  or _58444_ (_13499_, _13498_, _35723_);
  not _58445_ (_13500_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nand _58446_ (_13501_, _13498_, _13500_);
  and _58447_ (_13502_, _13501_, _11083_);
  and _58448_ (_13503_, _13502_, _13499_);
  or _58449_ (_13504_, _13442_, _33942_);
  or _58450_ (_13505_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _58451_ (_13506_, _13505_, _33662_);
  and _58452_ (_13507_, _13506_, _13504_);
  nor _58453_ (_13508_, _33661_, _13500_);
  or _58454_ (_13509_, _13508_, rst);
  or _58455_ (_13510_, _13509_, _13507_);
  or _58456_ (_39015_[6], _13510_, _13503_);
  and _58457_ (_13511_, _12701_, _11083_);
  and _58458_ (_13512_, _13511_, _13123_);
  not _58459_ (_13513_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _58460_ (_13514_, _11075_, _13513_);
  or _58461_ (_13515_, _13514_, _12705_);
  and _58462_ (_13516_, _13515_, _13512_);
  nor _58463_ (_13517_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _58464_ (_13518_, _13517_);
  nand _58465_ (_13519_, _13518_, _35722_);
  and _58466_ (_13520_, _13517_, _13513_);
  nor _58467_ (_13521_, _13520_, _13512_);
  and _58468_ (_13522_, _13521_, _13519_);
  or _58469_ (_13523_, _13522_, _34235_);
  or _58470_ (_13524_, _13523_, _13516_);
  nand _58471_ (_13525_, _34235_, _34221_);
  and _58472_ (_13526_, _13525_, _38997_);
  and _58473_ (_39016_[6], _13526_, _13524_);
  and _58474_ (_13527_, _34235_, _34122_);
  and _58475_ (_13528_, _13512_, _34253_);
  nand _58476_ (_13529_, _13528_, _35722_);
  or _58477_ (_13530_, _13528_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _58478_ (_13531_, _13530_, _34236_);
  and _58479_ (_13532_, _13531_, _13529_);
  or _58480_ (_13533_, _13532_, _13527_);
  and _58481_ (_39016_[0], _13533_, _38997_);
  and _58482_ (_13534_, _33930_, _33673_);
  not _58483_ (_13535_, _13534_);
  nor _58484_ (_13536_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _58485_ (_13537_, _13536_);
  and _58486_ (_13538_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not _58487_ (_13539_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _58488_ (_13540_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _13539_);
  not _58489_ (_13541_, _13540_);
  or _58490_ (_13542_, _13541_, _33987_);
  not _58491_ (_13543_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _58492_ (_13544_, _13543_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _58493_ (_13545_, _13544_);
  or _58494_ (_13546_, _13545_, _35601_);
  and _58495_ (_13547_, _13546_, _13542_);
  nor _58496_ (_13548_, _13544_, _13540_);
  or _58497_ (_13549_, _34131_, _13539_);
  nand _58498_ (_13550_, _13549_, _13548_);
  nand _58499_ (_13551_, _13550_, _13547_);
  nand _58500_ (_13552_, _13536_, _33778_);
  and _58501_ (_13553_, _13552_, _13551_);
  and _58502_ (_13554_, _13553_, _33815_);
  or _58503_ (_13555_, _13541_, _33951_);
  or _58504_ (_13556_, _13545_, _34035_);
  and _58505_ (_13557_, _13556_, _13555_);
  or _58506_ (_13558_, _34098_, _13539_);
  nand _58507_ (_13559_, _13558_, _13548_);
  nand _58508_ (_13560_, _13559_, _13557_);
  nand _58509_ (_13561_, _13536_, _34196_);
  and _58510_ (_13562_, _13561_, _13560_);
  and _58511_ (_13563_, _13562_, _33884_);
  and _58512_ (_13564_, _13563_, _13554_);
  and _58513_ (_13565_, _13553_, _33884_);
  and _58514_ (_13566_, _13562_, _33798_);
  nand _58515_ (_13567_, _13566_, _13565_);
  and _58516_ (_13568_, _13553_, _33798_);
  or _58517_ (_13569_, _13568_, _13563_);
  and _58518_ (_13570_, _13569_, _13567_);
  and _58519_ (_13571_, _13570_, _13564_);
  or _58520_ (_13572_, _13567_, _33765_);
  and _58521_ (_13573_, _13553_, _33766_);
  not _58522_ (_13574_, _13573_);
  nand _58523_ (_13575_, _13574_, _13567_);
  and _58524_ (_13576_, _13575_, _13566_);
  nand _58525_ (_13577_, _13576_, _13572_);
  or _58526_ (_13578_, _13573_, _13566_);
  and _58527_ (_13579_, _13578_, _13577_);
  and _58528_ (_13580_, _13579_, _13571_);
  not _58529_ (_13581_, _13576_);
  nand _58530_ (_13582_, _13561_, _13560_);
  or _58531_ (_13583_, _13582_, _33765_);
  nand _58532_ (_13584_, _13552_, _13551_);
  or _58533_ (_13585_, _13584_, _34180_);
  or _58534_ (_13586_, _13585_, _13583_);
  nand _58535_ (_13587_, _13585_, _13583_);
  and _58536_ (_13588_, _13587_, _13586_);
  nand _58537_ (_13589_, _13588_, _13581_);
  or _58538_ (_13590_, _13588_, _13581_);
  nand _58539_ (_13591_, _13590_, _13589_);
  nand _58540_ (_13592_, _13591_, _13580_);
  not _58541_ (_13593_, _33831_);
  and _58542_ (_13594_, _13562_, _13593_);
  and _58543_ (_13595_, _13553_, _33865_);
  nand _58544_ (_13596_, _13595_, _13594_);
  or _58545_ (_13597_, _13584_, _33831_);
  and _58546_ (_13598_, _13562_, _33865_);
  and _58547_ (_13599_, _13598_, _13597_);
  nand _58548_ (_13600_, _13599_, _13554_);
  nand _58549_ (_13601_, _13600_, _13596_);
  not _58550_ (_13602_, _13564_);
  and _58551_ (_13603_, _13562_, _33815_);
  or _58552_ (_13604_, _13603_, _13565_);
  and _58553_ (_13605_, _13604_, _13602_);
  nand _58554_ (_13606_, _13605_, _13601_);
  not _58555_ (_13607_, _13606_);
  not _58556_ (_13608_, _13571_);
  or _58557_ (_13609_, _13570_, _13564_);
  and _58558_ (_13610_, _13609_, _13608_);
  and _58559_ (_13611_, _13610_, _13607_);
  nand _58560_ (_13612_, _13579_, _13571_);
  or _58561_ (_13613_, _13579_, _13571_);
  and _58562_ (_13614_, _13613_, _13612_);
  nand _58563_ (_13615_, _13614_, _13611_);
  not _58564_ (_13616_, _13615_);
  or _58565_ (_13617_, _13591_, _13580_);
  and _58566_ (_13618_, _13617_, _13592_);
  nand _58567_ (_13619_, _13618_, _13616_);
  and _58568_ (_13620_, _13619_, _13592_);
  and _58569_ (_13621_, _13553_, _35711_);
  and _58570_ (_13622_, _13621_, _13594_);
  or _58571_ (_13623_, _13595_, _13594_);
  and _58572_ (_13624_, _13623_, _13596_);
  and _58573_ (_13625_, _13624_, _13622_);
  or _58574_ (_13626_, _13599_, _13554_);
  and _58575_ (_13627_, _13626_, _13600_);
  nand _58576_ (_13628_, _13627_, _13625_);
  not _58577_ (_13629_, _13628_);
  or _58578_ (_13630_, _13605_, _13601_);
  and _58579_ (_13631_, _13630_, _13606_);
  nand _58580_ (_13632_, _13631_, _13629_);
  not _58581_ (_13633_, _13632_);
  nand _58582_ (_13634_, _13610_, _13607_);
  or _58583_ (_13635_, _13610_, _13607_);
  and _58584_ (_13636_, _13635_, _13634_);
  nand _58585_ (_13637_, _13636_, _13633_);
  not _58586_ (_13638_, _13637_);
  or _58587_ (_13639_, _13614_, _13611_);
  and _58588_ (_13640_, _13639_, _13615_);
  and _58589_ (_13641_, _13618_, _13640_);
  nand _58590_ (_13642_, _13641_, _13638_);
  nand _58591_ (_13643_, _13642_, _13620_);
  and _58592_ (_13644_, _13562_, _35707_);
  and _58593_ (_13645_, _13644_, _13574_);
  and _58594_ (_13646_, _13588_, _13576_);
  and _58595_ (_13647_, _13646_, _13645_);
  nor _58596_ (_13648_, _13646_, _13645_);
  nor _58597_ (_13649_, _13648_, _13647_);
  nand _58598_ (_13650_, _13649_, _13643_);
  not _58599_ (_13651_, _13647_);
  and _58600_ (_13652_, _13651_, _13586_);
  nand _58601_ (_13653_, _13652_, _13650_);
  nand _58602_ (_13654_, _13653_, _13538_);
  and _58603_ (_13655_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  or _58604_ (_13656_, _13649_, _13643_);
  and _58605_ (_13657_, _13656_, _13650_);
  nand _58606_ (_13658_, _13657_, _13655_);
  or _58607_ (_13659_, _13653_, _13538_);
  nand _58608_ (_13660_, _13659_, _13654_);
  or _58609_ (_13661_, _13660_, _13658_);
  nand _58610_ (_13662_, _13661_, _13654_);
  and _58611_ (_13663_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _58612_ (_13664_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _58613_ (_13665_, _13664_, _13663_);
  and _58614_ (_13666_, _13665_, _13662_);
  and _58615_ (_13667_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  nand _58616_ (_13668_, _13640_, _13638_);
  nand _58617_ (_13669_, _13668_, _13615_);
  nand _58618_ (_13670_, _13618_, _13669_);
  or _58619_ (_13671_, _13618_, _13669_);
  and _58620_ (_13672_, _13671_, _13670_);
  nand _58621_ (_13673_, _13672_, _13667_);
  or _58622_ (_13674_, _13672_, _13667_);
  nand _58623_ (_13675_, _13674_, _13673_);
  and _58624_ (_13676_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or _58625_ (_13677_, _13640_, _13638_);
  and _58626_ (_13678_, _13677_, _13668_);
  nand _58627_ (_13679_, _13678_, _13676_);
  or _58628_ (_13680_, _13678_, _13676_);
  and _58629_ (_13681_, _13680_, _13679_);
  and _58630_ (_13682_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  or _58631_ (_13683_, _13636_, _13633_);
  and _58632_ (_13684_, _13683_, _13637_);
  nand _58633_ (_13685_, _13684_, _13682_);
  or _58634_ (_13686_, _13684_, _13682_);
  nand _58635_ (_13687_, _13686_, _13685_);
  and _58636_ (_13688_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or _58637_ (_13689_, _13631_, _13629_);
  and _58638_ (_13690_, _13689_, _13632_);
  nand _58639_ (_13691_, _13690_, _13688_);
  and _58640_ (_13692_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or _58641_ (_13693_, _13627_, _13625_);
  and _58642_ (_13694_, _13693_, _13628_);
  nand _58643_ (_13695_, _13694_, _13692_);
  and _58644_ (_13696_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand _58645_ (_13697_, _13624_, _13622_);
  or _58646_ (_13698_, _13624_, _13622_);
  and _58647_ (_13699_, _13698_, _13697_);
  and _58648_ (_13700_, _13699_, _13696_);
  not _58649_ (_13701_, _13700_);
  or _58650_ (_13702_, _13694_, _13692_);
  nand _58651_ (_13703_, _13702_, _13695_);
  or _58652_ (_13704_, _13703_, _13701_);
  and _58653_ (_13705_, _13704_, _13695_);
  or _58654_ (_13706_, _13690_, _13688_);
  nand _58655_ (_13707_, _13706_, _13691_);
  or _58656_ (_13708_, _13707_, _13705_);
  and _58657_ (_13709_, _13708_, _13691_);
  or _58658_ (_13710_, _13709_, _13687_);
  nand _58659_ (_13711_, _13710_, _13685_);
  nand _58660_ (_13712_, _13711_, _13681_);
  and _58661_ (_13713_, _13712_, _13679_);
  or _58662_ (_13714_, _13713_, _13675_);
  and _58663_ (_13715_, _13714_, _13673_);
  or _58664_ (_13716_, _13657_, _13655_);
  and _58665_ (_13717_, _13716_, _13658_);
  and _58666_ (_13718_, _13659_, _13654_);
  and _58667_ (_13719_, _13718_, _13717_);
  nand _58668_ (_13720_, _13665_, _13719_);
  nor _58669_ (_13721_, _13720_, _13715_);
  or _58670_ (_13722_, _13721_, _13666_);
  and _58671_ (_13723_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _58672_ (_13724_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _58673_ (_13725_, _13724_, _13723_);
  and _58674_ (_13726_, _13725_, _13722_);
  and _58675_ (_13727_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and _58676_ (_13728_, _13727_, _13726_);
  and _58677_ (_13729_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor _58678_ (_13730_, _13729_, _13728_);
  and _58679_ (_13731_, _13728_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  or _58680_ (_13732_, _13731_, _13730_);
  or _58681_ (_13733_, _13732_, _13535_);
  nor _58682_ (_13734_, _13727_, _13726_);
  nor _58683_ (_13735_, _13734_, _13728_);
  and _58684_ (_13736_, _13723_, _13722_);
  nor _58685_ (_13737_, _13724_, _13736_);
  nor _58686_ (_13738_, _13737_, _13726_);
  not _58687_ (_13739_, _13717_);
  or _58688_ (_13740_, _13739_, _13715_);
  not _58689_ (_13741_, _13740_);
  and _58690_ (_13742_, _13739_, _13715_);
  nor _58691_ (_13743_, _13742_, _13741_);
  and _58692_ (_13744_, _13740_, _13658_);
  or _58693_ (_13745_, _13660_, _13744_);
  nand _58694_ (_13746_, _13660_, _13744_);
  and _58695_ (_13747_, _13746_, _13745_);
  or _58696_ (_13748_, _13747_, _13743_);
  nand _58697_ (_13749_, _13745_, _13654_);
  nand _58698_ (_13750_, _13749_, _13663_);
  or _58699_ (_13751_, _13749_, _13663_);
  and _58700_ (_13752_, _13751_, _13750_);
  or _58701_ (_13753_, _13752_, _13748_);
  nor _58702_ (_13754_, _13723_, _13722_);
  nor _58703_ (_13755_, _13754_, _13736_);
  or _58704_ (_13756_, _13755_, _13753_);
  or _58705_ (_13757_, _13756_, _13738_);
  or _58706_ (_13758_, _13757_, _13735_);
  and _58707_ (_13759_, _13758_, _13534_);
  or _58708_ (_13760_, _35634_, _35632_);
  not _58709_ (_13761_, _35584_);
  nand _58710_ (_13762_, _35632_, _13761_);
  and _58711_ (_13763_, _13762_, _35582_);
  and _58712_ (_13764_, _13763_, _13760_);
  not _58713_ (_13765_, _35672_);
  nor _58714_ (_13766_, _13765_, _35670_);
  and _58715_ (_13767_, _13765_, _35670_);
  or _58716_ (_13768_, _13767_, _13766_);
  and _58717_ (_13769_, _13768_, _35637_);
  nor _58718_ (_13770_, _34131_, _34098_);
  and _58719_ (_13771_, _35601_, _34035_);
  and _58720_ (_13772_, _13771_, _13770_);
  and _58721_ (_13773_, _33778_, _34196_);
  and _58722_ (_13774_, _33921_, _33913_);
  and _58723_ (_13775_, _33987_, _33951_);
  and _58724_ (_13776_, _13775_, _13774_);
  and _58725_ (_13777_, _13776_, _13773_);
  nand _58726_ (_13778_, _13777_, _13772_);
  nand _58727_ (_13779_, _13778_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _58728_ (_13780_, _13779_, _13769_);
  nor _58729_ (_13781_, _13780_, _13764_);
  not _58730_ (_13782_, _13664_);
  and _58731_ (_13783_, _13782_, _13750_);
  nor _58732_ (_13784_, _13783_, _13722_);
  nand _58733_ (_13785_, _13784_, _13534_);
  nand _58734_ (_13786_, _13785_, _13781_);
  nor _58735_ (_13787_, _13786_, _13759_);
  nand _58736_ (_13788_, _13787_, _13733_);
  nor _58737_ (_13789_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _58738_ (_13790_, _13789_, _13512_);
  and _58739_ (_13791_, _13790_, _13788_);
  and _58740_ (_13792_, _11344_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _58741_ (_13793_, _13792_, _11345_);
  and _58742_ (_13794_, _13793_, _13512_);
  or _58743_ (_13795_, _13794_, _34235_);
  or _58744_ (_13796_, _13795_, _13791_);
  or _58745_ (_13797_, _34236_, _34089_);
  and _58746_ (_13798_, _13797_, _38997_);
  and _58747_ (_39016_[1], _13798_, _13796_);
  and _58748_ (_13799_, _13512_, _11356_);
  nand _58749_ (_13800_, _13799_, _35722_);
  or _58750_ (_13801_, _13799_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _58751_ (_13802_, _13801_, _34236_);
  and _58752_ (_13803_, _13802_, _13800_);
  or _58753_ (_13804_, _13803_, _34282_);
  and _58754_ (_39016_[2], _13804_, _38997_);
  and _58755_ (_13805_, _13512_, _11370_);
  nand _58756_ (_13806_, _13805_, _35722_);
  or _58757_ (_13807_, _13805_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _58758_ (_13808_, _13807_, _34236_);
  and _58759_ (_13809_, _13808_, _13806_);
  or _58760_ (_13810_, _13809_, _34238_);
  and _58761_ (_39016_[3], _13810_, _38997_);
  and _58762_ (_13811_, _34235_, _33978_);
  and _58763_ (_13812_, _13512_, _11383_);
  nand _58764_ (_13813_, _13812_, _35722_);
  or _58765_ (_13814_, _13812_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _58766_ (_13815_, _13814_, _34236_);
  and _58767_ (_13816_, _13815_, _13813_);
  or _58768_ (_13817_, _13816_, _13811_);
  and _58769_ (_39016_[4], _13817_, _38997_);
  and _58770_ (_13818_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _58771_ (_13819_, _13818_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _58772_ (_13820_, _35628_, _35582_);
  and _58773_ (_13821_, _35658_, _35637_);
  nand _58774_ (_13822_, _33935_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _58775_ (_13823_, _13822_, _13818_);
  or _58776_ (_13824_, _13823_, _13821_);
  or _58777_ (_13825_, _13824_, _13820_);
  and _58778_ (_13826_, _13825_, _13819_);
  or _58779_ (_13827_, _13826_, _13512_);
  not _58780_ (_13828_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _58781_ (_13829_, _11392_, _13828_);
  nand _58782_ (_13830_, _13829_, _13512_);
  or _58783_ (_13831_, _13830_, _12080_);
  and _58784_ (_13832_, _13831_, _13827_);
  or _58785_ (_13833_, _13832_, _34235_);
  or _58786_ (_13834_, _34236_, _33942_);
  and _58787_ (_13835_, _13834_, _38997_);
  and _58788_ (_39016_[5], _13835_, _13833_);
  nand _58789_ (_13836_, _11074_, _33665_);
  not _58790_ (_13837_, _13774_);
  nor _58791_ (_13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _58792_ (_13839_, _13838_, _34180_);
  nor _58793_ (_13840_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not _58794_ (_13841_, _13840_);
  and _58795_ (_13842_, _13841_, _13839_);
  not _58796_ (_13843_, _13842_);
  or _58797_ (_13844_, _34131_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _58798_ (_13845_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _58799_ (_13846_, _34062_, _13845_);
  and _58800_ (_13847_, _13846_, _13844_);
  or _58801_ (_13848_, _13847_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _58802_ (_13849_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _58803_ (_13850_, _34007_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _58804_ (_13851_, _33778_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _58805_ (_13852_, _13851_, _13850_);
  or _58806_ (_13853_, _13852_, _13849_);
  and _58807_ (_13854_, _13853_, _13848_);
  nor _58808_ (_13855_, _13854_, _13843_);
  and _58809_ (_13856_, _13854_, _13843_);
  nand _58810_ (_13857_, _13838_, _33765_);
  nor _58811_ (_13858_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not _58812_ (_13859_, _13858_);
  and _58813_ (_13860_, _13859_, _13857_);
  not _58814_ (_13861_, _13860_);
  and _58815_ (_13862_, _34098_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _58816_ (_13863_, _13862_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _58817_ (_13864_, _34035_, _13845_);
  nand _58818_ (_13865_, _33951_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _58819_ (_13866_, _13865_, _13864_);
  or _58820_ (_13867_, _13866_, _13849_);
  and _58821_ (_13868_, _13867_, _13863_);
  or _58822_ (_13869_, _13868_, _13861_);
  nor _58823_ (_13870_, _13869_, _13856_);
  nor _58824_ (_13871_, _13870_, _13855_);
  nor _58825_ (_13872_, _13856_, _13855_);
  nand _58826_ (_13873_, _13868_, _13861_);
  and _58827_ (_13874_, _13873_, _13869_);
  and _58828_ (_13875_, _13874_, _13872_);
  nand _58829_ (_13876_, _13838_, _33797_);
  nor _58830_ (_13877_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not _58831_ (_13878_, _13877_);
  and _58832_ (_13879_, _13878_, _13876_);
  and _58833_ (_13880_, _34131_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _58834_ (_13881_, _13880_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _58835_ (_13882_, _34062_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _58836_ (_13883_, _34007_, _13845_);
  and _58837_ (_13884_, _13883_, _13882_);
  or _58838_ (_13885_, _13884_, _13849_);
  nand _58839_ (_13886_, _13885_, _13881_);
  and _58840_ (_13887_, _13886_, _13879_);
  not _58841_ (_13888_, _13887_);
  or _58842_ (_13889_, _34098_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _58843_ (_13890_, _34035_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _58844_ (_13891_, _13890_, _13889_);
  and _58845_ (_13892_, _13891_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _58846_ (_13893_, _13892_);
  nand _58847_ (_13894_, _13838_, _33883_);
  nor _58848_ (_13895_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not _58849_ (_13896_, _13895_);
  and _58850_ (_13897_, _13896_, _13894_);
  and _58851_ (_13898_, _13897_, _13893_);
  not _58852_ (_13899_, _13898_);
  nor _58853_ (_13900_, _13886_, _13879_);
  or _58854_ (_13901_, _13900_, _13887_);
  or _58855_ (_13902_, _13901_, _13899_);
  nand _58856_ (_13903_, _13902_, _13888_);
  nand _58857_ (_13904_, _13903_, _13875_);
  and _58858_ (_13905_, _13904_, _13871_);
  and _58859_ (_13906_, _13847_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _58860_ (_13907_, _13906_);
  nor _58861_ (_13908_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not _58862_ (_13909_, _13908_);
  nand _58863_ (_13910_, _13838_, _33814_);
  and _58864_ (_13911_, _13910_, _13909_);
  nand _58865_ (_13912_, _13911_, _13907_);
  or _58866_ (_13913_, _13911_, _13907_);
  nand _58867_ (_13914_, _13913_, _13912_);
  and _58868_ (_13915_, _13862_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _58869_ (_13916_, _13915_);
  not _58870_ (_13917_, _13838_);
  or _58871_ (_13918_, _13917_, _33865_);
  nor _58872_ (_13919_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not _58873_ (_13920_, _13919_);
  and _58874_ (_13921_, _13920_, _13918_);
  nand _58875_ (_13922_, _13921_, _13916_);
  and _58876_ (_13923_, _13880_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _58877_ (_13924_, _13923_);
  nand _58878_ (_13925_, _13838_, _33831_);
  nor _58879_ (_13926_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not _58880_ (_13927_, _13926_);
  and _58881_ (_13928_, _13927_, _13925_);
  nor _58882_ (_13929_, _13928_, _13924_);
  or _58883_ (_13930_, _13921_, _13916_);
  nand _58884_ (_13931_, _13930_, _13922_);
  or _58885_ (_13932_, _13931_, _13929_);
  and _58886_ (_13933_, _13932_, _13922_);
  or _58887_ (_13934_, _13933_, _13914_);
  nand _58888_ (_13935_, _13934_, _13912_);
  or _58889_ (_13936_, _13897_, _13893_);
  and _58890_ (_13937_, _13936_, _13899_);
  not _58891_ (_13938_, _13901_);
  and _58892_ (_13939_, _13938_, _13937_);
  and _58893_ (_13940_, _13939_, _13875_);
  nand _58894_ (_13941_, _13940_, _13935_);
  nand _58895_ (_13942_, _13941_, _13905_);
  nor _58896_ (_13943_, _13891_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _58897_ (_13944_, _33951_, _13845_);
  and _58898_ (_13945_, _34196_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _58899_ (_13946_, _13945_, _13944_);
  nor _58900_ (_13947_, _13946_, _13849_);
  nor _58901_ (_13948_, _13947_, _13943_);
  not _58902_ (_13949_, _13948_);
  nor _58903_ (_13950_, _13773_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _58904_ (_13951_, _13866_, _13852_);
  nor _58905_ (_13952_, _13946_, _13884_);
  and _58906_ (_13953_, _13952_, _13951_);
  nor _58907_ (_13954_, _13953_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _58908_ (_13955_, _13954_, _13950_);
  and _58909_ (_13956_, _13955_, _13949_);
  and _58910_ (_13957_, _13956_, _13942_);
  nor _58911_ (_13958_, _13957_, _13843_);
  not _58912_ (_13959_, _13874_);
  and _58913_ (_13960_, _13937_, _13935_);
  nor _58914_ (_13961_, _13960_, _13898_);
  or _58915_ (_13962_, _13961_, _13900_);
  and _58916_ (_13963_, _13962_, _13888_);
  or _58917_ (_13964_, _13963_, _13959_);
  and _58918_ (_13965_, _13964_, _13869_);
  nand _58919_ (_13966_, _13965_, _13872_);
  or _58920_ (_13967_, _13965_, _13872_);
  nand _58921_ (_13968_, _13967_, _13966_);
  and _58922_ (_13969_, _13968_, _13957_);
  nor _58923_ (_13970_, _13969_, _13958_);
  not _58924_ (_13971_, _13854_);
  and _58925_ (_13972_, _13963_, _13959_);
  not _58926_ (_13973_, _13972_);
  nand _58927_ (_13974_, _13973_, _13964_);
  nand _58928_ (_13975_, _13974_, _13957_);
  nor _58929_ (_13976_, _13957_, _13860_);
  not _58930_ (_13977_, _13976_);
  and _58931_ (_13978_, _13977_, _13975_);
  nand _58932_ (_13979_, _13978_, _13971_);
  or _58933_ (_13980_, _13978_, _13971_);
  and _58934_ (_13981_, _13980_, _13979_);
  not _58935_ (_13982_, _13868_);
  nand _58936_ (_13983_, _13901_, _13961_);
  or _58937_ (_13984_, _13901_, _13961_);
  nand _58938_ (_13985_, _13984_, _13983_);
  nand _58939_ (_13986_, _13985_, _13957_);
  nor _58940_ (_13987_, _13957_, _13879_);
  not _58941_ (_13988_, _13987_);
  and _58942_ (_13989_, _13988_, _13986_);
  and _58943_ (_13990_, _13989_, _13982_);
  not _58944_ (_13991_, _13957_);
  nor _58945_ (_13992_, _13937_, _13935_);
  nor _58946_ (_13993_, _13992_, _13960_);
  nor _58947_ (_13994_, _13993_, _13991_);
  nor _58948_ (_13995_, _13957_, _13897_);
  nor _58949_ (_13996_, _13995_, _13994_);
  and _58950_ (_13997_, _13996_, _13886_);
  not _58951_ (_13998_, _13997_);
  nor _58952_ (_13999_, _13989_, _13982_);
  or _58953_ (_14000_, _13990_, _13999_);
  nor _58954_ (_14001_, _14000_, _13998_);
  or _58955_ (_14002_, _14001_, _13990_);
  and _58956_ (_14003_, _13933_, _13914_);
  not _58957_ (_14004_, _14003_);
  and _58958_ (_14005_, _14004_, _13934_);
  or _58959_ (_14006_, _14005_, _13991_);
  or _58960_ (_14007_, _13957_, _13911_);
  and _58961_ (_14008_, _14007_, _14006_);
  nor _58962_ (_14009_, _14008_, _13893_);
  not _58963_ (_14010_, _14009_);
  nand _58964_ (_14011_, _13991_, _13928_);
  nor _58965_ (_14012_, _13928_, _13923_);
  and _58966_ (_14013_, _13928_, _13923_);
  nor _58967_ (_14014_, _14013_, _14012_);
  nand _58968_ (_14015_, _13957_, _14014_);
  nand _58969_ (_14016_, _14015_, _14011_);
  nand _58970_ (_14017_, _14016_, _13916_);
  or _58971_ (_14018_, _14016_, _13916_);
  nand _58972_ (_14019_, _14018_, _14017_);
  nor _58973_ (_14020_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and _58974_ (_14021_, _13838_, _33848_);
  nor _58975_ (_14022_, _14021_, _14020_);
  nor _58976_ (_14023_, _14022_, _13924_);
  or _58977_ (_14024_, _14023_, _14019_);
  and _58978_ (_14025_, _14024_, _14017_);
  and _58979_ (_14026_, _13931_, _13929_);
  not _58980_ (_14027_, _14026_);
  and _58981_ (_14028_, _14027_, _13932_);
  or _58982_ (_14029_, _14028_, _13991_);
  or _58983_ (_14030_, _13957_, _13921_);
  and _58984_ (_14031_, _14030_, _14029_);
  nand _58985_ (_14032_, _14031_, _13907_);
  or _58986_ (_14033_, _14031_, _13907_);
  and _58987_ (_14034_, _14033_, _14032_);
  not _58988_ (_14035_, _14034_);
  or _58989_ (_14036_, _14035_, _14025_);
  and _58990_ (_14037_, _14008_, _13893_);
  not _58991_ (_14038_, _14037_);
  and _58992_ (_14039_, _14038_, _14032_);
  nand _58993_ (_14040_, _14039_, _14036_);
  and _58994_ (_14041_, _14040_, _14010_);
  nor _58995_ (_14042_, _13996_, _13886_);
  nor _58996_ (_14043_, _14042_, _13997_);
  not _58997_ (_14044_, _14000_);
  and _58998_ (_14045_, _14044_, _14043_);
  and _58999_ (_14046_, _14045_, _14041_);
  or _59000_ (_14047_, _14046_, _14002_);
  nand _59001_ (_14048_, _14047_, _13981_);
  or _59002_ (_14049_, _13970_, _13948_);
  and _59003_ (_14050_, _14049_, _13979_);
  nand _59004_ (_14051_, _14050_, _14048_);
  and _59005_ (_14052_, _13970_, _13948_);
  not _59006_ (_14053_, _14052_);
  and _59007_ (_14054_, _14053_, _13955_);
  and _59008_ (_14055_, _14054_, _14051_);
  or _59009_ (_14056_, _14055_, _13970_);
  nand _59010_ (_14057_, _14054_, _14051_);
  and _59011_ (_14058_, _14053_, _14049_);
  and _59012_ (_14059_, _14048_, _13979_);
  or _59013_ (_14060_, _14059_, _14058_);
  nand _59014_ (_14061_, _14059_, _14058_);
  and _59015_ (_14062_, _14061_, _14060_);
  or _59016_ (_14063_, _14062_, _14057_);
  and _59017_ (_14064_, _14063_, _14056_);
  or _59018_ (_14065_, _14064_, _13837_);
  nor _59019_ (_14066_, _34183_, _34180_);
  nor _59020_ (_14067_, _14066_, _35691_);
  and _59021_ (_14068_, _14067_, _33734_);
  nor _59022_ (_14069_, _14068_, _35693_);
  and _59023_ (_14070_, _14069_, _34180_);
  nor _59024_ (_14071_, _14069_, _34180_);
  nor _59025_ (_14072_, _14071_, _14070_);
  nor _59026_ (_14073_, _14072_, _35696_);
  and _59027_ (_14074_, _35712_, _33888_);
  not _59028_ (_14075_, _14074_);
  and _59029_ (_14076_, _33935_, _35707_);
  not _59030_ (_14077_, _14076_);
  and _59031_ (_14078_, _35681_, _35711_);
  nor _59032_ (_14079_, _14078_, _33929_);
  and _59033_ (_14080_, _14079_, _14077_);
  and _59034_ (_14081_, _14080_, _34212_);
  and _59035_ (_14082_, _14081_, _34209_);
  and _59036_ (_14083_, _14082_, _14075_);
  not _59037_ (_14084_, _14083_);
  nor _59038_ (_14085_, _14084_, _14073_);
  and _59039_ (_14086_, _14085_, _34203_);
  and _59040_ (_14087_, _35632_, _35639_);
  nor _59041_ (_14088_, _35632_, _35639_);
  nor _59042_ (_14089_, _14088_, _14087_);
  and _59043_ (_14090_, _14089_, _35582_);
  and _59044_ (_14091_, _35670_, _35639_);
  not _59045_ (_14092_, _14091_);
  nor _59046_ (_14093_, _35671_, _35638_);
  and _59047_ (_14094_, _14093_, _14092_);
  nor _59048_ (_14095_, _14094_, _14090_);
  and _59049_ (_14096_, _14095_, _14086_);
  and _59050_ (_14097_, _14096_, _13733_);
  and _59051_ (_14098_, _14097_, _14065_);
  nor _59052_ (_14099_, _14098_, _13836_);
  and _59053_ (_14100_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _33129_);
  and _59054_ (_14101_, _14100_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _59055_ (_14102_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _59056_ (_14103_, _14102_, _14101_);
  or _59057_ (_14104_, _14103_, _14099_);
  nor _59058_ (_14105_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not _59059_ (_14106_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _59060_ (_14107_, _14106_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _59061_ (_14108_, _14107_, _14105_);
  nor _59062_ (_14109_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not _59063_ (_14110_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _59064_ (_14111_, _14110_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _59065_ (_14112_, _14111_, _14109_);
  not _59066_ (_14113_, _14112_);
  nor _59067_ (_14114_, _14113_, _35672_);
  nor _59068_ (_14115_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not _59069_ (_14116_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _59070_ (_14117_, _14116_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _59071_ (_14118_, _14117_, _14115_);
  and _59072_ (_14119_, _14118_, _14114_);
  nor _59073_ (_14120_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not _59074_ (_14121_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _59075_ (_14122_, _14121_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _59076_ (_14123_, _14122_, _14120_);
  and _59077_ (_14124_, _14123_, _14119_);
  and _59078_ (_14125_, _14124_, _14108_);
  nor _59079_ (_14126_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not _59080_ (_14127_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _59081_ (_14128_, _14127_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _59082_ (_14129_, _14128_, _14126_);
  and _59083_ (_14130_, _14129_, _14125_);
  nor _59084_ (_14131_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not _59085_ (_14132_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _59086_ (_14133_, _14132_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _59087_ (_14134_, _14133_, _14131_);
  and _59088_ (_14135_, _14134_, _14130_);
  nor _59089_ (_14136_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not _59090_ (_14137_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _59091_ (_14138_, _14137_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _59092_ (_14139_, _14138_, _14136_);
  nand _59093_ (_14140_, _14139_, _14135_);
  nor _59094_ (_14141_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not _59095_ (_14142_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _59096_ (_14143_, _14142_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _59097_ (_14144_, _14143_, _14141_);
  and _59098_ (_14145_, _14144_, _14140_);
  nor _59099_ (_14146_, _14144_, _14140_);
  or _59100_ (_14147_, _14146_, _14145_);
  nand _59101_ (_14148_, _14147_, _35637_);
  and _59102_ (_14149_, _13713_, _13675_);
  not _59103_ (_14150_, _14149_);
  and _59104_ (_14151_, _14150_, _13714_);
  and _59105_ (_14152_, _14151_, _13534_);
  nor _59106_ (_14153_, _34132_, _34180_);
  and _59107_ (_14154_, _14153_, _34181_);
  and _59108_ (_14155_, _14154_, _34098_);
  and _59109_ (_14156_, _14155_, _34062_);
  and _59110_ (_14157_, _35623_, _33734_);
  and _59111_ (_14158_, _14157_, _14156_);
  nor _59112_ (_14159_, _35587_, _33734_);
  and _59113_ (_14160_, _34184_, _34180_);
  and _59114_ (_14161_, _13772_, _14160_);
  and _59115_ (_14162_, _14161_, _33987_);
  and _59116_ (_14163_, _14162_, _14159_);
  or _59117_ (_14164_, _14163_, _14158_);
  and _59118_ (_14165_, _33951_, _33734_);
  and _59119_ (_14166_, _33987_, _33734_);
  nor _59120_ (_14167_, _14166_, _14165_);
  and _59121_ (_14168_, _14167_, _14164_);
  and _59122_ (_14169_, _33778_, _33734_);
  nor _59123_ (_14170_, _14169_, _33779_);
  and _59124_ (_14171_, _14170_, _14168_);
  and _59125_ (_14172_, _14171_, _34197_);
  nor _59126_ (_14173_, _14171_, _34197_);
  nor _59127_ (_14174_, _14173_, _14172_);
  and _59128_ (_14175_, _14174_, _33899_);
  and _59129_ (_14176_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and _59130_ (_14177_, _34197_, _33734_);
  nor _59131_ (_14178_, _14177_, _35697_);
  nor _59132_ (_14179_, _14178_, _34006_);
  and _59133_ (_14180_, _35708_, _33815_);
  and _59134_ (_14181_, _33935_, _34197_);
  or _59135_ (_14182_, _14181_, _14180_);
  or _59136_ (_14183_, _14182_, _14179_);
  nor _59137_ (_14184_, _14183_, _14176_);
  not _59138_ (_14185_, _14184_);
  nor _59139_ (_14186_, _14185_, _14175_);
  not _59140_ (_14187_, _14186_);
  nor _59141_ (_14188_, _14187_, _14152_);
  and _59142_ (_14189_, _14188_, _14148_);
  nand _59143_ (_14190_, _14189_, _14101_);
  and _59144_ (_14191_, _14190_, _38997_);
  and _59145_ (_38993_[7], _14191_, _14104_);
  and _59146_ (_14192_, _11342_, _33665_);
  nor _59147_ (_14193_, _14192_, _14101_);
  not _59148_ (_14194_, _14193_);
  nand _59149_ (_14195_, _14194_, _14098_);
  or _59150_ (_14196_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _59151_ (_14197_, _14196_, _38997_);
  and _59152_ (_38994_[7], _14197_, _14195_);
  not _59153_ (_14198_, _14022_);
  and _59154_ (_14199_, _14055_, _13923_);
  nor _59155_ (_14200_, _14199_, _14198_);
  and _59156_ (_14201_, _14199_, _14198_);
  or _59157_ (_14202_, _14201_, _14200_);
  nand _59158_ (_14203_, _14202_, _13774_);
  and _59159_ (_14204_, _13743_, _13534_);
  and _59160_ (_14205_, _35648_, _33734_);
  nor _59161_ (_14206_, _14205_, _35649_);
  nand _59162_ (_14207_, _14206_, _35582_);
  nor _59163_ (_14208_, _35696_, _33848_);
  and _59164_ (_14209_, _35708_, _33888_);
  nor _59165_ (_14210_, _14209_, _14208_);
  nand _59166_ (_14211_, _14206_, _35637_);
  and _59167_ (_14212_, _35675_, _35707_);
  or _59168_ (_14213_, _34213_, _33831_);
  nand _59169_ (_14214_, _33935_, _35711_);
  nand _59170_ (_14215_, _14214_, _14213_);
  nor _59171_ (_14216_, _14215_, _14212_);
  and _59172_ (_14217_, _14216_, _34145_);
  and _59173_ (_14218_, _14217_, _14211_);
  and _59174_ (_14219_, _14218_, _14210_);
  and _59175_ (_14220_, _14219_, _14207_);
  not _59176_ (_14221_, _14220_);
  nor _59177_ (_14222_, _14221_, _14204_);
  nand _59178_ (_14223_, _14222_, _14203_);
  not _59179_ (_14224_, _14223_);
  nor _59180_ (_14225_, _14224_, _13836_);
  and _59181_ (_14226_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _59182_ (_14227_, _14226_, _14101_);
  or _59183_ (_14228_, _14227_, _14225_);
  not _59184_ (_14229_, _14101_);
  and _59185_ (_14230_, _34131_, _33935_);
  and _59186_ (_14231_, _35708_, _33884_);
  nor _59187_ (_14232_, _35697_, _34200_);
  not _59188_ (_14233_, _14232_);
  nor _59189_ (_14234_, _14233_, _34186_);
  nor _59190_ (_14235_, _14234_, _34131_);
  and _59191_ (_14236_, _14234_, _34131_);
  or _59192_ (_14237_, _14236_, _34100_);
  nor _59193_ (_14238_, _14237_, _14235_);
  nor _59194_ (_14239_, _34006_, _33848_);
  or _59195_ (_14240_, _14239_, _14238_);
  or _59196_ (_14241_, _14240_, _14231_);
  and _59197_ (_14242_, _14055_, _13774_);
  and _59198_ (_14243_, _14113_, _35672_);
  nor _59199_ (_14244_, _14243_, _14114_);
  and _59200_ (_14245_, _14244_, _35637_);
  and _59201_ (_14246_, _13621_, _13534_);
  or _59202_ (_14247_, _14246_, _14245_);
  or _59203_ (_14248_, _14247_, _14242_);
  or _59204_ (_14249_, _14248_, _14241_);
  or _59205_ (_14250_, _14249_, _14230_);
  or _59206_ (_14251_, _14250_, _14229_);
  and _59207_ (_14252_, _14251_, _38997_);
  and _59208_ (_38993_[0], _14252_, _14228_);
  nand _59209_ (_14253_, _13747_, _13534_);
  and _59210_ (_14254_, _14023_, _14019_);
  not _59211_ (_14255_, _14254_);
  and _59212_ (_14256_, _14255_, _14024_);
  or _59213_ (_14257_, _14256_, _14057_);
  or _59214_ (_14258_, _14055_, _14016_);
  and _59215_ (_14259_, _14258_, _14257_);
  nand _59216_ (_14260_, _14259_, _13774_);
  nor _59217_ (_14261_, _34134_, _34111_);
  or _59218_ (_14262_, _14261_, _35641_);
  and _59219_ (_14263_, _14262_, _35649_);
  nor _59220_ (_14264_, _14262_, _35649_);
  or _59221_ (_14265_, _14264_, _14263_);
  and _59222_ (_14266_, _14265_, _35637_);
  nor _59223_ (_14267_, _35619_, _35618_);
  nor _59224_ (_14268_, _14267_, _35620_);
  nor _59225_ (_14269_, _14268_, _35583_);
  nor _59226_ (_14270_, _14269_, _14266_);
  nor _59227_ (_14271_, _35690_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _59228_ (_14272_, _14271_, _13593_);
  nor _59229_ (_14273_, _14271_, _13593_);
  nor _59230_ (_14274_, _14273_, _14272_);
  nor _59231_ (_14275_, _14274_, _35696_);
  or _59232_ (_14276_, _33928_, _33848_);
  nand _59233_ (_14277_, _33934_, _33865_);
  not _59234_ (_14278_, _14277_);
  and _59235_ (_14279_, _33935_, _13593_);
  nor _59236_ (_14280_, _14279_, _14278_);
  and _59237_ (_14281_, _14280_, _14276_);
  and _59238_ (_14282_, _14281_, _34116_);
  and _59239_ (_14283_, _14282_, _34113_);
  not _59240_ (_14284_, _14283_);
  nor _59241_ (_14285_, _14284_, _14275_);
  and _59242_ (_14286_, _14285_, _34106_);
  and _59243_ (_14287_, _14286_, _14270_);
  and _59244_ (_14288_, _14287_, _14260_);
  nand _59245_ (_14289_, _14288_, _14253_);
  not _59246_ (_14290_, _14289_);
  nor _59247_ (_14291_, _14290_, _13836_);
  and _59248_ (_14292_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _59249_ (_14293_, _14292_, _14101_);
  or _59250_ (_14294_, _14293_, _14291_);
  nor _59251_ (_14295_, _14118_, _14114_);
  nor _59252_ (_14296_, _14295_, _14119_);
  and _59253_ (_14297_, _14296_, _35637_);
  not _59254_ (_14298_, _14297_);
  and _59255_ (_14299_, _13957_, _13774_);
  not _59256_ (_14300_, _14299_);
  and _59257_ (_14301_, _14154_, _33734_);
  and _59258_ (_14302_, _34132_, _14160_);
  and _59259_ (_14303_, _14302_, _33888_);
  nor _59260_ (_14304_, _14303_, _14301_);
  nor _59261_ (_14305_, _14304_, _34098_);
  and _59262_ (_14306_, _14304_, _34098_);
  nor _59263_ (_14307_, _14306_, _14305_);
  nor _59264_ (_14308_, _14307_, _34100_);
  and _59265_ (_14309_, _34098_, _33935_);
  and _59266_ (_14310_, _13562_, _35711_);
  not _59267_ (_14311_, _14310_);
  and _59268_ (_14312_, _14311_, _13597_);
  nor _59269_ (_14313_, _14312_, _13622_);
  and _59270_ (_14314_, _14313_, _13534_);
  and _59271_ (_14315_, _35708_, _33798_);
  nor _59272_ (_14316_, _34006_, _33831_);
  or _59273_ (_14317_, _14316_, _14315_);
  or _59274_ (_14318_, _14317_, _14314_);
  nor _59275_ (_14319_, _14318_, _14309_);
  not _59276_ (_14320_, _14319_);
  nor _59277_ (_14321_, _14320_, _14308_);
  and _59278_ (_14322_, _14321_, _14300_);
  and _59279_ (_14323_, _14322_, _14298_);
  nand _59280_ (_14324_, _14323_, _14101_);
  and _59281_ (_14325_, _14324_, _38997_);
  and _59282_ (_38993_[1], _14325_, _14294_);
  nand _59283_ (_14326_, _13752_, _13534_);
  not _59284_ (_14327_, _14036_);
  and _59285_ (_14328_, _14035_, _14025_);
  nor _59286_ (_14329_, _14328_, _14327_);
  or _59287_ (_14330_, _14329_, _14057_);
  or _59288_ (_14331_, _14055_, _14031_);
  and _59289_ (_14332_, _14331_, _14330_);
  nand _59290_ (_14333_, _14332_, _13774_);
  nor _59291_ (_14334_, _35620_, _35615_);
  nor _59292_ (_14335_, _14334_, _35621_);
  nor _59293_ (_14336_, _14335_, _35583_);
  or _59294_ (_14337_, _34213_, _33814_);
  and _59295_ (_14338_, _33935_, _33865_);
  nor _59296_ (_14339_, _34117_, _14338_);
  and _59297_ (_14340_, _14339_, _14337_);
  and _59298_ (_14341_, _14340_, _34082_);
  and _59299_ (_14342_, _14341_, _34079_);
  not _59300_ (_14343_, _14342_);
  nor _59301_ (_14344_, _14343_, _14336_);
  nor _59302_ (_14345_, _35652_, _35650_);
  nor _59303_ (_14346_, _14345_, _35638_);
  and _59304_ (_14347_, _14346_, _35654_);
  and _59305_ (_14348_, _35689_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _59306_ (_14349_, _14273_, _34064_);
  nor _59307_ (_14350_, _14349_, _14348_);
  nor _59308_ (_14351_, _14350_, _35696_);
  nor _59309_ (_14352_, _14351_, _14347_);
  and _59310_ (_14353_, _14352_, _14344_);
  and _59311_ (_14354_, _14353_, _34073_);
  and _59312_ (_14355_, _14354_, _14333_);
  and _59313_ (_14356_, _14355_, _14326_);
  nor _59314_ (_14357_, _14356_, _13836_);
  and _59315_ (_14358_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _59316_ (_14359_, _14358_, _14101_);
  or _59317_ (_14360_, _14359_, _14357_);
  nor _59318_ (_14361_, _14123_, _14119_);
  nor _59319_ (_14362_, _14361_, _14124_);
  and _59320_ (_14363_, _14362_, _35637_);
  not _59321_ (_14364_, _14363_);
  and _59322_ (_14365_, _14302_, _34107_);
  and _59323_ (_14366_, _14365_, _33888_);
  and _59324_ (_14367_, _14155_, _33734_);
  nor _59325_ (_14368_, _14367_, _14366_);
  and _59326_ (_14369_, _14368_, _35601_);
  nor _59327_ (_14370_, _14368_, _35601_);
  or _59328_ (_14371_, _14370_, _34100_);
  nor _59329_ (_14372_, _14371_, _14369_);
  nor _59330_ (_14373_, _13699_, _13696_);
  nor _59331_ (_14374_, _14373_, _13700_);
  and _59332_ (_14375_, _14374_, _13534_);
  and _59333_ (_14376_, _34062_, _33935_);
  and _59334_ (_14377_, _35708_, _33766_);
  and _59335_ (_14378_, _33674_, _33865_);
  and _59336_ (_14379_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or _59337_ (_14380_, _14379_, _14378_);
  or _59338_ (_14381_, _14380_, _14377_);
  nor _59339_ (_14382_, _14381_, _14376_);
  not _59340_ (_14383_, _14382_);
  nor _59341_ (_14384_, _14383_, _14375_);
  not _59342_ (_14385_, _14384_);
  nor _59343_ (_14386_, _14385_, _14372_);
  and _59344_ (_14387_, _14386_, _14364_);
  nand _59345_ (_14388_, _14387_, _14101_);
  and _59346_ (_14389_, _14388_, _38997_);
  and _59347_ (_38993_[2], _14389_, _14360_);
  not _59348_ (_14390_, _14008_);
  or _59349_ (_14391_, _14055_, _14390_);
  or _59350_ (_14392_, _14037_, _14009_);
  and _59351_ (_14393_, _14036_, _14032_);
  and _59352_ (_14394_, _14393_, _14392_);
  nor _59353_ (_14395_, _14393_, _14392_);
  or _59354_ (_14396_, _14395_, _14394_);
  or _59355_ (_14397_, _14396_, _14057_);
  nand _59356_ (_14398_, _14397_, _14391_);
  nand _59357_ (_14399_, _14398_, _13774_);
  nor _59358_ (_14400_, _35621_, _35612_);
  nor _59359_ (_14401_, _14400_, _35622_);
  nor _59360_ (_14402_, _14401_, _35583_);
  not _59361_ (_14403_, _14402_);
  and _59362_ (_14404_, _35654_, _35647_);
  or _59363_ (_14405_, _14404_, _35638_);
  nor _59364_ (_14406_, _14405_, _35655_);
  not _59365_ (_14407_, _14406_);
  nor _59366_ (_14408_, _35689_, _13828_);
  nor _59367_ (_14409_, _14408_, _33815_);
  and _59368_ (_14410_, _33935_, _33815_);
  nor _59369_ (_14411_, _35690_, _35696_);
  nor _59370_ (_14412_, _14411_, _14410_);
  nor _59371_ (_14413_, _14412_, _14409_);
  or _59372_ (_14414_, _34213_, _33883_);
  not _59373_ (_14415_, _34083_);
  and _59374_ (_14416_, _14415_, _14414_);
  not _59375_ (_14417_, _14416_);
  nor _59376_ (_14418_, _14417_, _14413_);
  and _59377_ (_14419_, _14418_, _34051_);
  and _59378_ (_14420_, _14419_, _14407_);
  and _59379_ (_14421_, _14420_, _14403_);
  and _59380_ (_14422_, _14421_, _14399_);
  and _59381_ (_14423_, _14422_, _13785_);
  nor _59382_ (_14424_, _14423_, _13836_);
  and _59383_ (_14425_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _59384_ (_14426_, _14425_, _14101_);
  or _59385_ (_14427_, _14426_, _14424_);
  nor _59386_ (_14428_, _14124_, _14108_);
  not _59387_ (_14429_, _14428_);
  nor _59388_ (_14430_, _14125_, _35638_);
  and _59389_ (_14431_, _14430_, _14429_);
  not _59390_ (_14432_, _14431_);
  and _59391_ (_14433_, _13703_, _13701_);
  not _59392_ (_14434_, _14433_);
  and _59393_ (_14435_, _14434_, _13704_);
  and _59394_ (_14436_, _14435_, _13534_);
  not _59395_ (_14437_, _14436_);
  and _59396_ (_14438_, _14156_, _33734_);
  and _59397_ (_14439_, _14365_, _35601_);
  and _59398_ (_14440_, _14439_, _33888_);
  nor _59399_ (_14441_, _14440_, _14438_);
  nor _59400_ (_14442_, _14441_, _34035_);
  not _59401_ (_14443_, _14442_);
  and _59402_ (_14444_, _14441_, _34035_);
  nor _59403_ (_14445_, _14444_, _34100_);
  and _59404_ (_14446_, _14445_, _14443_);
  and _59405_ (_14447_, _35623_, _33935_);
  nor _59406_ (_14448_, _34006_, _33814_);
  and _59407_ (_14449_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or _59408_ (_14450_, _14449_, _14448_);
  or _59409_ (_14451_, _14450_, _35709_);
  nor _59410_ (_14452_, _14451_, _14447_);
  not _59411_ (_14453_, _14452_);
  nor _59412_ (_14454_, _14453_, _14446_);
  and _59413_ (_14455_, _14454_, _14437_);
  and _59414_ (_14456_, _14455_, _14432_);
  nand _59415_ (_14457_, _14456_, _14101_);
  and _59416_ (_14458_, _14457_, _38997_);
  and _59417_ (_38993_[3], _14458_, _14427_);
  nand _59418_ (_14459_, _14043_, _14041_);
  or _59419_ (_14460_, _14043_, _14041_);
  and _59420_ (_14461_, _14460_, _14459_);
  and _59421_ (_14462_, _14461_, _14055_);
  and _59422_ (_14463_, _14057_, _13996_);
  or _59423_ (_14464_, _14463_, _14462_);
  nand _59424_ (_14465_, _14464_, _13774_);
  nand _59425_ (_14466_, _13755_, _13534_);
  nor _59426_ (_14467_, _35628_, _33991_);
  and _59427_ (_14468_, _35628_, _33991_);
  nor _59428_ (_14469_, _14468_, _14467_);
  and _59429_ (_14470_, _14469_, _35582_);
  not _59430_ (_14471_, _14470_);
  not _59431_ (_14472_, _35659_);
  nor _59432_ (_14473_, _35658_, _33991_);
  nor _59433_ (_14474_, _14473_, _35638_);
  and _59434_ (_14475_, _14474_, _14472_);
  nor _59435_ (_14476_, _35691_, _33884_);
  not _59436_ (_14477_, _14476_);
  nor _59437_ (_14478_, _35692_, _35696_);
  and _59438_ (_14479_, _14478_, _14477_);
  and _59439_ (_14480_, _33935_, _33884_);
  not _59440_ (_14481_, _14480_);
  or _59441_ (_14482_, _34213_, _33797_);
  not _59442_ (_14483_, _34020_);
  and _59443_ (_14484_, _14483_, _14482_);
  and _59444_ (_14485_, _14484_, _14481_);
  and _59445_ (_14486_, _14485_, _33993_);
  not _59446_ (_14487_, _14486_);
  nor _59447_ (_14488_, _14487_, _14479_);
  and _59448_ (_14489_, _14488_, _34016_);
  not _59449_ (_14490_, _14489_);
  nor _59450_ (_14491_, _14490_, _14475_);
  and _59451_ (_14492_, _14491_, _14471_);
  and _59452_ (_14493_, _14492_, _14466_);
  nand _59453_ (_14494_, _14493_, _14465_);
  not _59454_ (_14495_, _14494_);
  nor _59455_ (_14496_, _14495_, _13836_);
  and _59456_ (_14497_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _59457_ (_14498_, _14497_, _14101_);
  or _59458_ (_14499_, _14498_, _14496_);
  nor _59459_ (_14500_, _14129_, _14125_);
  nor _59460_ (_14501_, _14500_, _14130_);
  and _59461_ (_14502_, _14501_, _35637_);
  not _59462_ (_14503_, _14502_);
  and _59463_ (_14504_, _13707_, _13705_);
  not _59464_ (_14505_, _14504_);
  and _59465_ (_14506_, _14505_, _13708_);
  and _59466_ (_14507_, _14506_, _13534_);
  and _59467_ (_14508_, _14161_, _33888_);
  nor _59468_ (_14509_, _14508_, _14158_);
  and _59469_ (_14510_, _14509_, _33987_);
  nor _59470_ (_14511_, _14509_, _33987_);
  nor _59471_ (_14512_, _14511_, _14510_);
  and _59472_ (_14513_, _14512_, _33899_);
  nor _59473_ (_14514_, _33884_, _33734_);
  not _59474_ (_14515_, _14514_);
  nor _59475_ (_14516_, _14166_, _34006_);
  and _59476_ (_14517_, _14516_, _14515_);
  and _59477_ (_14518_, _34007_, _33935_);
  and _59478_ (_14519_, _35708_, _35711_);
  and _59479_ (_14520_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or _59480_ (_14521_, _14520_, _14519_);
  nor _59481_ (_14522_, _14521_, _14518_);
  not _59482_ (_14523_, _14522_);
  nor _59483_ (_14524_, _14523_, _14517_);
  not _59484_ (_14525_, _14524_);
  nor _59485_ (_14526_, _14525_, _14513_);
  not _59486_ (_14527_, _14526_);
  nor _59487_ (_14528_, _14527_, _14507_);
  and _59488_ (_14529_, _14528_, _14503_);
  nand _59489_ (_14530_, _14529_, _14101_);
  and _59490_ (_14531_, _14530_, _38997_);
  and _59491_ (_38993_[4], _14531_, _14499_);
  nand _59492_ (_14532_, _14057_, _13989_);
  and _59493_ (_14533_, _14459_, _13998_);
  nand _59494_ (_14534_, _14533_, _14044_);
  or _59495_ (_14535_, _14533_, _14044_);
  nand _59496_ (_14536_, _14535_, _14534_);
  nand _59497_ (_14537_, _14536_, _14055_);
  nand _59498_ (_14538_, _14537_, _14532_);
  nand _59499_ (_14539_, _14538_, _13774_);
  nand _59500_ (_14540_, _13738_, _13534_);
  nor _59501_ (_14541_, _35629_, _35599_);
  nor _59502_ (_14542_, _14541_, _35630_);
  nor _59503_ (_14543_, _14542_, _35583_);
  not _59504_ (_14544_, _14543_);
  nor _59505_ (_14545_, _33990_, _33967_);
  or _59506_ (_14546_, _14545_, _35662_);
  and _59507_ (_14547_, _14546_, _14472_);
  or _59508_ (_14548_, _14547_, _35638_);
  nor _59509_ (_14549_, _14548_, _35660_);
  nor _59510_ (_14550_, _14068_, _35692_);
  and _59511_ (_14551_, _14550_, _33797_);
  nor _59512_ (_14552_, _14550_, _33797_);
  nor _59513_ (_14553_, _14552_, _14551_);
  nor _59514_ (_14554_, _14553_, _35696_);
  and _59515_ (_14555_, _33935_, _33798_);
  not _59516_ (_14556_, _14555_);
  or _59517_ (_14557_, _34213_, _33765_);
  not _59518_ (_14558_, _33994_);
  and _59519_ (_14559_, _14558_, _14557_);
  and _59520_ (_14560_, _14559_, _14556_);
  and _59521_ (_14561_, _14560_, _33972_);
  and _59522_ (_14562_, _14561_, _33969_);
  not _59523_ (_14563_, _14562_);
  nor _59524_ (_14564_, _14563_, _14554_);
  and _59525_ (_14565_, _14564_, _33963_);
  not _59526_ (_14566_, _14565_);
  nor _59527_ (_14567_, _14566_, _14549_);
  and _59528_ (_14568_, _14567_, _14544_);
  and _59529_ (_14569_, _14568_, _14540_);
  and _59530_ (_14570_, _14569_, _14539_);
  nor _59531_ (_14571_, _14570_, _13836_);
  and _59532_ (_14572_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _59533_ (_14573_, _14572_, _14101_);
  or _59534_ (_14574_, _14573_, _14571_);
  nor _59535_ (_14575_, _14134_, _14130_);
  nor _59536_ (_14576_, _14575_, _14135_);
  and _59537_ (_14577_, _14576_, _35637_);
  not _59538_ (_14578_, _14577_);
  and _59539_ (_14579_, _13709_, _13687_);
  not _59540_ (_14580_, _14579_);
  and _59541_ (_14581_, _14580_, _13710_);
  and _59542_ (_14582_, _14581_, _13534_);
  nor _59543_ (_14583_, _14162_, _14158_);
  nor _59544_ (_14584_, _14583_, _14166_);
  and _59545_ (_14585_, _14584_, _33951_);
  nor _59546_ (_14586_, _14584_, _33951_);
  or _59547_ (_14587_, _14586_, _14585_);
  and _59548_ (_14588_, _14587_, _33899_);
  and _59549_ (_14589_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor _59550_ (_14590_, _33798_, _33734_);
  or _59551_ (_14591_, _14590_, _34006_);
  nor _59552_ (_14592_, _14591_, _14165_);
  and _59553_ (_14593_, _35708_, _13593_);
  and _59554_ (_14594_, _35587_, _33935_);
  or _59555_ (_14595_, _14594_, _14593_);
  or _59556_ (_14596_, _14595_, _14592_);
  nor _59557_ (_14597_, _14596_, _14589_);
  not _59558_ (_14598_, _14597_);
  nor _59559_ (_14599_, _14598_, _14588_);
  not _59560_ (_14600_, _14599_);
  nor _59561_ (_14601_, _14600_, _14582_);
  and _59562_ (_14602_, _14601_, _14578_);
  nand _59563_ (_14603_, _14602_, _14101_);
  and _59564_ (_14604_, _14603_, _38997_);
  and _59565_ (_38993_[5], _14604_, _14574_);
  or _59566_ (_14605_, _14047_, _13981_);
  and _59567_ (_14606_, _14605_, _14048_);
  or _59568_ (_14607_, _14606_, _14057_);
  or _59569_ (_14608_, _14055_, _13978_);
  and _59570_ (_14609_, _14608_, _14607_);
  and _59571_ (_14610_, _14609_, _13774_);
  and _59572_ (_14611_, _13735_, _13534_);
  or _59573_ (_14612_, _35666_, _35660_);
  nor _59574_ (_14613_, _35667_, _35638_);
  and _59575_ (_14614_, _14613_, _14612_);
  nor _59576_ (_14615_, _35630_, _35596_);
  nor _59577_ (_14616_, _14615_, _35631_);
  nor _59578_ (_14617_, _14616_, _35583_);
  nor _59579_ (_14618_, _14551_, _33765_);
  and _59580_ (_14619_, _14551_, _33765_);
  or _59581_ (_14620_, _14619_, _14618_);
  and _59582_ (_14621_, _14620_, _35688_);
  and _59583_ (_14622_, _33935_, _33766_);
  or _59584_ (_14623_, _33973_, _34214_);
  nor _59585_ (_14624_, _14623_, _14622_);
  and _59586_ (_14625_, _14624_, _33926_);
  nand _59587_ (_14626_, _14625_, _33918_);
  nor _59588_ (_14627_, _14626_, _14621_);
  nand _59589_ (_14628_, _14627_, _33903_);
  or _59590_ (_14629_, _14628_, _14617_);
  or _59591_ (_14630_, _14629_, _14614_);
  or _59592_ (_14631_, _14630_, _14611_);
  or _59593_ (_14632_, _14631_, _14610_);
  or _59594_ (_14633_, _14632_, _13836_);
  not _59595_ (_14634_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nand _59596_ (_14635_, _13836_, _14634_);
  and _59597_ (_14636_, _14635_, _14633_);
  or _59598_ (_14637_, _14636_, _14101_);
  or _59599_ (_14638_, _14139_, _14135_);
  and _59600_ (_14639_, _14638_, _14140_);
  and _59601_ (_14640_, _14639_, _35637_);
  or _59602_ (_14641_, _13711_, _13681_);
  and _59603_ (_14642_, _14641_, _13712_);
  and _59604_ (_14643_, _14642_, _13534_);
  and _59605_ (_14644_, _14168_, _33778_);
  nor _59606_ (_14645_, _14168_, _33778_);
  or _59607_ (_14646_, _14645_, _14644_);
  and _59608_ (_14647_, _14646_, _33899_);
  or _59609_ (_14648_, _33766_, _33734_);
  nor _59610_ (_14649_, _14169_, _34006_);
  and _59611_ (_14650_, _14649_, _14648_);
  and _59612_ (_14651_, _35708_, _33865_);
  and _59613_ (_14652_, _35585_, _33935_);
  and _59614_ (_14653_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  or _59615_ (_14654_, _14653_, _14652_);
  or _59616_ (_14655_, _14654_, _14651_);
  or _59617_ (_14656_, _14655_, _14650_);
  or _59618_ (_14657_, _14656_, _14647_);
  or _59619_ (_14658_, _14657_, _14643_);
  or _59620_ (_14659_, _14658_, _14640_);
  or _59621_ (_14660_, _14659_, _14229_);
  and _59622_ (_14661_, _14660_, _38997_);
  and _59623_ (_38993_[6], _14661_, _14637_);
  or _59624_ (_14662_, _14223_, _14193_);
  or _59625_ (_14663_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _59626_ (_14664_, _14663_, _38997_);
  and _59627_ (_38994_[0], _14664_, _14662_);
  or _59628_ (_14665_, _14289_, _14193_);
  or _59629_ (_14666_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _59630_ (_14667_, _14666_, _38997_);
  and _59631_ (_38994_[1], _14667_, _14665_);
  nand _59632_ (_14668_, _14356_, _14194_);
  or _59633_ (_14669_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _59634_ (_14670_, _14669_, _38997_);
  and _59635_ (_38994_[2], _14670_, _14668_);
  nand _59636_ (_14671_, _14423_, _14194_);
  or _59637_ (_14672_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _59638_ (_14673_, _14672_, _38997_);
  and _59639_ (_38994_[3], _14673_, _14671_);
  or _59640_ (_14674_, _14494_, _14193_);
  or _59641_ (_14675_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _59642_ (_14676_, _14675_, _38997_);
  and _59643_ (_38994_[4], _14676_, _14674_);
  nand _59644_ (_14677_, _14570_, _14194_);
  or _59645_ (_14678_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _59646_ (_14679_, _14678_, _38997_);
  and _59647_ (_38994_[5], _14679_, _14677_);
  or _59648_ (_14680_, _14632_, _14193_);
  or _59649_ (_14681_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _59650_ (_14682_, _14681_, _38997_);
  and _59651_ (_38994_[6], _14682_, _14680_);
  and _59652_ (_36923_, _33533_, _38997_);
  and _59653_ (_39017_, _36923_, _33475_);
  and _59654_ (_39018_[7], _34223_, _38997_);
  nand _59655_ (_39018_[0], _34466_, _38997_);
  nand _59656_ (_39018_[1], _34557_, _38997_);
  nand _59657_ (_39018_[2], _34766_, _38997_);
  and _59658_ (_39018_[3], _34401_, _38997_);
  and _59659_ (_39018_[4], _34525_, _38997_);
  nor _59660_ (_39018_[5], _34615_, rst);
  nor _59661_ (_39018_[6], _34649_, rst);
  not _59662_ (_14683_, _14098_);
  nand _59663_ (_14684_, _13158_, _34231_);
  or _59664_ (_14685_, _14684_, _14683_);
  not _59665_ (_14686_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _59666_ (_14687_, _14684_, _14686_);
  and _59667_ (_14688_, _14687_, _33662_);
  and _59668_ (_14689_, _14688_, _14685_);
  nor _59669_ (_14690_, _33661_, _14686_);
  nor _59670_ (_14691_, _33630_, _33591_);
  and _59671_ (_14692_, _14691_, _13123_);
  and _59672_ (_14693_, _14692_, _11075_);
  nand _59673_ (_14694_, _14693_, _35722_);
  or _59674_ (_14695_, _14693_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _59675_ (_14696_, _14695_, _11083_);
  and _59676_ (_14697_, _14696_, _14694_);
  or _59677_ (_14698_, _14697_, _14690_);
  or _59678_ (_14699_, _14698_, _14689_);
  and _59679_ (_38992_[7], _14699_, _38997_);
  or _59680_ (_14700_, _14684_, _14223_);
  not _59681_ (_14701_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _59682_ (_14702_, _14684_, _14701_);
  and _59683_ (_14703_, _14702_, _33662_);
  and _59684_ (_14704_, _14703_, _14700_);
  nor _59685_ (_14705_, _33661_, _14701_);
  or _59686_ (_14706_, _14684_, _35723_);
  and _59687_ (_14707_, _14702_, _11083_);
  and _59688_ (_14708_, _14707_, _14706_);
  or _59689_ (_14709_, _14708_, _14705_);
  or _59690_ (_14710_, _14709_, _14704_);
  and _59691_ (_38992_[0], _14710_, _38997_);
  or _59692_ (_14711_, _14684_, _14289_);
  not _59693_ (_14712_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _59694_ (_14713_, _14684_, _14712_);
  and _59695_ (_14714_, _14713_, _33662_);
  and _59696_ (_14715_, _14714_, _14711_);
  nor _59697_ (_14716_, _33661_, _14712_);
  and _59698_ (_14717_, _14692_, _34253_);
  nand _59699_ (_14718_, _14717_, _35722_);
  or _59700_ (_14719_, _14717_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _59701_ (_14720_, _14719_, _11083_);
  and _59702_ (_14721_, _14720_, _14718_);
  or _59703_ (_14722_, _14721_, _14716_);
  or _59704_ (_14723_, _14722_, _14715_);
  and _59705_ (_38992_[1], _14723_, _38997_);
  not _59706_ (_14724_, _14356_);
  or _59707_ (_14725_, _14684_, _14724_);
  not _59708_ (_14726_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _59709_ (_14727_, _14684_, _14726_);
  and _59710_ (_14728_, _14727_, _33662_);
  and _59711_ (_14729_, _14728_, _14725_);
  nor _59712_ (_14730_, _33661_, _14726_);
  nand _59713_ (_14731_, _14692_, _11359_);
  and _59714_ (_14732_, _14731_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _59715_ (_14733_, _34252_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _59716_ (_14734_, _14733_, _11345_);
  and _59717_ (_14735_, _14734_, _14692_);
  or _59718_ (_14736_, _14735_, _14732_);
  and _59719_ (_14737_, _14736_, _11083_);
  or _59720_ (_14738_, _14737_, _14730_);
  or _59721_ (_14739_, _14738_, _14729_);
  and _59722_ (_38992_[2], _14739_, _38997_);
  not _59723_ (_14740_, _14423_);
  or _59724_ (_14741_, _14684_, _14740_);
  not _59725_ (_14742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _59726_ (_14743_, _14684_, _14742_);
  and _59727_ (_14744_, _14743_, _33662_);
  and _59728_ (_14745_, _14744_, _14741_);
  nor _59729_ (_14746_, _33661_, _14742_);
  and _59730_ (_14747_, _14692_, _11356_);
  nand _59731_ (_14748_, _14747_, _35722_);
  or _59732_ (_14749_, _14747_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _59733_ (_14750_, _14749_, _11083_);
  and _59734_ (_14751_, _14750_, _14748_);
  or _59735_ (_14752_, _14751_, _14746_);
  or _59736_ (_14753_, _14752_, _14745_);
  and _59737_ (_38992_[3], _14753_, _38997_);
  or _59738_ (_14754_, _14684_, _14494_);
  not _59739_ (_14755_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _59740_ (_14756_, _14684_, _14755_);
  and _59741_ (_14757_, _14756_, _33662_);
  and _59742_ (_14758_, _14757_, _14754_);
  nor _59743_ (_14759_, _33661_, _14755_);
  and _59744_ (_14760_, _14692_, _11370_);
  nand _59745_ (_14761_, _14760_, _35722_);
  or _59746_ (_14762_, _14760_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _59747_ (_14763_, _14762_, _11083_);
  and _59748_ (_14764_, _14763_, _14761_);
  or _59749_ (_14765_, _14764_, _14759_);
  or _59750_ (_14766_, _14765_, _14758_);
  and _59751_ (_38992_[4], _14766_, _38997_);
  not _59752_ (_14767_, _14570_);
  or _59753_ (_14768_, _14684_, _14767_);
  not _59754_ (_14769_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _59755_ (_14770_, _14684_, _14769_);
  and _59756_ (_14771_, _14770_, _33662_);
  and _59757_ (_14772_, _14771_, _14768_);
  nor _59758_ (_14773_, _33661_, _14769_);
  and _59759_ (_14774_, _14692_, _11383_);
  nand _59760_ (_14775_, _14774_, _35722_);
  or _59761_ (_14776_, _14774_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _59762_ (_14777_, _14776_, _11083_);
  and _59763_ (_14778_, _14777_, _14775_);
  or _59764_ (_14779_, _14778_, _14773_);
  or _59765_ (_14780_, _14779_, _14772_);
  and _59766_ (_38992_[5], _14780_, _38997_);
  or _59767_ (_14781_, _14684_, _14632_);
  not _59768_ (_14782_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _59769_ (_14783_, _14684_, _14782_);
  and _59770_ (_14784_, _14783_, _33662_);
  and _59771_ (_14785_, _14784_, _14781_);
  nor _59772_ (_14786_, _33661_, _14782_);
  nand _59773_ (_14787_, _14692_, _11392_);
  or _59774_ (_14788_, _14787_, _35723_);
  nand _59775_ (_14789_, _14787_, _14782_);
  and _59776_ (_14790_, _14789_, _11083_);
  and _59777_ (_14791_, _14790_, _14788_);
  or _59778_ (_14792_, _14791_, _14786_);
  or _59779_ (_14793_, _14792_, _14785_);
  and _59780_ (_38992_[6], _14793_, _38997_);
  nor _59781_ (_14794_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _59782_ (_14795_, _14794_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _59783_ (_14796_, _12066_, _34231_);
  and _59784_ (_14797_, _14796_, _34257_);
  and _59785_ (_14798_, _14797_, _33662_);
  nor _59786_ (_14799_, _14798_, _14795_);
  or _59787_ (_14800_, _14799_, _14098_);
  not _59788_ (_14801_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _59789_ (_14802_, _14100_, _14801_);
  not _59790_ (_14803_, _14802_);
  and _59791_ (_14804_, _14691_, _11083_);
  and _59792_ (_14805_, _14804_, _13106_);
  and _59793_ (_14806_, _14805_, _11075_);
  and _59794_ (_14807_, _14806_, _35722_);
  nor _59795_ (_14808_, _14806_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _59796_ (_14809_, _14808_);
  nand _59797_ (_14810_, _14809_, _14799_);
  or _59798_ (_14811_, _14810_, _14807_);
  and _59799_ (_14812_, _14811_, _14803_);
  and _59800_ (_14813_, _14812_, _14800_);
  and _59801_ (_14814_, _14802_, _14189_);
  or _59802_ (_14815_, _14814_, _14813_);
  nor _59803_ (_38991_[7], _14815_, rst);
  or _59804_ (_14816_, _14799_, _14223_);
  nor _59805_ (_14817_, _34229_, _34128_);
  nor _59806_ (_14818_, _14817_, _11315_);
  or _59807_ (_14819_, _14802_, _14795_);
  nor _59808_ (_14820_, _14819_, _14798_);
  and _59809_ (_14821_, _14820_, _14805_);
  not _59810_ (_14822_, _14821_);
  nor _59811_ (_14823_, _14822_, _14818_);
  not _59812_ (_14824_, _14799_);
  nor _59813_ (_14825_, _14805_, _34128_);
  nor _59814_ (_14826_, _14825_, _14824_);
  not _59815_ (_14827_, _14826_);
  nor _59816_ (_14828_, _14827_, _14823_);
  nor _59817_ (_14829_, _14828_, _14802_);
  nand _59818_ (_14830_, _14829_, _14816_);
  nand _59819_ (_14831_, _14802_, _14250_);
  nand _59820_ (_14832_, _14831_, _14830_);
  and _59821_ (_38991_[0], _14832_, _38997_);
  nor _59822_ (_14833_, _14803_, _14323_);
  not _59823_ (_14834_, _14833_);
  or _59824_ (_14835_, _14799_, _14289_);
  not _59825_ (_14836_, _14805_);
  nor _59826_ (_14837_, _34253_, _34095_);
  nor _59827_ (_14838_, _14837_, _11326_);
  nor _59828_ (_14839_, _14838_, _14836_);
  nor _59829_ (_14840_, _14805_, _34095_);
  nor _59830_ (_14841_, _14840_, _14824_);
  not _59831_ (_14842_, _14841_);
  nor _59832_ (_14843_, _14842_, _14839_);
  nor _59833_ (_14844_, _14843_, _14802_);
  nand _59834_ (_14845_, _14844_, _14835_);
  nand _59835_ (_14846_, _14845_, _14834_);
  and _59836_ (_38991_[1], _14846_, _38997_);
  or _59837_ (_14847_, _14799_, _14356_);
  and _59838_ (_14848_, _14805_, _11343_);
  and _59839_ (_14849_, _14848_, _35722_);
  nor _59840_ (_14850_, _14848_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not _59841_ (_14851_, _14850_);
  nand _59842_ (_14852_, _14851_, _14799_);
  or _59843_ (_14853_, _14852_, _14849_);
  and _59844_ (_14854_, _14853_, _14803_);
  nand _59845_ (_14855_, _14854_, _14847_);
  and _59846_ (_14856_, _14802_, _14387_);
  not _59847_ (_14857_, _14856_);
  and _59848_ (_14858_, _14857_, _14855_);
  and _59849_ (_38991_[2], _14858_, _38997_);
  or _59850_ (_14859_, _14799_, _14423_);
  and _59851_ (_14860_, _14821_, _11357_);
  and _59852_ (_14861_, _14805_, _11356_);
  nand _59853_ (_14862_, _14799_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _59854_ (_14863_, _14862_, _14861_);
  or _59855_ (_14864_, _14863_, _14802_);
  nor _59856_ (_14865_, _14864_, _14860_);
  nand _59857_ (_14866_, _14865_, _14859_);
  and _59858_ (_14867_, _14802_, _14456_);
  not _59859_ (_14868_, _14867_);
  and _59860_ (_14869_, _14868_, _14866_);
  and _59861_ (_38991_[3], _14869_, _38997_);
  nor _59862_ (_14870_, _14803_, _14529_);
  not _59863_ (_14871_, _14870_);
  or _59864_ (_14872_, _14799_, _14494_);
  nor _59865_ (_14873_, _11370_, _33984_);
  nor _59866_ (_14874_, _14873_, _11376_);
  nor _59867_ (_14875_, _14874_, _14822_);
  nor _59868_ (_14876_, _14805_, _33984_);
  nor _59869_ (_14877_, _14876_, _14824_);
  not _59870_ (_14878_, _14877_);
  nor _59871_ (_14879_, _14878_, _14875_);
  nor _59872_ (_14880_, _14879_, _14802_);
  nand _59873_ (_14881_, _14880_, _14872_);
  nand _59874_ (_14882_, _14881_, _14871_);
  and _59875_ (_38991_[4], _14882_, _38997_);
  or _59876_ (_14883_, _14799_, _14570_);
  nand _59877_ (_14884_, _14821_, _11383_);
  or _59878_ (_14885_, _14884_, _35722_);
  and _59879_ (_14886_, _14805_, _11383_);
  nand _59880_ (_14887_, _14799_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _59881_ (_14888_, _14887_, _14886_);
  and _59882_ (_14889_, _14888_, _14803_);
  and _59883_ (_14890_, _14889_, _14885_);
  nand _59884_ (_14891_, _14890_, _14883_);
  and _59885_ (_14892_, _14802_, _14602_);
  not _59886_ (_14893_, _14892_);
  and _59887_ (_14894_, _14893_, _14891_);
  and _59888_ (_38991_[5], _14894_, _38997_);
  and _59889_ (_14895_, _14824_, _14632_);
  and _59890_ (_14896_, _14821_, _12080_);
  nand _59891_ (_14897_, _14805_, _11392_);
  and _59892_ (_14898_, _14799_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _59893_ (_14899_, _14898_, _14897_);
  or _59894_ (_14900_, _14899_, _14802_);
  or _59895_ (_14901_, _14900_, _14896_);
  or _59896_ (_14902_, _14901_, _14895_);
  or _59897_ (_14903_, _14803_, _14659_);
  and _59898_ (_14904_, _14903_, _14902_);
  and _59899_ (_38991_[6], _14904_, _38997_);
  and _59900_ (_14905_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _59901_ (_14906_, _14905_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _59902_ (_14907_, _14905_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _59903_ (_14908_, _14907_, _14906_);
  and _59904_ (_36859_[1], _14908_, _38997_);
  and _59905_ (_36860_[5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _38997_);
  nor _59906_ (_36861_[7], _14064_, rst);
  and _59907_ (_36860_[0], _14055_, _38997_);
  and _59908_ (_36860_[1], _13957_, _38997_);
  and _59909_ (_36860_[2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _38997_);
  and _59910_ (_36860_[3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _38997_);
  and _59911_ (_36860_[4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _38997_);
  or _59912_ (_14909_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _59913_ (_14910_, _14905_, rst);
  and _59914_ (_36859_[0], _14910_, _14909_);
  and _59915_ (_36861_[0], _14202_, _38997_);
  and _59916_ (_36861_[1], _14259_, _38997_);
  and _59917_ (_36861_[2], _14332_, _38997_);
  and _59918_ (_36861_[3], _14398_, _38997_);
  and _59919_ (_36861_[4], _14464_, _38997_);
  and _59920_ (_36861_[5], _14538_, _38997_);
  and _59921_ (_36861_[6], _14609_, _38997_);
  nand _59922_ (_14911_, _13548_, _13534_);
  or _59923_ (_14912_, _13534_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _59924_ (_14913_, _14912_, _38997_);
  and _59925_ (_36862_[1], _14913_, _14911_);
  nor _59926_ (_36863_[15], _13732_, rst);
  nor _59927_ (_14914_, _13534_, _13543_);
  and _59928_ (_14915_, _13534_, _13543_);
  or _59929_ (_14916_, _14915_, _14914_);
  and _59930_ (_36862_[0], _14916_, _38997_);
  and _59931_ (_36863_[0], _13621_, _38997_);
  and _59932_ (_36863_[1], _14313_, _38997_);
  and _59933_ (_36863_[2], _14374_, _38997_);
  and _59934_ (_36863_[3], _14435_, _38997_);
  and _59935_ (_36863_[4], _14506_, _38997_);
  and _59936_ (_36863_[5], _14581_, _38997_);
  and _59937_ (_36863_[6], _14642_, _38997_);
  and _59938_ (_36863_[7], _14151_, _38997_);
  and _59939_ (_36863_[8], _13743_, _38997_);
  and _59940_ (_36863_[9], _13747_, _38997_);
  and _59941_ (_36863_[10], _13752_, _38997_);
  and _59942_ (_36863_[11], _13784_, _38997_);
  and _59943_ (_36863_[12], _13755_, _38997_);
  and _59944_ (_36863_[13], _13738_, _38997_);
  and _59945_ (_36863_[14], _13735_, _38997_);
  nor _59946_ (_36867_[2], _33497_, rst);
  and _59947_ (_14917_, _33387_, _33410_);
  and _59948_ (_14918_, _33371_, _33252_);
  nor _59949_ (_14919_, _14918_, _14917_);
  and _59950_ (_14920_, _33371_, _33385_);
  not _59951_ (_14921_, _14920_);
  and _59952_ (_14922_, _14921_, _14919_);
  and _59953_ (_14923_, _33135_, _38997_);
  not _59954_ (_14924_, _14923_);
  or _59955_ (_14925_, _14924_, _14917_);
  or _59956_ (_36868_[2], _14925_, _14922_);
  and _59957_ (_14926_, _33197_, _33172_);
  not _59958_ (_14927_, _33222_);
  nor _59959_ (_14928_, _33246_, _14927_);
  and _59960_ (_14929_, _14928_, _14926_);
  not _59961_ (_14930_, _33295_);
  not _59962_ (_14931_, _33319_);
  and _59963_ (_14932_, _33344_, _14931_);
  and _59964_ (_14933_, _14932_, _14930_);
  and _59965_ (_14934_, _14933_, _14929_);
  not _59966_ (_14935_, _33271_);
  nor _59967_ (_14936_, _33197_, _14935_);
  and _59968_ (_14937_, _14932_, _33295_);
  and _59969_ (_14938_, _14937_, _14936_);
  not _59970_ (_14939_, _33246_);
  not _59971_ (_14940_, _33172_);
  and _59972_ (_14941_, _33197_, _14940_);
  and _59973_ (_14942_, _14941_, _14939_);
  nor _59974_ (_14943_, _33344_, _33319_);
  nor _59975_ (_14944_, _33295_, _14935_);
  and _59976_ (_14945_, _14944_, _14943_);
  and _59977_ (_14946_, _14945_, _14942_);
  or _59978_ (_14947_, _14946_, _14938_);
  nor _59979_ (_14948_, _14947_, _14934_);
  and _59980_ (_14949_, _14943_, _14930_);
  and _59981_ (_14950_, _33246_, _33271_);
  and _59982_ (_14951_, _14950_, _14941_);
  or _59983_ (_14952_, _14951_, _14936_);
  and _59984_ (_14953_, _14952_, _14949_);
  and _59985_ (_14954_, _33344_, _33319_);
  and _59986_ (_14955_, _14954_, _33271_);
  and _59987_ (_14956_, _14955_, _14929_);
  nor _59988_ (_14957_, _14956_, _14953_);
  nand _59989_ (_14958_, _14957_, _14948_);
  and _59990_ (_14959_, _14941_, _14928_);
  and _59991_ (_14960_, _14959_, _14935_);
  and _59992_ (_14961_, _14960_, _14943_);
  and _59993_ (_14962_, _33295_, _14935_);
  and _59994_ (_14963_, _14962_, _14943_);
  and _59995_ (_14964_, _14963_, _14929_);
  and _59996_ (_14965_, _14926_, _33246_);
  and _59997_ (_14966_, _14965_, _33222_);
  nor _59998_ (_14967_, _33344_, _14931_);
  and _59999_ (_14968_, _14967_, _33295_);
  and _60000_ (_14969_, _14968_, _14966_);
  nor _60001_ (_14970_, _14969_, _14964_);
  not _60002_ (_14971_, _14970_);
  or _60003_ (_14972_, _14971_, _14961_);
  or _60004_ (_14973_, _14972_, _14958_);
  and _60005_ (_14974_, _33295_, _33271_);
  and _60006_ (_14975_, _14967_, _14974_);
  nor _60007_ (_14976_, _33295_, _33271_);
  and _60008_ (_14977_, _14967_, _14976_);
  or _60009_ (_14978_, _14977_, _14975_);
  and _60010_ (_14979_, _14978_, _14929_);
  and _60011_ (_14980_, _14974_, _14932_);
  and _60012_ (_14981_, _14942_, _14927_);
  and _60013_ (_14982_, _14981_, _14980_);
  nor _60014_ (_14983_, _14982_, _14979_);
  and _60015_ (_14984_, _14926_, _14939_);
  not _60016_ (_14985_, _14984_);
  and _60017_ (_14986_, _14976_, _14954_);
  nor _60018_ (_14987_, _14986_, _14927_);
  nor _60019_ (_14988_, _14987_, _14985_);
  not _60020_ (_14989_, _14988_);
  and _60021_ (_14990_, _14962_, _14954_);
  and _60022_ (_14991_, _14990_, _14929_);
  and _60023_ (_14992_, _14967_, _14944_);
  and _60024_ (_14993_, _14992_, _14929_);
  nor _60025_ (_14994_, _14993_, _14991_);
  and _60026_ (_14995_, _14994_, _14989_);
  and _60027_ (_14996_, _14954_, _14944_);
  and _60028_ (_14997_, _14965_, _14927_);
  and _60029_ (_14998_, _14997_, _14996_);
  and _60030_ (_14999_, _14967_, _14930_);
  and _60031_ (_15000_, _14999_, _14966_);
  or _60032_ (_15001_, _15000_, _14998_);
  and _60033_ (_15002_, _14943_, _33295_);
  and _60034_ (_15003_, _14997_, _15002_);
  and _60035_ (_15004_, _14965_, _14933_);
  or _60036_ (_15005_, _15004_, _15003_);
  nor _60037_ (_15006_, _15005_, _15001_);
  and _60038_ (_15007_, _15006_, _14995_);
  nand _60039_ (_15008_, _15007_, _14983_);
  or _60040_ (_15009_, _15008_, _14973_);
  and _60041_ (_15010_, _15009_, _33136_);
  not _60042_ (_15011_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _60043_ (_15012_, _33134_, _33129_);
  and _60044_ (_15013_, _15012_, _33456_);
  nor _60045_ (_15014_, _15013_, _15011_);
  or _60046_ (_15015_, _15014_, rst);
  or _60047_ (_36869_[1], _15015_, _15010_);
  nand _60048_ (_15016_, _33319_, _33130_);
  or _60049_ (_15017_, _33130_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _60050_ (_15018_, _15017_, _38997_);
  and _60051_ (_36870_[7], _15018_, _15016_);
  and _60052_ (_15019_, \oc8051_top_1.oc8051_sfr1.wait_data , _38997_);
  and _60053_ (_15020_, _15019_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _60054_ (_15021_, _33252_, _33381_);
  nor _60055_ (_15022_, _15021_, _33459_);
  and _60056_ (_15023_, _33423_, _33410_);
  nor _60057_ (_15024_, _15023_, _34354_);
  nand _60058_ (_15025_, _15024_, _15022_);
  and _60059_ (_15026_, _33388_, _33410_);
  and _60060_ (_15027_, _33478_, _33372_);
  or _60061_ (_15028_, _15027_, _15026_);
  and _60062_ (_15029_, _33388_, _33252_);
  nor _60063_ (_15030_, _15029_, _34349_);
  nand _60064_ (_15031_, _15030_, _33362_);
  or _60065_ (_15032_, _15031_, _15028_);
  or _60066_ (_15033_, _15032_, _15025_);
  and _60067_ (_15034_, _15033_, _14923_);
  or _60068_ (_36871_, _15034_, _15020_);
  not _60069_ (_15035_, _33485_);
  and _60070_ (_15036_, _33437_, _33252_);
  or _60071_ (_15037_, _15036_, _15035_);
  and _60072_ (_15038_, _33443_, _33417_);
  or _60073_ (_15039_, _15038_, _33521_);
  and _60074_ (_15040_, _33365_, _33366_);
  and _60075_ (_15041_, _15040_, _33423_);
  or _60076_ (_15042_, _15041_, _15039_);
  or _60077_ (_15043_, _15042_, _15037_);
  and _60078_ (_15044_, _15043_, _33135_);
  and _60079_ (_15045_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _60080_ (_15046_, _33467_, _15011_);
  not _60081_ (_15047_, _33481_);
  and _60082_ (_15048_, _15047_, _15046_);
  or _60083_ (_15049_, _15048_, _15045_);
  or _60084_ (_15050_, _15049_, _15044_);
  and _60085_ (_36872_[1], _15050_, _38997_);
  and _60086_ (_15051_, _15019_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _60087_ (_15052_, _33478_, _33395_);
  or _60088_ (_15053_, _33395_, _33418_);
  and _60089_ (_15054_, _15053_, _33368_);
  or _60090_ (_15055_, _15054_, _15052_);
  and _60091_ (_15056_, _15040_, _33359_);
  or _60092_ (_15057_, _15056_, _15055_);
  and _60093_ (_15058_, _15053_, _33201_);
  and _60094_ (_15059_, _33201_, _33275_);
  and _60095_ (_15060_, _15059_, _33358_);
  or _60096_ (_15061_, _15060_, _15058_);
  and _60097_ (_15062_, _15059_, _33375_);
  nor _60098_ (_15063_, _15062_, _33504_);
  not _60099_ (_15064_, _15063_);
  and _60100_ (_15065_, _33374_, _33275_);
  and _60101_ (_15066_, _33478_, _15065_);
  or _60102_ (_15067_, _15066_, _33506_);
  or _60103_ (_15068_, _15067_, _15064_);
  or _60104_ (_15069_, _15068_, _15037_);
  or _60105_ (_15070_, _15069_, _15061_);
  or _60106_ (_15071_, _15070_, _15057_);
  and _60107_ (_15072_, _15071_, _14923_);
  or _60108_ (_36873_[1], _15072_, _15051_);
  and _60109_ (_15073_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _60110_ (_15074_, _33436_, _33135_);
  or _60111_ (_15075_, _15074_, _15073_);
  or _60112_ (_15076_, _15075_, _15048_);
  and _60113_ (_36874_[2], _15076_, _38997_);
  and _60114_ (_15077_, _33367_, _33202_);
  and _60115_ (_15078_, _33391_, _33358_);
  nor _60116_ (_15079_, _15078_, _15077_);
  nor _60117_ (_15080_, _15079_, _33354_);
  and _60118_ (_15081_, _15026_, _33131_);
  nor _60119_ (_15082_, _15081_, _15080_);
  nor _60120_ (_15083_, _15082_, _33467_);
  nor _60121_ (_15084_, _14917_, _33354_);
  nor _60122_ (_15085_, _15084_, _14922_);
  and _60123_ (_15086_, _15085_, _15046_);
  or _60124_ (_15087_, _15086_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _60125_ (_15088_, _15087_, _15083_);
  or _60126_ (_15089_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _33129_);
  and _60127_ (_15090_, _15089_, _38997_);
  and _60128_ (_36875_[2], _15090_, _15088_);
  and _60129_ (_15091_, _15019_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or _60130_ (_15092_, _15060_, _15035_);
  and _60131_ (_15093_, _33418_, _33201_);
  or _60132_ (_15094_, _15093_, _33419_);
  or _60133_ (_15095_, _15094_, _15092_);
  or _60134_ (_15096_, _34356_, _34354_);
  or _60135_ (_15097_, _15096_, _33434_);
  or _60136_ (_15098_, _33359_, _33423_);
  and _60137_ (_15099_, _15098_, _33398_);
  or _60138_ (_15100_, _15056_, _15038_);
  or _60139_ (_15101_, _15100_, _34348_);
  or _60140_ (_15102_, _15101_, _15099_);
  or _60141_ (_15103_, _15102_, _15097_);
  or _60142_ (_15104_, _15103_, _15095_);
  and _60143_ (_15105_, _15104_, _14923_);
  or _60144_ (_36876_[1], _15105_, _15091_);
  and _60145_ (_15106_, _15019_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _60146_ (_15107_, _33398_, _33418_);
  not _60147_ (_15108_, _33511_);
  and _60148_ (_15109_, _33515_, _33380_);
  or _60149_ (_15110_, _15109_, _15108_);
  or _60150_ (_15111_, _15110_, _15107_);
  and _60151_ (_15112_, _15040_, _33429_);
  and _60152_ (_15113_, _33349_, _33410_);
  or _60153_ (_15114_, _15113_, _15041_);
  or _60154_ (_15115_, _15114_, _15112_);
  or _60155_ (_15116_, _15115_, _15061_);
  or _60156_ (_15117_, _15116_, _15111_);
  and _60157_ (_15118_, _33403_, _33465_);
  or _60158_ (_15119_, _15118_, _33411_);
  or _60159_ (_15120_, _15119_, _34359_);
  and _60160_ (_15121_, _33478_, _33403_);
  or _60161_ (_15122_, _15121_, _15120_);
  and _60162_ (_15123_, _33443_, _33380_);
  and _60163_ (_15124_, _33443_, _33407_);
  or _60164_ (_15125_, _15124_, _15123_);
  or _60165_ (_15126_, _33506_, _33430_);
  or _60166_ (_15127_, _33416_, _33406_);
  or _60167_ (_15128_, _15127_, _15126_);
  or _60168_ (_15129_, _15128_, _15125_);
  or _60169_ (_15130_, _15129_, _15057_);
  or _60170_ (_15131_, _15130_, _15122_);
  or _60171_ (_15132_, _15131_, _15117_);
  and _60172_ (_15133_, _15132_, _14923_);
  or _60173_ (_36877_[3], _15133_, _15106_);
  and _60174_ (_15134_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nor _60175_ (_15135_, _33481_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _60176_ (_15136_, _15135_, _15134_);
  and _60177_ (_15137_, _15136_, _38997_);
  and _60178_ (_15138_, _33398_, _33350_);
  and _60179_ (_15139_, _15059_, _33387_);
  or _60180_ (_15140_, _15139_, _15138_);
  and _60181_ (_15141_, _15040_, _33350_);
  or _60182_ (_15142_, _15141_, _15140_);
  and _60183_ (_15143_, _15040_, _33437_);
  and _60184_ (_15144_, _33350_, _33201_);
  or _60185_ (_15145_, _15144_, _33522_);
  or _60186_ (_15146_, _15145_, _15143_);
  or _60187_ (_15147_, _15146_, _15142_);
  and _60188_ (_15148_, _15147_, _14923_);
  or _60189_ (_36878_[1], _15148_, _15137_);
  or _60190_ (_15149_, _34351_, _33436_);
  or _60191_ (_15150_, _15149_, _34350_);
  or _60192_ (_15151_, _15054_, _33432_);
  or _60193_ (_15152_, _15151_, _15150_);
  or _60194_ (_15153_, _34355_, _33434_);
  and _60195_ (_15154_, _33359_, _33465_);
  and _60196_ (_15155_, _33370_, _33275_);
  and _60197_ (_15156_, _15155_, _33368_);
  or _60198_ (_15157_, _15156_, _33420_);
  or _60199_ (_15158_, _15157_, _15154_);
  or _60200_ (_15159_, _15158_, _15119_);
  or _60201_ (_15160_, _15159_, _15153_);
  or _60202_ (_15161_, _15160_, _15152_);
  and _60203_ (_15162_, _33397_, _33201_);
  and _60204_ (_15163_, _15059_, _33370_);
  or _60205_ (_15164_, _15163_, _15162_);
  or _60206_ (_15165_, _15164_, _15039_);
  or _60207_ (_15166_, _15165_, _15061_);
  and _60208_ (_15167_, _33398_, _33275_);
  and _60209_ (_15168_, _15167_, _33370_);
  or _60210_ (_15169_, _15168_, _33506_);
  or _60211_ (_15170_, _15169_, _33399_);
  and _60212_ (_15171_, _33388_, _33201_);
  and _60213_ (_15172_, _15077_, _33275_);
  or _60214_ (_15173_, _15172_, _33507_);
  or _60215_ (_15174_, _15173_, _15171_);
  or _60216_ (_15175_, _15174_, _33386_);
  or _60217_ (_15176_, _15175_, _15170_);
  or _60218_ (_15177_, _15176_, _15166_);
  or _60219_ (_15178_, _15177_, _15161_);
  and _60220_ (_15179_, _15178_, _33135_);
  and _60221_ (_15180_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and _60222_ (_15181_, _33461_, _33359_);
  and _60223_ (_15182_, _15080_, _33458_);
  or _60224_ (_15183_, _15182_, _15048_);
  or _60225_ (_15184_, _15183_, _15181_);
  or _60226_ (_15185_, _15184_, _15180_);
  or _60227_ (_15186_, _15185_, _15179_);
  and _60228_ (_36879_, _15186_, _38997_);
  and _60229_ (_36867_[0], _33530_, _38997_);
  and _60230_ (_36867_[1], _33472_, _38997_);
  nand _60231_ (_36868_[0], _15085_, _14923_);
  or _60232_ (_36868_[1], _14924_, _14919_);
  or _60233_ (_15187_, _15000_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _60234_ (_15188_, _15187_, _15003_);
  or _60235_ (_15189_, _15188_, _14961_);
  and _60236_ (_15190_, _15189_, _15013_);
  nor _60237_ (_15191_, _15012_, _33456_);
  or _60238_ (_15192_, _15191_, rst);
  or _60239_ (_36869_[0], _15192_, _15190_);
  nand _60240_ (_15193_, _33222_, _33130_);
  or _60241_ (_15194_, _33130_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _60242_ (_15195_, _15194_, _38997_);
  and _60243_ (_36870_[0], _15195_, _15193_);
  or _60244_ (_15196_, _33246_, _33490_);
  or _60245_ (_15197_, _33130_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _60246_ (_15198_, _15197_, _38997_);
  and _60247_ (_36870_[1], _15198_, _15196_);
  nand _60248_ (_15199_, _33172_, _33130_);
  or _60249_ (_15200_, _33130_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _60250_ (_15201_, _15200_, _38997_);
  and _60251_ (_36870_[2], _15201_, _15199_);
  nand _60252_ (_15202_, _33197_, _33130_);
  or _60253_ (_15203_, _33130_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _60254_ (_15204_, _15203_, _38997_);
  and _60255_ (_36870_[3], _15204_, _15202_);
  or _60256_ (_15205_, _33271_, _33490_);
  or _60257_ (_15206_, _33130_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _60258_ (_15207_, _15206_, _38997_);
  and _60259_ (_36870_[4], _15207_, _15205_);
  nand _60260_ (_15208_, _33295_, _33130_);
  or _60261_ (_15209_, _33130_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _60262_ (_15210_, _15209_, _38997_);
  and _60263_ (_36870_[5], _15210_, _15208_);
  or _60264_ (_15211_, _33344_, _33490_);
  or _60265_ (_15212_, _33130_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _60266_ (_15213_, _15212_, _38997_);
  and _60267_ (_36870_[6], _15213_, _15211_);
  and _60268_ (_15214_, _15059_, _33381_);
  or _60269_ (_15215_, _15214_, _15144_);
  or _60270_ (_15216_, _15215_, _15143_);
  or _60271_ (_15217_, _33359_, _33418_);
  and _60272_ (_15218_, _15217_, _33478_);
  or _60273_ (_15219_, _15218_, _15052_);
  and _60274_ (_15220_, _33478_, _33408_);
  and _60275_ (_15221_, _33371_, _33275_);
  and _60276_ (_15222_, _15221_, _33478_);
  and _60277_ (_15223_, _15040_, _33382_);
  or _60278_ (_15224_, _15223_, _15222_);
  or _60279_ (_15225_, _15224_, _15220_);
  or _60280_ (_15226_, _15225_, _15219_);
  or _60281_ (_15227_, _15226_, _15216_);
  and _60282_ (_15228_, _15040_, _33403_);
  or _60283_ (_15229_, _15228_, _15036_);
  and _60284_ (_15230_, _33443_, _33371_);
  and _60285_ (_15231_, _33443_, _33381_);
  or _60286_ (_15232_, _15231_, _33522_);
  or _60287_ (_15233_, _15232_, _15230_);
  or _60288_ (_15234_, _15233_, _15142_);
  or _60289_ (_15235_, _15234_, _15229_);
  or _60290_ (_15236_, _15124_, _15112_);
  and _60291_ (_15237_, _15167_, _33381_);
  and _60292_ (_15238_, _15040_, _33372_);
  or _60293_ (_15239_, _15238_, _15237_);
  or _60294_ (_15240_, _15239_, _15236_);
  nand _60295_ (_15241_, _33511_, _33485_);
  not _60296_ (_15242_, _33518_);
  or _60297_ (_15243_, _15113_, _15242_);
  or _60298_ (_15244_, _15243_, _15241_);
  or _60299_ (_15245_, _15244_, _15240_);
  or _60300_ (_15246_, _15245_, _15235_);
  or _60301_ (_15247_, _15246_, _15227_);
  and _60302_ (_15248_, _15247_, _33135_);
  and _60303_ (_15249_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _60304_ (_15250_, _15249_, _15086_);
  or _60305_ (_15251_, _15250_, _15248_);
  and _60306_ (_36872_[0], _15251_, _38997_);
  and _60307_ (_15252_, _15019_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _60308_ (_15253_, _15125_, _15028_);
  and _60309_ (_15254_, _33478_, _33383_);
  or _60310_ (_15255_, _15254_, _15229_);
  or _60311_ (_15256_, _15255_, _15253_);
  and _60312_ (_15257_, _33429_, _33465_);
  and _60313_ (_15258_, _33478_, _33429_);
  or _60314_ (_15259_, _15258_, _15064_);
  or _60315_ (_15260_, _15259_, _15257_);
  or _60316_ (_15261_, _15066_, _15118_);
  or _60317_ (_15262_, _15261_, _33435_);
  or _60318_ (_15263_, _15262_, _15260_);
  or _60319_ (_15264_, _15263_, _15111_);
  or _60320_ (_15265_, _15264_, _15256_);
  and _60321_ (_15266_, _15265_, _14923_);
  or _60322_ (_36873_[0], _15266_, _15252_);
  or _60323_ (_15267_, _15175_, _15161_);
  and _60324_ (_15268_, _15267_, _33135_);
  and _60325_ (_15269_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _60326_ (_15270_, _15269_, _15184_);
  or _60327_ (_15271_, _15270_, _15268_);
  and _60328_ (_36874_[0], _15271_, _38997_);
  and _60329_ (_15272_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _60330_ (_15273_, _15272_, _15183_);
  nand _60331_ (_15274_, _33431_, _33354_);
  nand _60332_ (_15275_, _15274_, _33520_);
  or _60333_ (_15276_, _15275_, _15080_);
  or _60334_ (_15277_, _15276_, _15170_);
  and _60335_ (_15278_, _15277_, _33135_);
  or _60336_ (_15279_, _15278_, _15273_);
  and _60337_ (_36874_[1], _15279_, _38997_);
  or _60338_ (_15280_, _14917_, _33480_);
  and _60339_ (_15281_, _15141_, _33275_);
  or _60340_ (_15282_, _15281_, _15223_);
  or _60341_ (_15283_, _15282_, _15280_);
  or _60342_ (_15284_, _15220_, _15258_);
  and _60343_ (_15285_, _15221_, _33368_);
  and _60344_ (_15286_, _15141_, _33354_);
  or _60345_ (_15287_, _15286_, _15285_);
  or _60346_ (_15288_, _15287_, _15284_);
  or _60347_ (_15289_, _15288_, _15080_);
  or _60348_ (_15290_, _15289_, _15283_);
  and _60349_ (_15291_, _15040_, _33376_);
  or _60350_ (_15292_, _15291_, _15027_);
  or _60351_ (_15293_, _15222_, _33479_);
  or _60352_ (_15294_, _15293_, _15292_);
  or _60353_ (_15295_, _15294_, _15219_);
  and _60354_ (_15296_, _33478_, _33423_);
  or _60355_ (_15297_, _15113_, _15296_);
  or _60356_ (_15298_, _15297_, _15216_);
  nor _60357_ (_15299_, _15163_, _33522_);
  nand _60358_ (_15300_, _15299_, _33484_);
  or _60359_ (_15301_, _15168_, _15121_);
  or _60360_ (_15302_, _15301_, _15300_);
  or _60361_ (_15303_, _15140_, _15237_);
  and _60362_ (_15304_, _33386_, _33464_);
  or _60363_ (_15305_, _15304_, _15303_);
  or _60364_ (_15306_, _15305_, _15302_);
  or _60365_ (_15307_, _15306_, _15298_);
  or _60366_ (_15308_, _15307_, _15295_);
  or _60367_ (_15309_, _15308_, _15290_);
  and _60368_ (_15310_, _15309_, _33135_);
  and _60369_ (_15311_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _60370_ (_15312_, _33481_, _33131_);
  and _60371_ (_15313_, _33372_, _33252_);
  or _60372_ (_15314_, _15026_, _33482_);
  nor _60373_ (_15315_, _33201_, _33275_);
  and _60374_ (_15316_, _33371_, _33389_);
  and _60375_ (_15317_, _15316_, _15315_);
  or _60376_ (_15318_, _15317_, _15314_);
  or _60377_ (_15319_, _15318_, _15313_);
  and _60378_ (_15320_, _15319_, _15046_);
  or _60379_ (_15321_, _15320_, _15312_);
  or _60380_ (_15322_, _15321_, _15311_);
  or _60381_ (_15323_, _15322_, _15310_);
  and _60382_ (_36875_[0], _15323_, _38997_);
  and _60383_ (_15324_, _15059_, _33371_);
  or _60384_ (_15325_, _15156_, _15036_);
  or _60385_ (_15326_, _15325_, _15324_);
  or _60386_ (_15327_, _15326_, _33384_);
  or _60387_ (_15328_, _15327_, _15303_);
  and _60388_ (_15329_, _33429_, _33410_);
  and _60389_ (_15330_, _15221_, _33398_);
  or _60390_ (_15331_, _15330_, _33386_);
  or _60391_ (_15332_, _15331_, _15329_);
  or _60392_ (_15333_, _33522_, _33480_);
  or _60393_ (_15334_, _15333_, _33482_);
  not _60394_ (_15335_, _33484_);
  or _60395_ (_15336_, _15335_, _33411_);
  or _60396_ (_15337_, _15336_, _15334_);
  or _60397_ (_15338_, _15337_, _15332_);
  or _60398_ (_15339_, _15338_, _15328_);
  or _60399_ (_15340_, _15298_, _15295_);
  or _60400_ (_15341_, _15340_, _15339_);
  and _60401_ (_15342_, _15341_, _33135_);
  and _60402_ (_15343_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _60403_ (_15344_, _15343_, _15321_);
  or _60404_ (_15345_, _15344_, _15342_);
  and _60405_ (_36875_[1], _15345_, _38997_);
  and _60406_ (_15346_, _15019_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _60407_ (_15347_, _15095_, _34362_);
  or _60408_ (_15348_, _15347_, _15153_);
  or _60409_ (_15349_, _33410_, _33201_);
  and _60410_ (_15350_, _15349_, _33351_);
  and _60411_ (_15351_, _33478_, _33418_);
  and _60412_ (_15352_, _33376_, _33410_);
  or _60413_ (_15353_, _15352_, _15351_);
  and _60414_ (_15354_, _15217_, _33410_);
  or _60415_ (_15355_, _15354_, _15353_);
  or _60416_ (_15356_, _15355_, _15350_);
  and _60417_ (_15357_, _15167_, _33350_);
  or _60418_ (_15358_, _15281_, _15357_);
  or _60419_ (_15359_, _15139_, _15038_);
  or _60420_ (_15360_, _15143_, _15056_);
  or _60421_ (_15361_, _15360_, _15359_);
  or _60422_ (_15362_, _15361_, _15358_);
  or _60423_ (_15363_, _33522_, _34351_);
  or _60424_ (_15364_, _15363_, _15099_);
  or _60425_ (_15365_, _15364_, _15362_);
  or _60426_ (_15366_, _15365_, _15356_);
  or _60427_ (_15367_, _15366_, _15348_);
  and _60428_ (_15368_, _15367_, _14923_);
  or _60429_ (_36876_[0], _15368_, _15346_);
  or _60430_ (_15369_, _15109_, _15041_);
  or _60431_ (_15370_, _15286_, _15107_);
  or _60432_ (_15371_, _15370_, _15369_);
  nor _60433_ (_15372_, _15123_, _33404_);
  nand _60434_ (_15373_, _15372_, _33486_);
  or _60435_ (_15374_, _15373_, _15371_);
  and _60436_ (_15375_, _33359_, _33410_);
  and _60437_ (_15376_, _33351_, _33410_);
  or _60438_ (_15377_, _15351_, _15376_);
  or _60439_ (_15378_, _15377_, _15375_);
  or _60440_ (_15379_, _15378_, _15283_);
  or _60441_ (_15380_, _15379_, _15374_);
  nor _60442_ (_15381_, _34358_, _33386_);
  not _60443_ (_15382_, _15381_);
  or _60444_ (_15383_, _33503_, _15382_);
  or _60445_ (_15384_, _15383_, _15215_);
  or _60446_ (_15385_, _15384_, _15122_);
  or _60447_ (_15386_, _15385_, _15380_);
  and _60448_ (_15387_, _15386_, _14923_);
  and _60449_ (_15388_, _15019_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _60450_ (_15389_, _33492_, _38997_);
  or _60451_ (_15390_, _15389_, _15388_);
  or _60452_ (_36877_[0], _15390_, _15387_);
  and _60453_ (_15391_, _33350_, _33410_);
  or _60454_ (_15392_, _15391_, _15361_);
  or _60455_ (_15393_, _33504_, _33405_);
  or _60456_ (_15394_, _15393_, _15062_);
  not _60457_ (_15395_, _33523_);
  or _60458_ (_15396_, _15041_, _15395_);
  or _60459_ (_15397_, _15396_, _15394_);
  or _60460_ (_15398_, _15397_, _15392_);
  not _60461_ (_15399_, _15223_);
  and _60462_ (_15400_, _15399_, _15381_);
  not _60463_ (_15401_, _15400_);
  or _60464_ (_15402_, _15401_, _15055_);
  or _60465_ (_15403_, _15402_, _15398_);
  or _60466_ (_15404_, _15214_, _15061_);
  or _60467_ (_15405_, _15222_, _34347_);
  or _60468_ (_15406_, _15405_, _15292_);
  nor _60469_ (_15407_, _33506_, _15237_);
  not _60470_ (_15408_, _15407_);
  or _60471_ (_15409_, _15408_, _15406_);
  or _60472_ (_15410_, _15409_, _15404_);
  or _60473_ (_15411_, _15410_, _15403_);
  and _60474_ (_15412_, _15411_, _33135_);
  and _60475_ (_15413_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _60476_ (_15414_, _15413_, _33491_);
  or _60477_ (_15415_, _15414_, _15412_);
  and _60478_ (_36877_[1], _15415_, _38997_);
  and _60479_ (_15416_, _33358_, _33410_);
  or _60480_ (_15417_, _15039_, _33434_);
  or _60481_ (_15418_, _15417_, _15416_);
  or _60482_ (_15419_, _15418_, _15055_);
  or _60483_ (_15420_, _15419_, _15401_);
  or _60484_ (_15421_, _33479_, _33416_);
  or _60485_ (_15422_, _15421_, _33420_);
  or _60486_ (_15423_, _15422_, _15218_);
  or _60487_ (_15424_, _15408_, _15405_);
  or _60488_ (_15425_, _15424_, _15423_);
  or _60489_ (_15426_, _15425_, _15404_);
  or _60490_ (_15427_, _15426_, _15420_);
  and _60491_ (_15428_, _15427_, _14923_);
  and _60492_ (_15429_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _60493_ (_15430_, _15429_, _33493_);
  and _60494_ (_15431_, _15430_, _38997_);
  or _60495_ (_36877_[2], _15431_, _15428_);
  and _60496_ (_15432_, _15019_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not _60497_ (_15433_, _33202_);
  and _60498_ (_15434_, _33376_, _15433_);
  or _60499_ (_15435_, _15434_, _34356_);
  or _60500_ (_15436_, _15376_, _15023_);
  or _60501_ (_15437_, _15436_, _15435_);
  or _60502_ (_15438_, _15437_, _15355_);
  or _60503_ (_15439_, _15147_, _34362_);
  or _60504_ (_15440_, _15439_, _15438_);
  and _60505_ (_15441_, _15440_, _14923_);
  or _60506_ (_36878_[0], _15441_, _15432_);
  nor _60507_ (_36864_[7], _33319_, rst);
  nor _60508_ (_36865_[7], _34342_, rst);
  and _60509_ (_15442_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and _60510_ (_15443_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and _60511_ (_15444_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _60512_ (_15445_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _60513_ (_15446_, _15445_, _15444_);
  and _60514_ (_15447_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _60515_ (_15448_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _60516_ (_15449_, _15448_, _15447_);
  and _60517_ (_15450_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  not _60518_ (_15451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _60519_ (_15452_, _33146_, _15451_);
  nor _60520_ (_15453_, _15452_, _15450_);
  and _60521_ (_15454_, _15453_, _15449_);
  and _60522_ (_15455_, _15454_, _15446_);
  nor _60523_ (_15456_, _15455_, _33140_);
  nor _60524_ (_15457_, _15456_, _15443_);
  nor _60525_ (_15458_, _15457_, _34325_);
  nor _60526_ (_15459_, _15458_, _15442_);
  nor _60527_ (_36866_[7], _15459_, rst);
  nor _60528_ (_36864_[0], _33222_, rst);
  and _60529_ (_36864_[1], _33246_, _38997_);
  nor _60530_ (_36864_[2], _33172_, rst);
  nor _60531_ (_36864_[3], _33197_, rst);
  and _60532_ (_36864_[4], _33271_, _38997_);
  nor _60533_ (_36864_[5], _33295_, rst);
  and _60534_ (_36864_[6], _33344_, _38997_);
  nor _60535_ (_36865_[0], _34457_, rst);
  nor _60536_ (_36865_[1], _34575_, rst);
  nor _60537_ (_36865_[2], _34757_, rst);
  nor _60538_ (_36865_[3], _34417_, rst);
  nor _60539_ (_36865_[4], _34495_, rst);
  nor _60540_ (_36865_[5], _34603_, rst);
  nor _60541_ (_36865_[6], _34685_, rst);
  and _60542_ (_15460_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and _60543_ (_15461_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _60544_ (_15462_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _60545_ (_15463_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _60546_ (_15464_, _15463_, _15462_);
  and _60547_ (_15465_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _60548_ (_15466_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _60549_ (_15467_, _15466_, _15465_);
  and _60550_ (_15468_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  not _60551_ (_15469_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _60552_ (_15470_, _33146_, _15469_);
  nor _60553_ (_15471_, _15470_, _15468_);
  and _60554_ (_15472_, _15471_, _15467_);
  and _60555_ (_15473_, _15472_, _15464_);
  nor _60556_ (_15474_, _15473_, _33140_);
  nor _60557_ (_15475_, _15474_, _15461_);
  nor _60558_ (_15476_, _15475_, _34325_);
  nor _60559_ (_15477_, _15476_, _15460_);
  nor _60560_ (_36866_[0], _15477_, rst);
  and _60561_ (_15478_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and _60562_ (_15479_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and _60563_ (_15480_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _60564_ (_15481_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _60565_ (_15482_, _15481_, _15480_);
  and _60566_ (_15483_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _60567_ (_15484_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _60568_ (_15485_, _15484_, _15483_);
  and _60569_ (_15486_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _60570_ (_15487_, _33236_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _60571_ (_15488_, _15487_, _15486_);
  and _60572_ (_15489_, _15488_, _15485_);
  and _60573_ (_15490_, _15489_, _15482_);
  nor _60574_ (_15491_, _15490_, _33140_);
  nor _60575_ (_15492_, _15491_, _15479_);
  nor _60576_ (_15493_, _15492_, _34325_);
  nor _60577_ (_15494_, _15493_, _15478_);
  nor _60578_ (_36866_[1], _15494_, rst);
  and _60579_ (_15495_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and _60580_ (_15496_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and _60581_ (_15497_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _60582_ (_15498_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _60583_ (_15499_, _15498_, _15497_);
  and _60584_ (_15500_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  not _60585_ (_15501_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _60586_ (_15502_, _33146_, _15501_);
  nor _60587_ (_15503_, _15502_, _15500_);
  and _60588_ (_15504_, _15503_, _15499_);
  and _60589_ (_15505_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _60590_ (_15506_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _60591_ (_15507_, _15506_, _15505_);
  and _60592_ (_15508_, _15507_, _15504_);
  nor _60593_ (_15509_, _15508_, _33140_);
  nor _60594_ (_15510_, _15509_, _15496_);
  nor _60595_ (_15511_, _15510_, _34325_);
  nor _60596_ (_15512_, _15511_, _15495_);
  nor _60597_ (_36866_[2], _15512_, rst);
  and _60598_ (_15513_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and _60599_ (_15514_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and _60600_ (_15515_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _60601_ (_15516_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _60602_ (_15517_, _15516_, _15515_);
  and _60603_ (_15518_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _60604_ (_15519_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _60605_ (_15520_, _15519_, _15518_);
  and _60606_ (_15521_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  not _60607_ (_15522_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _60608_ (_15523_, _33146_, _15522_);
  nor _60609_ (_15524_, _15523_, _15521_);
  and _60610_ (_15525_, _15524_, _15520_);
  and _60611_ (_15526_, _15525_, _15517_);
  nor _60612_ (_15527_, _15526_, _33140_);
  nor _60613_ (_15528_, _15527_, _15514_);
  nor _60614_ (_15529_, _15528_, _34325_);
  nor _60615_ (_15530_, _15529_, _15513_);
  nor _60616_ (_36866_[3], _15530_, rst);
  and _60617_ (_15531_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and _60618_ (_15532_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and _60619_ (_15533_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _60620_ (_15534_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _60621_ (_15535_, _15534_, _15533_);
  and _60622_ (_15536_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _60623_ (_15537_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _60624_ (_15538_, _15537_, _15536_);
  and _60625_ (_15539_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  not _60626_ (_15540_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _60627_ (_15541_, _33146_, _15540_);
  nor _60628_ (_15542_, _15541_, _15539_);
  and _60629_ (_15543_, _15542_, _15538_);
  and _60630_ (_15544_, _15543_, _15535_);
  nor _60631_ (_15545_, _15544_, _33140_);
  nor _60632_ (_15546_, _15545_, _15532_);
  nor _60633_ (_15547_, _15546_, _34325_);
  nor _60634_ (_15548_, _15547_, _15531_);
  nor _60635_ (_36866_[4], _15548_, rst);
  and _60636_ (_15549_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and _60637_ (_15550_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and _60638_ (_15551_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _60639_ (_15552_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _60640_ (_15553_, _15552_, _15551_);
  and _60641_ (_15554_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  not _60642_ (_15555_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _60643_ (_15556_, _33146_, _15555_);
  nor _60644_ (_15557_, _15556_, _15554_);
  and _60645_ (_15558_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and _60646_ (_15559_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor _60647_ (_15560_, _15559_, _15558_);
  and _60648_ (_15561_, _15560_, _15557_);
  and _60649_ (_15562_, _15561_, _15553_);
  nor _60650_ (_15563_, _15562_, _33140_);
  nor _60651_ (_15564_, _15563_, _15550_);
  nor _60652_ (_15565_, _15564_, _34325_);
  nor _60653_ (_15566_, _15565_, _15549_);
  nor _60654_ (_36866_[5], _15566_, rst);
  and _60655_ (_15567_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and _60656_ (_15568_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and _60657_ (_15569_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _60658_ (_15570_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _60659_ (_15571_, _15570_, _15569_);
  and _60660_ (_15572_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _60661_ (_15573_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _60662_ (_15574_, _15573_, _15572_);
  and _60663_ (_15575_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  not _60664_ (_15576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _60665_ (_15577_, _33146_, _15576_);
  nor _60666_ (_15578_, _15577_, _15575_);
  and _60667_ (_15579_, _15578_, _15574_);
  and _60668_ (_15580_, _15579_, _15571_);
  nor _60669_ (_15581_, _15580_, _33140_);
  nor _60670_ (_15582_, _15581_, _15568_);
  nor _60671_ (_15583_, _15582_, _34325_);
  nor _60672_ (_15584_, _15583_, _15567_);
  nor _60673_ (_36866_[6], _15584_, rst);
  and _60674_ (_15585_, _33136_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or _60675_ (_15586_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _60676_ (_15587_, _15585_, _14142_);
  and _60677_ (_15588_, _15587_, _38997_);
  and _60678_ (_36889_[15], _15588_, _15586_);
  not _60679_ (_15589_, _15585_);
  or _60680_ (_15590_, _15589_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _60681_ (_00006_, _15585_, _38997_);
  and _60682_ (_15591_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _38997_);
  or _60683_ (_15592_, _15591_, _00006_);
  and _60684_ (_36890_[15], _15592_, _15590_);
  and _60685_ (_36891_, _34346_, _38997_);
  nor _60686_ (_36892_[4], _34239_, rst);
  and _60687_ (_36893_[7], _34320_, _38997_);
  nor _60688_ (_15593_, _34529_, _34227_);
  and _60689_ (_15594_, _34529_, _34227_);
  nor _60690_ (_15595_, _15594_, _15593_);
  nor _60691_ (_15596_, _34637_, _34232_);
  and _60692_ (_15597_, _34637_, _34232_);
  nor _60693_ (_15598_, _15597_, _15596_);
  and _60694_ (_15599_, _15598_, _15595_);
  nor _60695_ (_15600_, _34421_, _34251_);
  and _60696_ (_15601_, _34421_, _34251_);
  nor _60697_ (_15602_, _15601_, _15600_);
  nor _60698_ (_15603_, _34691_, _33631_);
  and _60699_ (_15604_, _34691_, _33631_);
  nor _60700_ (_15605_, _15604_, _15603_);
  and _60701_ (_15606_, _15605_, _34710_);
  and _60702_ (_15607_, _15606_, _15602_);
  and _60703_ (_15608_, _15607_, _15599_);
  and _60704_ (_15609_, _34579_, _11341_);
  nor _60705_ (_15610_, _34579_, _11341_);
  or _60706_ (_15611_, _15610_, _15609_);
  nor _60707_ (_15612_, _34471_, _33558_);
  and _60708_ (_15613_, _34471_, _33558_);
  nor _60709_ (_15614_, _15613_, _15612_);
  nor _60710_ (_15615_, _15614_, _15611_);
  nor _60711_ (_15616_, _34770_, _33644_);
  and _60712_ (_15617_, _34770_, _33644_);
  nor _60713_ (_15618_, _15617_, _15616_);
  nor _60714_ (_15619_, _15618_, _13118_);
  and _60715_ (_15620_, _15619_, _15615_);
  and _60716_ (_15621_, _15620_, _15608_);
  nor _60717_ (_15622_, _33618_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _60718_ (_15623_, _15622_, _15621_);
  not _60719_ (_15624_, _15623_);
  not _60720_ (_15625_, _33462_);
  and _60721_ (_15626_, _15625_, _33362_);
  nor _60722_ (_15627_, _15626_, _33467_);
  and _60723_ (_15628_, _15627_, _15625_);
  nor _60724_ (_15629_, _11075_, _11089_);
  and _60725_ (_15630_, _15629_, _15608_);
  and _60726_ (_15631_, _15630_, _15628_);
  not _60727_ (_15632_, _15631_);
  nor _60728_ (_15633_, _15022_, _33275_);
  not _60729_ (_15634_, _33361_);
  not _60730_ (_15635_, _14089_);
  not _60731_ (_15636_, _15627_);
  and _60732_ (_15637_, _15636_, _33463_);
  nor _60733_ (_15638_, _14206_, _35617_);
  and _60734_ (_15639_, _15638_, _14335_);
  and _60735_ (_15640_, _15639_, _14401_);
  not _60736_ (_15641_, _15640_);
  nor _60737_ (_15642_, _15641_, _14469_);
  and _60738_ (_15643_, _15642_, _14542_);
  and _60739_ (_15644_, _15643_, _14616_);
  and _60740_ (_15645_, _15644_, _15637_);
  and _60741_ (_15646_, _15645_, _15635_);
  not _60742_ (_15647_, _15646_);
  and _60743_ (_15648_, _15628_, _33728_);
  nor _60744_ (_15649_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _60745_ (_15650_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _60746_ (_15651_, _15650_, _15649_);
  nor _60747_ (_15652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _60748_ (_15653_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _60749_ (_15654_, _15653_, _15652_);
  and _60750_ (_15655_, _15654_, _15651_);
  and _60751_ (_15656_, _15655_, _33460_);
  and _60752_ (_15657_, _33462_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _60753_ (_15658_, _15657_, _15656_);
  nor _60754_ (_15659_, _15658_, _15648_);
  and _60755_ (_15660_, _15659_, _15647_);
  or _60756_ (_15661_, _15660_, _15634_);
  nor _60757_ (_15662_, _15661_, _15633_);
  or _60758_ (_15663_, _33382_, _33408_);
  and _60759_ (_15664_, _15663_, _33252_);
  not _60760_ (_15665_, _15664_);
  and _60761_ (_15666_, _15063_, _33353_);
  and _60762_ (_15667_, _15666_, _15665_);
  not _60763_ (_15668_, _15093_);
  nor _60764_ (_15669_, _15291_, _33419_);
  and _60765_ (_15670_, _15669_, _15668_);
  and _60766_ (_15671_, _15670_, _15667_);
  and _60767_ (_15672_, _15671_, _15660_);
  nor _60768_ (_15673_, _15672_, _15662_);
  nor _60769_ (_15674_, _15029_, _15335_);
  and _60770_ (_15675_, _15674_, _33510_);
  not _60771_ (_15676_, _15675_);
  nor _60772_ (_15677_, _15676_, _15673_);
  nor _60773_ (_15678_, _15677_, _34367_);
  not _60774_ (_15679_, _15678_);
  nor _60775_ (_15680_, _15079_, _33477_);
  nor _60776_ (_15681_, _15680_, _33469_);
  and _60777_ (_15682_, _15681_, _15679_);
  and _60778_ (_15683_, _14820_, _14836_);
  not _60779_ (_15684_, _15683_);
  and _60780_ (_15685_, _15684_, _33460_);
  not _60781_ (_15686_, _13512_);
  nor _60782_ (_15687_, _13518_, _34235_);
  and _60783_ (_15688_, _15687_, _15686_);
  not _60784_ (_15689_, _15688_);
  and _60785_ (_15690_, _15689_, _33462_);
  nor _60786_ (_15691_, _15690_, _15685_);
  not _60787_ (_15692_, _15691_);
  nor _60788_ (_15693_, _15692_, _15682_);
  and _60789_ (_15694_, _15693_, _15632_);
  and _60790_ (_15695_, _15694_, _15624_);
  and _60791_ (_15696_, _15695_, _33470_);
  and _60792_ (_36896_, _15696_, _38997_);
  and _60793_ (_36897_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _38997_);
  and _60794_ (_36898_[7], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _38997_);
  nor _60795_ (_15697_, _33161_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _60796_ (_15698_, _15697_, _34325_);
  nor _60797_ (_15699_, _15698_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not _60798_ (_15700_, _15699_);
  and _60799_ (_15701_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _60800_ (_15702_, _15701_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _60801_ (_15703_, _15702_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _60802_ (_15704_, _15703_, _15700_);
  and _60803_ (_15705_, _15704_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _60804_ (_15706_, _15705_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _60805_ (_15707_, _15706_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _60806_ (_15708_, _15707_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _60807_ (_15709_, _15708_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _60808_ (_15710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _60809_ (_15711_, _15710_, _15709_);
  and _60810_ (_15712_, _15711_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _60811_ (_15713_, _15712_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _60812_ (_15714_, _15713_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand _60813_ (_15715_, _15713_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _60814_ (_15716_, _15715_, _15714_);
  or _60815_ (_15717_, _15716_, _15695_);
  and _60816_ (_15718_, _15717_, _38997_);
  and _60817_ (_15719_, _15063_, _33362_);
  nand _60818_ (_15720_, _15719_, _15669_);
  nand _60819_ (_15721_, _15720_, _33458_);
  and _60820_ (_15722_, _33358_, _33465_);
  nand _60821_ (_15723_, _15722_, _33131_);
  and _60822_ (_15724_, _33350_, _33131_);
  and _60823_ (_15725_, _15724_, _33252_);
  nor _60824_ (_15726_, _15725_, _33469_);
  and _60825_ (_15727_, _15726_, _15723_);
  and _60826_ (_15728_, _15727_, _15721_);
  and _60827_ (_15729_, _15728_, _34342_);
  nand _60828_ (_15730_, _15727_, _15721_);
  and _60829_ (_15731_, _15730_, _15459_);
  nor _60830_ (_15732_, _15731_, _15729_);
  and _60831_ (_15733_, _15732_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _60832_ (_15734_, _15732_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _60833_ (_15735_, _15734_);
  and _60834_ (_15736_, _15728_, _34685_);
  and _60835_ (_15737_, _15730_, _15584_);
  nor _60836_ (_15738_, _15737_, _15736_);
  and _60837_ (_15739_, _15738_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not _60838_ (_15740_, _15739_);
  nor _60839_ (_15741_, _15738_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _60840_ (_15742_, _15741_, _15739_);
  and _60841_ (_15743_, _15728_, _34603_);
  and _60842_ (_15744_, _15730_, _15566_);
  nor _60843_ (_15745_, _15744_, _15743_);
  nor _60844_ (_15746_, _15745_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _60845_ (_15747_, _15745_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _60846_ (_15748_, _15728_, _34495_);
  and _60847_ (_15749_, _15730_, _15548_);
  nor _60848_ (_15750_, _15749_, _15748_);
  nand _60849_ (_15751_, _15750_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _60850_ (_15752_, _15728_, _34417_);
  and _60851_ (_15753_, _15730_, _15530_);
  nor _60852_ (_15754_, _15753_, _15752_);
  nor _60853_ (_15755_, _15754_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _60854_ (_15756_, _15754_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _60855_ (_15757_, _34757_);
  or _60856_ (_15758_, _15730_, _15757_);
  not _60857_ (_15759_, _15512_);
  or _60858_ (_15760_, _15728_, _15759_);
  and _60859_ (_15761_, _15760_, _15758_);
  and _60860_ (_15762_, _15761_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _60861_ (_15763_, _34575_);
  or _60862_ (_15764_, _15730_, _15763_);
  not _60863_ (_15765_, _15494_);
  or _60864_ (_15766_, _15728_, _15765_);
  and _60865_ (_15767_, _15766_, _15764_);
  nand _60866_ (_15768_, _15767_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _60867_ (_15769_, _15768_);
  not _60868_ (_15770_, _34457_);
  or _60869_ (_15771_, _15730_, _15770_);
  not _60870_ (_15772_, _15477_);
  or _60871_ (_15773_, _15728_, _15772_);
  and _60872_ (_15774_, _15773_, _15771_);
  and _60873_ (_15775_, _15774_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _60874_ (_15776_, _15767_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _60875_ (_15777_, _15776_, _15768_);
  and _60876_ (_15778_, _15777_, _15775_);
  or _60877_ (_15779_, _15778_, _15769_);
  not _60878_ (_15780_, _15762_);
  or _60879_ (_15781_, _15761_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _60880_ (_15782_, _15781_, _15780_);
  and _60881_ (_15783_, _15782_, _15779_);
  or _60882_ (_15784_, _15783_, _15762_);
  nor _60883_ (_15785_, _15784_, _15756_);
  nor _60884_ (_15786_, _15785_, _15755_);
  or _60885_ (_15787_, _15750_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _60886_ (_15788_, _15787_, _15751_);
  nand _60887_ (_15789_, _15788_, _15786_);
  nand _60888_ (_15790_, _15789_, _15751_);
  nor _60889_ (_15791_, _15790_, _15747_);
  nor _60890_ (_15792_, _15791_, _15746_);
  nand _60891_ (_15793_, _15792_, _15742_);
  nand _60892_ (_15794_, _15793_, _15740_);
  and _60893_ (_15795_, _15794_, _15735_);
  or _60894_ (_15796_, _15795_, _15733_);
  and _60895_ (_15797_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _60896_ (_15798_, _15797_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _60897_ (_15799_, _15798_, _15796_);
  and _60898_ (_15800_, _15799_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _60899_ (_15801_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _60900_ (_15802_, _15801_, _15800_);
  or _60901_ (_15803_, _15802_, _15732_);
  not _60902_ (_15804_, _15732_);
  or _60903_ (_15805_, _15796_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _60904_ (_15806_, _15805_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _60905_ (_15807_, _15806_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _60906_ (_15808_, _15807_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _60907_ (_15809_, _15808_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _60908_ (_15810_, _15809_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _60909_ (_15811_, _15810_, _15804_);
  nand _60910_ (_15812_, _15811_, _15803_);
  nor _60911_ (_15813_, _15732_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _60912_ (_15814_, _15732_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _60913_ (_15815_, _15814_, _15813_);
  or _60914_ (_15816_, _15815_, _15812_);
  nor _60915_ (_15817_, _15816_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _60916_ (_15818_, _15816_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or _60917_ (_15819_, _15818_, _15817_);
  and _60918_ (_15820_, _15063_, _15022_);
  and _60919_ (_15821_, _15820_, _33362_);
  and _60920_ (_15822_, _15821_, _15674_);
  and _60921_ (_15823_, _15822_, _15670_);
  nor _60922_ (_15824_, _15823_, _34367_);
  nor _60923_ (_15825_, _15824_, _15725_);
  nor _60924_ (_15826_, _33484_, _34367_);
  nor _60925_ (_15827_, _15826_, _15680_);
  not _60926_ (_15828_, _15827_);
  and _60927_ (_15829_, _15828_, _15728_);
  nor _60928_ (_15830_, _15829_, _15825_);
  and _60929_ (_15831_, _15830_, _15819_);
  nor _60930_ (_15832_, _14098_, _33470_);
  not _60931_ (_15833_, _15826_);
  nor _60932_ (_15834_, _15833_, _14189_);
  not _60933_ (_15835_, _34342_);
  and _60934_ (_15836_, _15828_, _15730_);
  and _60935_ (_15837_, _15836_, _15835_);
  and _60936_ (_15838_, _33252_, _33131_);
  and _60937_ (_15839_, _15838_, _33350_);
  not _60938_ (_15840_, _15839_);
  not _60939_ (_15841_, _33468_);
  nor _60940_ (_15842_, _15841_, _33442_);
  and _60941_ (_15843_, _15078_, _33131_);
  nor _60942_ (_15844_, _15843_, _15842_);
  and _60943_ (_15845_, _15844_, _15721_);
  and _60944_ (_15846_, _15845_, _15840_);
  nor _60945_ (_15847_, _15828_, _15824_);
  and _60946_ (_15848_, _15847_, _15846_);
  and _60947_ (_15849_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _60948_ (_15850_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _60949_ (_15851_, _15850_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _60950_ (_15852_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _60951_ (_15853_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _60952_ (_15854_, _15853_, _15852_);
  and _60953_ (_15855_, _15854_, _15851_);
  and _60954_ (_15856_, _15855_, _15798_);
  and _60955_ (_15857_, _15856_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _60956_ (_15858_, _15857_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _60957_ (_15859_, _15858_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _60958_ (_15860_, _15859_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _60959_ (_15861_, _15860_, _14142_);
  or _60960_ (_15862_, _15860_, _14142_);
  and _60961_ (_15863_, _15862_, _15861_);
  not _60962_ (_15864_, _15824_);
  and _60963_ (_15865_, _15829_, _15864_);
  and _60964_ (_15866_, _15865_, _15863_);
  or _60965_ (_15867_, _15866_, _15849_);
  or _60966_ (_15868_, _15867_, _15837_);
  nor _60967_ (_15869_, _15868_, _15834_);
  nand _60968_ (_15870_, _15869_, _15695_);
  or _60969_ (_15871_, _15870_, _15832_);
  or _60970_ (_15872_, _15871_, _15831_);
  and _60971_ (_36899_[15], _15872_, _15718_);
  and _60972_ (_15873_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _38997_);
  and _60973_ (_15874_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _60974_ (_15875_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _60975_ (_15876_, _33135_, _15875_);
  not _60976_ (_15877_, _15876_);
  not _60977_ (_15878_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _60978_ (_15879_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _60979_ (_15880_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _60980_ (_15881_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _60981_ (_15882_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _60982_ (_15883_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _60983_ (_15884_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _60984_ (_15885_, _15884_, _15882_);
  and _60985_ (_15886_, _15885_, _15883_);
  nor _60986_ (_15887_, _15886_, _15882_);
  nor _60987_ (_15888_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _60988_ (_15889_, _15888_, _15881_);
  not _60989_ (_15890_, _15889_);
  nor _60990_ (_15891_, _15890_, _15887_);
  nor _60991_ (_15892_, _15891_, _15881_);
  not _60992_ (_15893_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _60993_ (_15894_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not _60994_ (_15895_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _60995_ (_15896_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not _60996_ (_15897_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _60997_ (_15898_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _60998_ (_15899_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _60999_ (_15900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _61000_ (_15901_, _15900_, _15899_);
  and _61001_ (_15902_, _15901_, _15898_);
  and _61002_ (_15903_, _15902_, _15897_);
  and _61003_ (_15904_, _15903_, _15896_);
  and _61004_ (_15905_, _15904_, _15895_);
  and _61005_ (_15906_, _15905_, _15894_);
  and _61006_ (_15907_, _15906_, _15893_);
  and _61007_ (_15908_, _15907_, _15892_);
  and _61008_ (_15909_, _15908_, _15880_);
  and _61009_ (_15910_, _15909_, _15879_);
  and _61010_ (_15911_, _15910_, _15878_);
  nor _61011_ (_15912_, _15911_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _61012_ (_15913_, _15911_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _61013_ (_15914_, _15913_, _15912_);
  nor _61014_ (_15915_, _15910_, _15878_);
  nor _61015_ (_15916_, _15915_, _15911_);
  not _61016_ (_15917_, _15916_);
  nor _61017_ (_15918_, _15909_, _15879_);
  nor _61018_ (_15919_, _15918_, _15910_);
  not _61019_ (_15920_, _15919_);
  nor _61020_ (_15921_, _15908_, _15880_);
  nor _61021_ (_15922_, _15921_, _15909_);
  not _61022_ (_15923_, _15922_);
  and _61023_ (_15924_, _15892_, _15906_);
  nor _61024_ (_15925_, _15924_, _15893_);
  nor _61025_ (_15926_, _15925_, _15908_);
  not _61026_ (_15927_, _15926_);
  and _61027_ (_15928_, _15892_, _15904_);
  and _61028_ (_15929_, _15928_, _15895_);
  nor _61029_ (_15930_, _15929_, _15894_);
  or _61030_ (_15931_, _15930_, _15924_);
  nor _61031_ (_15932_, _15928_, _15895_);
  nor _61032_ (_15933_, _15932_, _15929_);
  not _61033_ (_15934_, _15933_);
  and _61034_ (_15935_, _15892_, _15902_);
  nor _61035_ (_15936_, _15935_, _15897_);
  and _61036_ (_15937_, _15892_, _15903_);
  nor _61037_ (_15938_, _15937_, _15936_);
  not _61038_ (_15939_, _15938_);
  and _61039_ (_15940_, _15892_, _15901_);
  nor _61040_ (_15941_, _15940_, _15898_);
  nor _61041_ (_15942_, _15941_, _15935_);
  not _61042_ (_15943_, _15942_);
  and _61043_ (_15944_, _15892_, _15900_);
  nor _61044_ (_15945_, _15944_, _15899_);
  nor _61045_ (_15946_, _15945_, _15940_);
  not _61046_ (_15947_, _15946_);
  not _61047_ (_15948_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _61048_ (_15949_, _15892_, _15948_);
  nor _61049_ (_15950_, _15892_, _15948_);
  nor _61050_ (_15951_, _15950_, _15949_);
  not _61051_ (_15952_, _15951_);
  not _61052_ (_15953_, _14966_);
  and _61053_ (_15954_, _14962_, _14932_);
  not _61054_ (_15955_, _15954_);
  and _61055_ (_15956_, _14954_, _14974_);
  nor _61056_ (_15957_, _15956_, _14980_);
  and _61057_ (_15958_, _15957_, _15955_);
  and _61058_ (_15959_, _14976_, _14943_);
  and _61059_ (_15960_, _14943_, _14974_);
  or _61060_ (_15961_, _15960_, _15959_);
  not _61061_ (_15962_, _15961_);
  nor _61062_ (_15963_, _14996_, _14945_);
  and _61063_ (_15964_, _15963_, _15962_);
  and _61064_ (_15965_, _15964_, _15958_);
  nor _61065_ (_15966_, _15965_, _15953_);
  not _61066_ (_15967_, _15966_);
  not _61067_ (_15968_, _14967_);
  and _61068_ (_15969_, _14959_, _14944_);
  nor _61069_ (_15970_, _15969_, _14981_);
  nor _61070_ (_15971_, _15970_, _15968_);
  not _61071_ (_15972_, _15971_);
  and _61072_ (_15973_, _15972_, _14995_);
  and _61073_ (_15974_, _15973_, _15967_);
  and _61074_ (_15975_, _15960_, _14929_);
  and _61075_ (_15976_, _14966_, _14963_);
  nor _61076_ (_15977_, _15976_, _15975_);
  nor _61077_ (_15978_, _14965_, _14942_);
  not _61078_ (_15979_, _15978_);
  and _61079_ (_15980_, _15979_, _14986_);
  and _61080_ (_15981_, _14976_, _14932_);
  and _61081_ (_15982_, _15981_, _14981_);
  nor _61082_ (_15983_, _15982_, _15980_);
  and _61083_ (_15984_, _15983_, _15977_);
  and _61084_ (_15985_, _14954_, _14930_);
  and _61085_ (_15986_, _15985_, _14951_);
  not _61086_ (_15987_, _15986_);
  and _61087_ (_15988_, _33246_, _14935_);
  and _61088_ (_15989_, _15988_, _14943_);
  and _61089_ (_15990_, _15989_, _14941_);
  nor _61090_ (_15991_, _15990_, _14938_);
  and _61091_ (_15992_, _15991_, _15987_);
  not _61092_ (_15993_, _33197_);
  and _61093_ (_15994_, _14963_, _15993_);
  and _61094_ (_15995_, _15956_, _14942_);
  nor _61095_ (_15996_, _15995_, _15994_);
  and _61096_ (_15997_, _15996_, _15992_);
  and _61097_ (_15998_, _15997_, _14957_);
  and _61098_ (_15999_, _15998_, _15984_);
  and _61099_ (_16000_, _14990_, _33222_);
  and _61100_ (_16001_, _16000_, _15979_);
  not _61101_ (_16002_, _16001_);
  and _61102_ (_16003_, _14997_, _14990_);
  not _61103_ (_16004_, _14959_);
  nor _61104_ (_16005_, _15960_, _14996_);
  nor _61105_ (_16006_, _16005_, _16004_);
  nor _61106_ (_16007_, _16006_, _16003_);
  and _61107_ (_16008_, _16007_, _16002_);
  and _61108_ (_16009_, _14945_, _14929_);
  nor _61109_ (_16010_, _15959_, _14996_);
  nor _61110_ (_16011_, _16010_, _33197_);
  nor _61111_ (_16012_, _16011_, _16009_);
  nor _61112_ (_16013_, _15959_, _14937_);
  not _61113_ (_16014_, _16013_);
  and _61114_ (_16015_, _16014_, _14929_);
  or _61115_ (_16016_, _14963_, _14996_);
  and _61116_ (_16017_, _16016_, _14981_);
  nor _61117_ (_16018_, _16017_, _16015_);
  and _61118_ (_16019_, _16018_, _16012_);
  and _61119_ (_16020_, _16019_, _16008_);
  and _61120_ (_16021_, _16020_, _15999_);
  and _61121_ (_16022_, _14981_, _14945_);
  and _61122_ (_16023_, _14997_, _15956_);
  nor _61123_ (_16024_, _16023_, _16022_);
  and _61124_ (_16025_, _14959_, _14945_);
  not _61125_ (_16026_, _16025_);
  and _61126_ (_16027_, _16026_, _14983_);
  and _61127_ (_16028_, _16027_, _16024_);
  not _61128_ (_16029_, _14981_);
  nor _61129_ (_16030_, _15954_, _15960_);
  and _61130_ (_16031_, _14944_, _14932_);
  nor _61131_ (_16032_, _16031_, _14990_);
  and _61132_ (_16033_, _16032_, _16030_);
  nor _61133_ (_16034_, _16033_, _16029_);
  not _61134_ (_16035_, _16034_);
  and _61135_ (_16036_, _14977_, _14959_);
  nor _61136_ (_16037_, _16036_, _14971_);
  and _61137_ (_16038_, _16037_, _16035_);
  and _61138_ (_16039_, _16038_, _16028_);
  and _61139_ (_16040_, _16039_, _16021_);
  and _61140_ (_16041_, _16040_, _15974_);
  nor _61141_ (_16042_, _15885_, _15883_);
  nor _61142_ (_16043_, _16042_, _15886_);
  not _61143_ (_16044_, _16043_);
  nor _61144_ (_16045_, _16044_, _16041_);
  not _61145_ (_16046_, _16045_);
  and _61146_ (_16047_, _14997_, _14986_);
  or _61147_ (_16048_, _16003_, _16047_);
  or _61148_ (_16049_, _16017_, _15975_);
  or _61149_ (_16050_, _14993_, _14969_);
  or _61150_ (_16051_, _16050_, _16049_);
  or _61151_ (_16052_, _16051_, _16048_);
  not _61152_ (_16053_, _14953_);
  nand _61153_ (_16054_, _16028_, _16053_);
  or _61154_ (_16055_, _16054_, _16052_);
  nor _61155_ (_16056_, _16055_, _16041_);
  not _61156_ (_16057_, _16056_);
  nor _61157_ (_16058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _61158_ (_16059_, _16058_, _15883_);
  and _61159_ (_16060_, _16059_, _16057_);
  and _61160_ (_16061_, _16044_, _16041_);
  nor _61161_ (_16062_, _16061_, _16045_);
  nand _61162_ (_16063_, _16062_, _16060_);
  and _61163_ (_16064_, _16063_, _16046_);
  not _61164_ (_16065_, _16064_);
  and _61165_ (_16066_, _15890_, _15887_);
  nor _61166_ (_16067_, _16066_, _15891_);
  and _61167_ (_16068_, _16067_, _16065_);
  and _61168_ (_16069_, _16068_, _15952_);
  not _61169_ (_16070_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _61170_ (_16071_, _15949_, _16070_);
  or _61171_ (_16072_, _16071_, _15944_);
  and _61172_ (_16073_, _16072_, _16069_);
  and _61173_ (_16074_, _16073_, _15947_);
  and _61174_ (_16075_, _16074_, _15943_);
  and _61175_ (_16076_, _16075_, _15939_);
  nor _61176_ (_16077_, _15937_, _15896_);
  or _61177_ (_16078_, _16077_, _15928_);
  and _61178_ (_16079_, _16078_, _16076_);
  and _61179_ (_16080_, _16079_, _15934_);
  and _61180_ (_16081_, _16080_, _15931_);
  and _61181_ (_16082_, _16081_, _15927_);
  and _61182_ (_16083_, _16082_, _15923_);
  and _61183_ (_16084_, _16083_, _15920_);
  and _61184_ (_16085_, _16084_, _15917_);
  or _61185_ (_16086_, _16085_, _15914_);
  nand _61186_ (_16087_, _16085_, _15914_);
  and _61187_ (_16088_, _16087_, _16086_);
  or _61188_ (_16089_, _16088_, _15877_);
  or _61189_ (_16090_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _61190_ (_16091_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and _61191_ (_16092_, _16091_, _16090_);
  and _61192_ (_16093_, _16092_, _16089_);
  or _61193_ (_36900_[15], _16093_, _15874_);
  nor _61194_ (_16094_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _61195_ (_36901_, _16094_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _61196_ (_36902_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _38997_);
  not _61197_ (_16095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor _61198_ (_16096_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _61199_ (_16097_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _61200_ (_16098_, _16097_, _16096_);
  not _61201_ (_16099_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor _61202_ (_16100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _61203_ (_16101_, _16100_, _16099_);
  and _61204_ (_16102_, _16101_, _16098_);
  and _61205_ (_16103_, _16102_, _16095_);
  and _61206_ (_16104_, \oc8051_top_1.oc8051_rom1.ea_int , _33132_);
  nand _61207_ (_16105_, _16104_, _33135_);
  nand _61208_ (_16106_, _16105_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _61209_ (_16107_, _16106_, _16103_);
  and _61210_ (_36903_, _16107_, _38997_);
  and _61211_ (_16108_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _61212_ (_16109_, _16108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _61213_ (_36904_[7], _16109_, _38997_);
  nor _61214_ (_16110_, _15699_, _34325_);
  nor _61215_ (_16111_, _16041_, _33148_);
  not _61216_ (_16112_, _16111_);
  nor _61217_ (_16113_, _16056_, _33144_);
  and _61218_ (_16114_, _16041_, _33148_);
  nor _61219_ (_16115_, _16114_, _16111_);
  nand _61220_ (_16116_, _16115_, _16113_);
  and _61221_ (_16117_, _16116_, _16112_);
  nor _61222_ (_16118_, _16117_, _34325_);
  and _61223_ (_16119_, _16118_, _33143_);
  nor _61224_ (_16120_, _16118_, _33143_);
  nor _61225_ (_16121_, _16120_, _16119_);
  nor _61226_ (_16122_, _16121_, _16110_);
  and _61227_ (_16123_, _33149_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _61228_ (_16124_, _16123_, _16110_);
  and _61229_ (_16125_, _16124_, _16055_);
  or _61230_ (_16126_, _16125_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _61231_ (_16127_, _16126_, _16122_);
  and _61232_ (_36905_[2], _16127_, _38997_);
  and _61233_ (_16128_, _33240_, _33265_);
  and _61234_ (_16129_, _33338_, _33313_);
  and _61235_ (_16130_, _16129_, _16128_);
  and _61236_ (_16131_, _33136_, _38997_);
  and _61237_ (_16132_, _16131_, _33191_);
  and _61238_ (_16133_, _16132_, _33217_);
  and _61239_ (_16134_, _33167_, _33290_);
  and _61240_ (_16135_, _16134_, _16133_);
  and _61241_ (_36908_, _16135_, _16130_);
  nor _61242_ (_16136_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and _61243_ (_16137_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _61244_ (_16138_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and _61245_ (_36910_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _38997_);
  and _61246_ (_16139_, _36910_, _16138_);
  or _61247_ (_36909_[7], _16139_, _16137_);
  not _61248_ (_16140_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _61249_ (_16141_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _61250_ (_16142_, _16141_, _16140_);
  and _61251_ (_16143_, _16141_, _16140_);
  nor _61252_ (_16144_, _16143_, _16142_);
  not _61253_ (_16145_, _16144_);
  and _61254_ (_16146_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _61255_ (_16147_, _16146_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _61256_ (_16148_, _16146_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _61257_ (_16149_, _16148_, _16147_);
  or _61258_ (_16150_, _16149_, _16141_);
  and _61259_ (_16151_, _16150_, _16145_);
  nor _61260_ (_16152_, _16142_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _61261_ (_16153_, _16142_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _61262_ (_16154_, _16153_, _16152_);
  or _61263_ (_16155_, _16147_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _61264_ (_36912_[3], _16155_, _38997_);
  and _61265_ (_16156_, _36912_[3], _16154_);
  and _61266_ (_36911_, _16156_, _16151_);
  not _61267_ (_16157_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor _61268_ (_16158_, _15699_, _16157_);
  and _61269_ (_16159_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not _61270_ (_16160_, _16158_);
  and _61271_ (_16161_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or _61272_ (_16162_, _16161_, _16159_);
  and _61273_ (_36913_[31], _16162_, _38997_);
  and _61274_ (_16163_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor _61275_ (_16164_, _16158_, _34334_);
  or _61276_ (_16165_, _16164_, _16163_);
  and _61277_ (_36914_[31], _16165_, _38997_);
  and _61278_ (_16166_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not _61279_ (_16167_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _61280_ (_16168_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _16167_);
  and _61281_ (_16169_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _61282_ (_16170_, _16169_, _16166_);
  and _61283_ (_36915_[7], _16170_, _38997_);
  and _61284_ (_16171_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  or _61285_ (_16172_, _16171_, _16168_);
  and _61286_ (_36916_, _16172_, _38997_);
  or _61287_ (_16173_, _16167_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and _61288_ (_36917_, _16173_, _38997_);
  not _61289_ (_16174_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _61290_ (_16175_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _61291_ (_16176_, _16175_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _61292_ (_16177_, _16167_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and _61293_ (_16178_, _16177_, _38997_);
  and _61294_ (_36918_[15], _16178_, _16176_);
  or _61295_ (_16179_, _16167_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _61296_ (_36919_, _16179_, _38997_);
  nor _61297_ (_16180_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _61298_ (_16181_, _16180_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _61299_ (_16182_, _16181_, _38997_);
  and _61300_ (_16183_, _36910_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _61301_ (_36920_, _16183_, _16182_);
  and _61302_ (_16184_, _16157_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _61303_ (_16185_, _16184_, _16181_);
  and _61304_ (_36921_, _16185_, _38997_);
  nand _61305_ (_16186_, _16181_, _14189_);
  or _61306_ (_16187_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and _61307_ (_16188_, _16187_, _38997_);
  and _61308_ (_36922_[15], _16188_, _16186_);
  and _61309_ (_16189_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _61310_ (_16190_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _61311_ (_16191_, _15585_, _16190_);
  or _61312_ (_16192_, _16191_, _16189_);
  and _61313_ (_36889_[0], _16192_, _38997_);
  and _61314_ (_16193_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _61315_ (_16194_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _61316_ (_16195_, _15585_, _16194_);
  or _61317_ (_16196_, _16195_, _16193_);
  and _61318_ (_36889_[1], _16196_, _38997_);
  and _61319_ (_16197_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _61320_ (_16198_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _61321_ (_16199_, _15585_, _16198_);
  or _61322_ (_16200_, _16199_, _16197_);
  and _61323_ (_36889_[2], _16200_, _38997_);
  and _61324_ (_16201_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _61325_ (_16202_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _61326_ (_16203_, _15585_, _16202_);
  or _61327_ (_16204_, _16203_, _16201_);
  and _61328_ (_36889_[3], _16204_, _38997_);
  and _61329_ (_16205_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not _61330_ (_16206_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _61331_ (_16207_, _15585_, _16206_);
  or _61332_ (_16208_, _16207_, _16205_);
  and _61333_ (_36889_[4], _16208_, _38997_);
  and _61334_ (_16209_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not _61335_ (_16210_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _61336_ (_16211_, _15585_, _16210_);
  or _61337_ (_16212_, _16211_, _16209_);
  and _61338_ (_36889_[5], _16212_, _38997_);
  and _61339_ (_16213_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not _61340_ (_16214_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _61341_ (_16215_, _15585_, _16214_);
  or _61342_ (_16216_, _16215_, _16213_);
  and _61343_ (_36889_[6], _16216_, _38997_);
  and _61344_ (_16217_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _61345_ (_16218_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _61346_ (_16219_, _15585_, _16218_);
  or _61347_ (_16220_, _16219_, _16217_);
  and _61348_ (_36889_[7], _16220_, _38997_);
  and _61349_ (_16221_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not _61350_ (_16222_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _61351_ (_16223_, _15585_, _16222_);
  or _61352_ (_16224_, _16223_, _16221_);
  and _61353_ (_36889_[8], _16224_, _38997_);
  and _61354_ (_16225_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not _61355_ (_16226_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _61356_ (_16227_, _15585_, _16226_);
  or _61357_ (_16228_, _16227_, _16225_);
  and _61358_ (_36889_[9], _16228_, _38997_);
  and _61359_ (_16229_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not _61360_ (_16230_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _61361_ (_16231_, _15585_, _16230_);
  or _61362_ (_16232_, _16231_, _16229_);
  and _61363_ (_36889_[10], _16232_, _38997_);
  and _61364_ (_16233_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not _61365_ (_16234_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _61366_ (_16235_, _15585_, _16234_);
  or _61367_ (_16236_, _16235_, _16233_);
  and _61368_ (_36889_[11], _16236_, _38997_);
  and _61369_ (_16237_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not _61370_ (_16238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor _61371_ (_16239_, _15585_, _16238_);
  or _61372_ (_16240_, _16239_, _16237_);
  and _61373_ (_36889_[12], _16240_, _38997_);
  and _61374_ (_16241_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not _61375_ (_16242_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _61376_ (_16243_, _15585_, _16242_);
  or _61377_ (_16244_, _16243_, _16241_);
  and _61378_ (_36889_[13], _16244_, _38997_);
  and _61379_ (_16245_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not _61380_ (_16246_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _61381_ (_16247_, _15585_, _16246_);
  or _61382_ (_16248_, _16247_, _16245_);
  and _61383_ (_36889_[14], _16248_, _38997_);
  or _61384_ (_16249_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand _61385_ (_16250_, _15585_, _16190_);
  and _61386_ (_16251_, _16250_, _38997_);
  and _61387_ (_36890_[0], _16251_, _16249_);
  or _61388_ (_16252_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nand _61389_ (_16253_, _15585_, _16194_);
  and _61390_ (_16254_, _16253_, _38997_);
  and _61391_ (_36890_[1], _16254_, _16252_);
  or _61392_ (_16255_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nand _61393_ (_16256_, _15585_, _16198_);
  and _61394_ (_16257_, _16256_, _38997_);
  and _61395_ (_36890_[2], _16257_, _16255_);
  or _61396_ (_16258_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nand _61397_ (_16259_, _15585_, _16202_);
  and _61398_ (_16260_, _16259_, _38997_);
  and _61399_ (_36890_[3], _16260_, _16258_);
  or _61400_ (_16261_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nand _61401_ (_16262_, _15585_, _16206_);
  and _61402_ (_16263_, _16262_, _38997_);
  and _61403_ (_36890_[4], _16263_, _16261_);
  or _61404_ (_16264_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nand _61405_ (_16265_, _15585_, _16210_);
  and _61406_ (_16266_, _16265_, _38997_);
  and _61407_ (_36890_[5], _16266_, _16264_);
  or _61408_ (_16267_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nand _61409_ (_16268_, _15585_, _16214_);
  and _61410_ (_16269_, _16268_, _38997_);
  and _61411_ (_36890_[6], _16269_, _16267_);
  or _61412_ (_16270_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nand _61413_ (_16271_, _15585_, _16218_);
  and _61414_ (_16272_, _16271_, _38997_);
  and _61415_ (_36890_[7], _16272_, _16270_);
  or _61416_ (_16273_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nand _61417_ (_16274_, _15585_, _16222_);
  and _61418_ (_16275_, _16274_, _38997_);
  and _61419_ (_36890_[8], _16275_, _16273_);
  or _61420_ (_16276_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nand _61421_ (_16277_, _15585_, _16226_);
  and _61422_ (_16278_, _16277_, _38997_);
  and _61423_ (_36890_[9], _16278_, _16276_);
  or _61424_ (_16279_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nand _61425_ (_16280_, _15585_, _16230_);
  and _61426_ (_16281_, _16280_, _38997_);
  and _61427_ (_36890_[10], _16281_, _16279_);
  or _61428_ (_16282_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nand _61429_ (_16283_, _15585_, _16234_);
  and _61430_ (_16284_, _16283_, _38997_);
  and _61431_ (_36890_[11], _16284_, _16282_);
  or _61432_ (_16285_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nand _61433_ (_16286_, _15585_, _16238_);
  and _61434_ (_16287_, _16286_, _38997_);
  and _61435_ (_36890_[12], _16287_, _16285_);
  or _61436_ (_16288_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nand _61437_ (_16289_, _15585_, _16242_);
  and _61438_ (_16290_, _16289_, _38997_);
  and _61439_ (_36890_[13], _16290_, _16288_);
  or _61440_ (_16291_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nand _61441_ (_16292_, _15585_, _16246_);
  and _61442_ (_16293_, _16292_, _38997_);
  and _61443_ (_36890_[14], _16293_, _16291_);
  and _61444_ (_36892_[0], _33226_, _38997_);
  and _61445_ (_36892_[1], _33250_, _38997_);
  and _61446_ (_36892_[2], _33177_, _38997_);
  nor _61447_ (_36892_[3], _34283_, rst);
  nor _61448_ (_16294_, _16158_, _15469_);
  and _61449_ (_16295_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or _61450_ (_16296_, _16295_, _16294_);
  and _61451_ (_36913_[0], _16296_, _38997_);
  and _61452_ (_16297_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _61453_ (_16298_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and _61454_ (_16299_, _16298_, _16158_);
  or _61455_ (_16300_, _16299_, _16297_);
  and _61456_ (_36913_[1], _16300_, _38997_);
  nor _61457_ (_16301_, _16158_, _15501_);
  and _61458_ (_16302_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or _61459_ (_16303_, _16302_, _16301_);
  and _61460_ (_36913_[2], _16303_, _38997_);
  nor _61461_ (_16304_, _16158_, _15522_);
  and _61462_ (_16305_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and _61463_ (_16306_, _16305_, _16158_);
  or _61464_ (_16307_, _16306_, _16304_);
  and _61465_ (_36913_[3], _16307_, _38997_);
  nor _61466_ (_16308_, _16158_, _15540_);
  and _61467_ (_16309_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or _61468_ (_16310_, _16309_, _16308_);
  and _61469_ (_36913_[4], _16310_, _38997_);
  nor _61470_ (_16311_, _16158_, _15555_);
  and _61471_ (_16312_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or _61472_ (_16313_, _16312_, _16311_);
  and _61473_ (_36913_[5], _16313_, _38997_);
  nor _61474_ (_16314_, _16158_, _15576_);
  and _61475_ (_16315_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and _61476_ (_16316_, _16315_, _16158_);
  or _61477_ (_16317_, _16316_, _16314_);
  and _61478_ (_36913_[6], _16317_, _38997_);
  nor _61479_ (_16318_, _16158_, _15451_);
  and _61480_ (_16319_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or _61481_ (_16320_, _16319_, _16318_);
  and _61482_ (_36913_[7], _16320_, _38997_);
  and _61483_ (_16321_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and _61484_ (_16322_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or _61485_ (_16323_, _16322_, _16321_);
  and _61486_ (_36913_[8], _16323_, _38997_);
  and _61487_ (_16324_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and _61488_ (_16325_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or _61489_ (_16326_, _16325_, _16324_);
  and _61490_ (_36913_[9], _16326_, _38997_);
  and _61491_ (_16327_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and _61492_ (_16328_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or _61493_ (_16329_, _16328_, _16327_);
  and _61494_ (_36913_[10], _16329_, _38997_);
  and _61495_ (_16330_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and _61496_ (_16331_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or _61497_ (_16332_, _16331_, _16330_);
  and _61498_ (_36913_[11], _16332_, _38997_);
  and _61499_ (_16333_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and _61500_ (_16334_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or _61501_ (_16335_, _16334_, _16333_);
  and _61502_ (_36913_[12], _16335_, _38997_);
  and _61503_ (_16336_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and _61504_ (_16337_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or _61505_ (_16338_, _16337_, _16336_);
  and _61506_ (_36913_[13], _16338_, _38997_);
  and _61507_ (_16339_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and _61508_ (_16340_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or _61509_ (_16341_, _16340_, _16339_);
  and _61510_ (_36913_[14], _16341_, _38997_);
  and _61511_ (_16342_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and _61512_ (_16343_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or _61513_ (_16344_, _16343_, _16342_);
  and _61514_ (_36913_[15], _16344_, _38997_);
  and _61515_ (_16345_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and _61516_ (_16346_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or _61517_ (_16347_, _16346_, _16345_);
  and _61518_ (_36913_[16], _16347_, _38997_);
  and _61519_ (_16348_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and _61520_ (_16349_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or _61521_ (_16350_, _16349_, _16348_);
  and _61522_ (_36913_[17], _16350_, _38997_);
  and _61523_ (_16351_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and _61524_ (_16352_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or _61525_ (_16353_, _16352_, _16351_);
  and _61526_ (_36913_[18], _16353_, _38997_);
  and _61527_ (_16354_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and _61528_ (_16355_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or _61529_ (_16356_, _16355_, _16354_);
  and _61530_ (_36913_[19], _16356_, _38997_);
  and _61531_ (_16357_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and _61532_ (_16358_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or _61533_ (_16359_, _16358_, _16357_);
  and _61534_ (_36913_[20], _16359_, _38997_);
  and _61535_ (_16360_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and _61536_ (_16361_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or _61537_ (_16362_, _16361_, _16360_);
  and _61538_ (_36913_[21], _16362_, _38997_);
  and _61539_ (_16363_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and _61540_ (_16364_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or _61541_ (_16365_, _16364_, _16363_);
  and _61542_ (_36913_[22], _16365_, _38997_);
  and _61543_ (_16366_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and _61544_ (_16367_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or _61545_ (_16368_, _16367_, _16366_);
  and _61546_ (_36913_[23], _16368_, _38997_);
  and _61547_ (_16369_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and _61548_ (_16370_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or _61549_ (_16371_, _16370_, _16369_);
  and _61550_ (_36913_[24], _16371_, _38997_);
  and _61551_ (_16372_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and _61552_ (_16373_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or _61553_ (_16374_, _16373_, _16372_);
  and _61554_ (_36913_[25], _16374_, _38997_);
  and _61555_ (_16375_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and _61556_ (_16376_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or _61557_ (_16377_, _16376_, _16375_);
  and _61558_ (_36913_[26], _16377_, _38997_);
  and _61559_ (_16378_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and _61560_ (_16379_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or _61561_ (_16380_, _16379_, _16378_);
  and _61562_ (_36913_[27], _16380_, _38997_);
  and _61563_ (_16381_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and _61564_ (_16382_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or _61565_ (_16383_, _16382_, _16381_);
  and _61566_ (_36913_[28], _16383_, _38997_);
  and _61567_ (_16384_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and _61568_ (_16385_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or _61569_ (_16386_, _16385_, _16384_);
  and _61570_ (_36913_[29], _16386_, _38997_);
  and _61571_ (_16387_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and _61572_ (_16388_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or _61573_ (_16389_, _16388_, _16387_);
  and _61574_ (_36913_[30], _16389_, _38997_);
  nor _61575_ (_36893_[0], _34441_, rst);
  nor _61576_ (_36893_[1], _34548_, rst);
  nor _61577_ (_36893_[2], _34741_, rst);
  nor _61578_ (_36893_[3], _34391_, rst);
  nor _61579_ (_36893_[4], _34517_, rst);
  nor _61580_ (_36893_[5], _34634_, rst);
  nor _61581_ (_36893_[6], _34669_, rst);
  and _61582_ (_36898_[0], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _38997_);
  and _61583_ (_36898_[1], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _38997_);
  and _61584_ (_36898_[2], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _38997_);
  and _61585_ (_36898_[3], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _38997_);
  and _61586_ (_36898_[4], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _38997_);
  and _61587_ (_36898_[5], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _38997_);
  and _61588_ (_36898_[6], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _38997_);
  not _61589_ (_16390_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _61590_ (_16391_, _15696_, _16390_);
  and _61591_ (_16392_, _15021_, _33458_);
  and _61592_ (_16393_, _15689_, _16392_);
  nor _61593_ (_16394_, _15680_, _15842_);
  and _61594_ (_16395_, _16394_, _15679_);
  nor _61595_ (_16396_, _16395_, _16393_);
  and _61596_ (_16397_, _16396_, _15632_);
  and _61597_ (_16398_, _15621_, _34706_);
  and _61598_ (_16399_, _16398_, _33658_);
  nor _61599_ (_16400_, _16399_, _15685_);
  and _61600_ (_16401_, _16400_, _16397_);
  or _61601_ (_16402_, _15848_, _15826_);
  and _61602_ (_16403_, _16402_, _14223_);
  nor _61603_ (_16404_, _15827_, _15844_);
  and _61604_ (_16405_, _16404_, _15772_);
  and _61605_ (_16406_, _15828_, _15846_);
  and _61606_ (_16407_, _16406_, _15864_);
  and _61607_ (_16408_, _16407_, _15770_);
  or _61608_ (_16409_, _16408_, _16405_);
  nor _61609_ (_16410_, _15824_, _15839_);
  nor _61610_ (_16411_, _16406_, _16410_);
  nor _61611_ (_16412_, _15774_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _61612_ (_16413_, _16412_, _15775_);
  and _61613_ (_16414_, _16413_, _16411_);
  or _61614_ (_16415_, _16414_, _16409_);
  or _61615_ (_16416_, _16415_, _16403_);
  and _61616_ (_16417_, _16416_, _16401_);
  or _61617_ (_16418_, _16417_, _16391_);
  and _61618_ (_36899_[0], _16418_, _38997_);
  nand _61619_ (_16419_, _16402_, _14289_);
  nand _61620_ (_16420_, _15842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nand _61621_ (_16421_, _16404_, _15765_);
  nand _61622_ (_16422_, _16407_, _15763_);
  and _61623_ (_16423_, _16422_, _16421_);
  and _61624_ (_16424_, _16423_, _16420_);
  or _61625_ (_16425_, _15777_, _15775_);
  nand _61626_ (_16426_, _16425_, _16411_);
  or _61627_ (_16427_, _16426_, _15778_);
  and _61628_ (_16428_, _16427_, _16424_);
  and _61629_ (_16429_, _16428_, _16419_);
  nand _61630_ (_16430_, _16429_, _16401_);
  or _61631_ (_16431_, _16401_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _61632_ (_16432_, _16431_, _38997_);
  and _61633_ (_36899_[1], _16432_, _16430_);
  and _61634_ (_16433_, _16402_, _14724_);
  and _61635_ (_16434_, _15842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _61636_ (_16435_, _16404_, _15759_);
  and _61637_ (_16436_, _16407_, _15757_);
  or _61638_ (_16437_, _16436_, _16435_);
  or _61639_ (_16438_, _16437_, _16434_);
  or _61640_ (_16439_, _16438_, _16433_);
  not _61641_ (_16440_, _15783_);
  or _61642_ (_16441_, _15782_, _15779_);
  and _61643_ (_16442_, _16441_, _16440_);
  nand _61644_ (_16443_, _16442_, _16411_);
  nand _61645_ (_16444_, _16443_, _16401_);
  or _61646_ (_16445_, _16444_, _16439_);
  not _61647_ (_16446_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _61648_ (_16447_, _15699_, _16446_);
  and _61649_ (_16448_, _15699_, _16446_);
  nor _61650_ (_16449_, _16448_, _16447_);
  or _61651_ (_16450_, _16449_, _16401_);
  and _61652_ (_16451_, _16450_, _38997_);
  and _61653_ (_36899_[2], _16451_, _16445_);
  and _61654_ (_16452_, _16402_, _14740_);
  not _61655_ (_16453_, _15530_);
  and _61656_ (_16454_, _16404_, _16453_);
  not _61657_ (_16455_, _34417_);
  and _61658_ (_16456_, _16407_, _16455_);
  or _61659_ (_16457_, _16456_, _16454_);
  or _61660_ (_16458_, _15755_, _15756_);
  not _61661_ (_16459_, _16458_);
  nand _61662_ (_16460_, _16459_, _15784_);
  or _61663_ (_16461_, _16459_, _15784_);
  and _61664_ (_16462_, _16461_, _16411_);
  and _61665_ (_16463_, _16462_, _16460_);
  or _61666_ (_16464_, _16463_, _16457_);
  or _61667_ (_16465_, _16464_, _16452_);
  nand _61668_ (_16466_, _15842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nand _61669_ (_16467_, _16466_, _16401_);
  or _61670_ (_16468_, _16467_, _16465_);
  and _61671_ (_16469_, _16447_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _61672_ (_16470_, _16447_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _61673_ (_16471_, _16470_, _16469_);
  or _61674_ (_16472_, _16471_, _16401_);
  and _61675_ (_16473_, _16472_, _38997_);
  and _61676_ (_36899_[3], _16473_, _16468_);
  and _61677_ (_16474_, _15702_, _15700_);
  nor _61678_ (_16475_, _16469_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _61679_ (_16476_, _16475_, _16474_);
  or _61680_ (_16477_, _16476_, _15695_);
  and _61681_ (_16478_, _16477_, _38997_);
  and _61682_ (_16479_, _16402_, _14494_);
  or _61683_ (_16480_, _15788_, _15786_);
  and _61684_ (_16481_, _15830_, _15789_);
  and _61685_ (_16482_, _16481_, _16480_);
  not _61686_ (_16483_, _15548_);
  and _61687_ (_16484_, _15836_, _16483_);
  not _61688_ (_16485_, _34495_);
  and _61689_ (_16486_, _15865_, _16485_);
  and _61690_ (_16487_, _33469_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _61691_ (_16488_, _16487_, _16486_);
  or _61692_ (_16489_, _16488_, _16484_);
  nor _61693_ (_16490_, _16489_, _16482_);
  nand _61694_ (_16491_, _16490_, _15695_);
  or _61695_ (_16492_, _16491_, _16479_);
  and _61696_ (_36899_[4], _16492_, _16478_);
  nor _61697_ (_16493_, _16474_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _61698_ (_16494_, _16493_, _15704_);
  or _61699_ (_16495_, _16494_, _15695_);
  and _61700_ (_16496_, _16495_, _38997_);
  and _61701_ (_16497_, _16402_, _14767_);
  or _61702_ (_16498_, _15746_, _15747_);
  and _61703_ (_16499_, _16498_, _15790_);
  nor _61704_ (_16500_, _16498_, _15790_);
  or _61705_ (_16501_, _16500_, _16499_);
  and _61706_ (_16502_, _16501_, _15830_);
  not _61707_ (_16503_, _15566_);
  and _61708_ (_16504_, _15836_, _16503_);
  not _61709_ (_16505_, _34603_);
  and _61710_ (_16506_, _15865_, _16505_);
  and _61711_ (_16507_, _33469_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _61712_ (_16508_, _16507_, _16506_);
  or _61713_ (_16509_, _16508_, _16504_);
  nor _61714_ (_16510_, _16509_, _16502_);
  nand _61715_ (_16511_, _16510_, _15695_);
  or _61716_ (_16512_, _16511_, _16497_);
  and _61717_ (_36899_[5], _16512_, _16496_);
  nor _61718_ (_16513_, _15704_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _61719_ (_16514_, _16513_, _15705_);
  or _61720_ (_16515_, _16514_, _15695_);
  and _61721_ (_16516_, _16515_, _38997_);
  and _61722_ (_16517_, _15842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _61723_ (_16518_, _16402_, _14632_);
  not _61724_ (_16519_, _15584_);
  and _61725_ (_16520_, _16404_, _16519_);
  and _61726_ (_16521_, _16407_, _34686_);
  or _61727_ (_16522_, _16521_, _16520_);
  or _61728_ (_16523_, _15792_, _15742_);
  and _61729_ (_16524_, _16411_, _15793_);
  and _61730_ (_16525_, _16524_, _16523_);
  or _61731_ (_16526_, _16525_, _16522_);
  or _61732_ (_16527_, _16526_, _16518_);
  nor _61733_ (_16528_, _16527_, _16517_);
  nand _61734_ (_16529_, _16528_, _16401_);
  and _61735_ (_36899_[6], _16529_, _16516_);
  nor _61736_ (_16530_, _15705_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _61737_ (_16531_, _16530_, _15706_);
  or _61738_ (_16532_, _16531_, _15695_);
  and _61739_ (_16533_, _16532_, _38997_);
  or _61740_ (_16534_, _15733_, _15734_);
  and _61741_ (_16535_, _16534_, _15794_);
  nor _61742_ (_16536_, _16534_, _15794_);
  or _61743_ (_16537_, _16536_, _16535_);
  and _61744_ (_16538_, _16537_, _16411_);
  and _61745_ (_16539_, _16402_, _14683_);
  and _61746_ (_16540_, _15842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _61747_ (_16541_, _15459_);
  and _61748_ (_16542_, _16404_, _16541_);
  and _61749_ (_16543_, _16407_, _15835_);
  or _61750_ (_16544_, _16543_, _16542_);
  or _61751_ (_16545_, _16544_, _16540_);
  or _61752_ (_16546_, _16545_, _16539_);
  nor _61753_ (_16547_, _16546_, _16538_);
  nand _61754_ (_16548_, _16547_, _16401_);
  and _61755_ (_36899_[7], _16548_, _16533_);
  nor _61756_ (_16549_, _15706_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _61757_ (_16550_, _16549_, _15707_);
  or _61758_ (_16551_, _16550_, _15695_);
  and _61759_ (_16552_, _16551_, _38997_);
  and _61760_ (_16553_, _15796_, _14110_);
  nor _61761_ (_16554_, _15796_, _14110_);
  nor _61762_ (_16555_, _16554_, _16553_);
  nor _61763_ (_16556_, _16555_, _15732_);
  and _61764_ (_16557_, _16555_, _15732_);
  or _61765_ (_16558_, _16557_, _16556_);
  and _61766_ (_16559_, _16558_, _15830_);
  and _61767_ (_16560_, _14223_, _33469_);
  and _61768_ (_16561_, _15826_, _14250_);
  nand _61769_ (_16562_, _15836_, _15770_);
  and _61770_ (_16563_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _61771_ (_16564_, _15865_, _14930_);
  nor _61772_ (_16565_, _16564_, _16563_);
  and _61773_ (_16566_, _16565_, _16562_);
  nand _61774_ (_16567_, _16566_, _15695_);
  or _61775_ (_16568_, _16567_, _16561_);
  or _61776_ (_16569_, _16568_, _16560_);
  or _61777_ (_16570_, _16569_, _16559_);
  and _61778_ (_36899_[8], _16570_, _16552_);
  nor _61779_ (_16571_, _15707_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _61780_ (_16572_, _16571_, _15708_);
  or _61781_ (_16573_, _16572_, _15695_);
  and _61782_ (_16574_, _16573_, _38997_);
  and _61783_ (_16575_, _15796_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _61784_ (_16576_, _16575_, _15804_);
  nor _61785_ (_16577_, _15805_, _15804_);
  nor _61786_ (_16578_, _16577_, _16576_);
  nand _61787_ (_16579_, _16578_, _14116_);
  or _61788_ (_16580_, _16578_, _14116_);
  and _61789_ (_16581_, _16580_, _15830_);
  and _61790_ (_16582_, _16581_, _16579_);
  and _61791_ (_16583_, _14289_, _33469_);
  nor _61792_ (_16584_, _15833_, _14323_);
  and _61793_ (_16585_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _61794_ (_16586_, _15836_, _15763_);
  or _61795_ (_16587_, _16586_, _16585_);
  and _61796_ (_16588_, _15865_, _33344_);
  or _61797_ (_16589_, _16588_, _16587_);
  nor _61798_ (_16590_, _16589_, _16584_);
  nand _61799_ (_16591_, _16590_, _15695_);
  or _61800_ (_16592_, _16591_, _16583_);
  or _61801_ (_16593_, _16592_, _16582_);
  and _61802_ (_36899_[9], _16593_, _16574_);
  nor _61803_ (_16594_, _15708_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _61804_ (_16595_, _16594_, _15709_);
  or _61805_ (_16596_, _16595_, _15695_);
  and _61806_ (_16597_, _16596_, _38997_);
  and _61807_ (_16598_, _16577_, _14116_);
  and _61808_ (_16599_, _16576_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _61809_ (_16600_, _16599_, _16598_);
  nand _61810_ (_16601_, _16600_, _14121_);
  or _61811_ (_16602_, _16600_, _14121_);
  and _61812_ (_16603_, _16602_, _15830_);
  and _61813_ (_16604_, _16603_, _16601_);
  nor _61814_ (_16605_, _14356_, _33470_);
  nor _61815_ (_16606_, _15833_, _14387_);
  and _61816_ (_16607_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _61817_ (_16608_, _15836_, _15757_);
  and _61818_ (_16609_, _15865_, _14931_);
  or _61819_ (_16610_, _16609_, _16608_);
  or _61820_ (_16611_, _16610_, _16607_);
  nor _61821_ (_16612_, _16611_, _16606_);
  nand _61822_ (_16613_, _16612_, _15695_);
  or _61823_ (_16614_, _16613_, _16605_);
  or _61824_ (_16615_, _16614_, _16604_);
  and _61825_ (_36899_[10], _16615_, _16597_);
  nor _61826_ (_16616_, _15709_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _61827_ (_16617_, _15709_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _61828_ (_16618_, _16617_, _16616_);
  or _61829_ (_16619_, _16618_, _15695_);
  and _61830_ (_16620_, _16619_, _38997_);
  and _61831_ (_16621_, _15799_, _15804_);
  nor _61832_ (_16622_, _15807_, _15804_);
  nor _61833_ (_16623_, _16622_, _16621_);
  nor _61834_ (_16624_, _16623_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _61835_ (_16625_, _16623_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _61836_ (_16626_, _16625_, _16624_);
  and _61837_ (_16627_, _16626_, _15830_);
  nor _61838_ (_16628_, _14423_, _33470_);
  nor _61839_ (_16629_, _15833_, _14456_);
  and _61840_ (_16630_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _61841_ (_16631_, _15836_, _16455_);
  or _61842_ (_16632_, _16631_, _16630_);
  nor _61843_ (_16633_, _15856_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _61844_ (_16634_, _16633_, _15857_);
  and _61845_ (_16635_, _16634_, _15865_);
  or _61846_ (_16636_, _16635_, _16632_);
  nor _61847_ (_16637_, _16636_, _16629_);
  nand _61848_ (_16638_, _16637_, _15695_);
  or _61849_ (_16639_, _16638_, _16628_);
  or _61850_ (_16640_, _16639_, _16627_);
  and _61851_ (_36899_[11], _16640_, _16620_);
  nor _61852_ (_16641_, _16617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _61853_ (_16642_, _16641_, _15711_);
  or _61854_ (_16643_, _16642_, _15695_);
  and _61855_ (_16644_, _16643_, _38997_);
  nor _61856_ (_16645_, _15808_, _15804_);
  and _61857_ (_16646_, _15800_, _15804_);
  or _61858_ (_16647_, _16646_, _16645_);
  nand _61859_ (_16648_, _16647_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _61860_ (_16649_, _16647_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _61861_ (_16650_, _16649_, _15830_);
  and _61862_ (_16651_, _16650_, _16648_);
  and _61863_ (_16652_, _14494_, _33469_);
  nor _61864_ (_16653_, _15833_, _14529_);
  and _61865_ (_16654_, _15836_, _16485_);
  and _61866_ (_16655_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _61867_ (_16656_, _15857_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _61868_ (_16657_, _16656_, _15858_);
  and _61869_ (_16658_, _16657_, _15865_);
  or _61870_ (_16659_, _16658_, _16655_);
  or _61871_ (_16660_, _16659_, _16654_);
  nor _61872_ (_16661_, _16660_, _16653_);
  nand _61873_ (_16662_, _16661_, _15695_);
  or _61874_ (_16663_, _16662_, _16652_);
  or _61875_ (_16664_, _16663_, _16651_);
  and _61876_ (_36899_[12], _16664_, _16644_);
  not _61877_ (_16665_, _16401_);
  or _61878_ (_16666_, _15809_, _15804_);
  nand _61879_ (_16667_, _16646_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _61880_ (_16668_, _16667_, _16666_);
  nor _61881_ (_16669_, _16668_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _61882_ (_16670_, _16668_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _61883_ (_16671_, _16670_, _16669_);
  and _61884_ (_16672_, _16671_, _15830_);
  nor _61885_ (_16673_, _14570_, _33470_);
  nor _61886_ (_16674_, _15833_, _14602_);
  and _61887_ (_16675_, _15836_, _16505_);
  and _61888_ (_16676_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _61889_ (_16677_, _15858_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _61890_ (_16678_, _16677_, _15859_);
  and _61891_ (_16679_, _16678_, _15865_);
  or _61892_ (_16680_, _16679_, _16676_);
  or _61893_ (_16681_, _16680_, _16675_);
  or _61894_ (_16682_, _16681_, _16674_);
  or _61895_ (_16683_, _16682_, _16673_);
  or _61896_ (_16684_, _16683_, _16672_);
  or _61897_ (_16685_, _16684_, _16665_);
  nor _61898_ (_16686_, _15711_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _61899_ (_16687_, _16686_, _15712_);
  or _61900_ (_16688_, _16687_, _16401_);
  and _61901_ (_16689_, _16688_, _38997_);
  and _61902_ (_36899_[13], _16689_, _16685_);
  and _61903_ (_16690_, _14632_, _33469_);
  and _61904_ (_16691_, _15826_, _14659_);
  and _61905_ (_16692_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _61906_ (_16693_, _15836_, _34686_);
  or _61907_ (_16694_, _16693_, _16692_);
  or _61908_ (_16695_, _15859_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _61909_ (_16696_, _16695_, _15860_);
  and _61910_ (_16697_, _16696_, _15865_);
  or _61911_ (_16698_, _16697_, _16694_);
  or _61912_ (_16699_, _16698_, _16691_);
  or _61913_ (_16700_, _16699_, _16690_);
  and _61914_ (_16701_, _15811_, _15803_);
  nor _61915_ (_16702_, _16701_, _14137_);
  and _61916_ (_16703_, _16701_, _14137_);
  or _61917_ (_16704_, _16703_, _16702_);
  and _61918_ (_16705_, _16704_, _16411_);
  or _61919_ (_16706_, _16705_, _16700_);
  or _61920_ (_16707_, _16706_, _16665_);
  nor _61921_ (_16708_, _15712_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _61922_ (_16709_, _16708_, _15713_);
  or _61923_ (_16710_, _16709_, _16401_);
  and _61924_ (_16711_, _16710_, _38997_);
  and _61925_ (_36899_[14], _16711_, _16707_);
  and _61926_ (_16712_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _61927_ (_16713_, _16059_, _16057_);
  nor _61928_ (_16714_, _16713_, _16060_);
  or _61929_ (_16715_, _16714_, _15877_);
  or _61930_ (_16716_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _61931_ (_16717_, _16716_, _16091_);
  and _61932_ (_16718_, _16717_, _16715_);
  or _61933_ (_36900_[0], _16718_, _16712_);
  and _61934_ (_16719_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _61935_ (_16720_, _16062_, _16060_);
  and _61936_ (_16721_, _16720_, _16063_);
  or _61937_ (_16722_, _16721_, _15877_);
  or _61938_ (_16723_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _61939_ (_16724_, _16723_, _16091_);
  and _61940_ (_16725_, _16724_, _16722_);
  or _61941_ (_36900_[1], _16725_, _16719_);
  and _61942_ (_16726_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _61943_ (_16727_, _16067_, _16065_);
  nor _61944_ (_16728_, _16727_, _16068_);
  or _61945_ (_16729_, _16728_, _15877_);
  or _61946_ (_16730_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _61947_ (_16731_, _16730_, _16091_);
  and _61948_ (_16732_, _16731_, _16729_);
  or _61949_ (_36900_[2], _16732_, _16726_);
  and _61950_ (_16733_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _61951_ (_16734_, _16068_, _15952_);
  nor _61952_ (_16735_, _16734_, _16069_);
  or _61953_ (_16736_, _16735_, _15877_);
  or _61954_ (_16737_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _61955_ (_16738_, _16737_, _16091_);
  and _61956_ (_16739_, _16738_, _16736_);
  or _61957_ (_36900_[3], _16739_, _16733_);
  nor _61958_ (_16740_, _16072_, _16069_);
  nor _61959_ (_16741_, _16740_, _16073_);
  or _61960_ (_16742_, _16741_, _15877_);
  or _61961_ (_16743_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _61962_ (_16744_, _16743_, _16091_);
  and _61963_ (_16745_, _16744_, _16742_);
  and _61964_ (_16746_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _61965_ (_36900_[4], _16746_, _16745_);
  nor _61966_ (_16747_, _16073_, _15947_);
  nor _61967_ (_16748_, _16747_, _16074_);
  or _61968_ (_16749_, _16748_, _15877_);
  or _61969_ (_16750_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _61970_ (_16751_, _16750_, _16091_);
  and _61971_ (_16752_, _16751_, _16749_);
  and _61972_ (_16753_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _61973_ (_36900_[5], _16753_, _16752_);
  nor _61974_ (_16754_, _16074_, _15943_);
  nor _61975_ (_16755_, _16754_, _16075_);
  or _61976_ (_16756_, _16755_, _15877_);
  or _61977_ (_16757_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _61978_ (_16758_, _16757_, _16091_);
  and _61979_ (_16759_, _16758_, _16756_);
  and _61980_ (_16760_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _61981_ (_36900_[6], _16760_, _16759_);
  and _61982_ (_16761_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _61983_ (_16762_, _16075_, _15939_);
  nor _61984_ (_16763_, _16762_, _16076_);
  or _61985_ (_16764_, _16763_, _15877_);
  or _61986_ (_16765_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _61987_ (_16766_, _16765_, _16091_);
  and _61988_ (_16767_, _16766_, _16764_);
  or _61989_ (_36900_[7], _16767_, _16761_);
  or _61990_ (_16768_, _16078_, _16076_);
  nor _61991_ (_16769_, _16079_, _15877_);
  and _61992_ (_16770_, _16769_, _16768_);
  nor _61993_ (_16771_, _15876_, _14110_);
  or _61994_ (_16772_, _16771_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _61995_ (_16773_, _16772_, _16770_);
  or _61996_ (_16774_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _33132_);
  and _61997_ (_16775_, _16774_, _38997_);
  and _61998_ (_36900_[8], _16775_, _16773_);
  nor _61999_ (_16776_, _16079_, _15934_);
  nor _62000_ (_16777_, _16776_, _16080_);
  or _62001_ (_16778_, _16777_, _15877_);
  or _62002_ (_16779_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _62003_ (_16780_, _16779_, _16091_);
  and _62004_ (_16781_, _16780_, _16778_);
  and _62005_ (_16782_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _62006_ (_36900_[9], _16782_, _16781_);
  nor _62007_ (_16783_, _16080_, _15931_);
  nor _62008_ (_16784_, _16783_, _16081_);
  or _62009_ (_16785_, _16784_, _15877_);
  or _62010_ (_16786_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _62011_ (_16787_, _16786_, _16091_);
  and _62012_ (_16788_, _16787_, _16785_);
  and _62013_ (_16789_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _62014_ (_36900_[10], _16789_, _16788_);
  and _62015_ (_16790_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _62016_ (_16791_, _16081_, _15927_);
  nor _62017_ (_16792_, _16791_, _16082_);
  or _62018_ (_16793_, _16792_, _15877_);
  or _62019_ (_16794_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _62020_ (_16795_, _16794_, _16091_);
  and _62021_ (_16796_, _16795_, _16793_);
  or _62022_ (_36900_[11], _16796_, _16790_);
  nor _62023_ (_16797_, _16082_, _15923_);
  nor _62024_ (_16798_, _16797_, _16083_);
  or _62025_ (_16799_, _16798_, _15877_);
  or _62026_ (_16800_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _62027_ (_16801_, _16800_, _16091_);
  and _62028_ (_16802_, _16801_, _16799_);
  and _62029_ (_16803_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _62030_ (_36900_[12], _16803_, _16802_);
  nor _62031_ (_16804_, _16083_, _15920_);
  nor _62032_ (_16805_, _16804_, _16084_);
  or _62033_ (_16806_, _16805_, _15877_);
  or _62034_ (_16807_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _62035_ (_16808_, _16807_, _16091_);
  and _62036_ (_16809_, _16808_, _16806_);
  and _62037_ (_16810_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _62038_ (_36900_[13], _16810_, _16809_);
  nor _62039_ (_16811_, _16084_, _15917_);
  nor _62040_ (_16812_, _16811_, _16085_);
  or _62041_ (_16813_, _16812_, _15877_);
  or _62042_ (_16814_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _62043_ (_16815_, _16814_, _16091_);
  and _62044_ (_16816_, _16815_, _16813_);
  and _62045_ (_16817_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _62046_ (_36900_[14], _16817_, _16816_);
  and _62047_ (_16818_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _62048_ (_16819_, _16818_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _62049_ (_36904_[0], _16819_, _38997_);
  and _62050_ (_16820_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _62051_ (_16821_, _16820_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _62052_ (_36904_[1], _16821_, _38997_);
  and _62053_ (_16822_, _16102_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or _62054_ (_16823_, _16822_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _62055_ (_36904_[2], _16823_, _38997_);
  and _62056_ (_16824_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _62057_ (_16825_, _16824_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _62058_ (_36904_[3], _16825_, _38997_);
  and _62059_ (_16826_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _62060_ (_16827_, _16826_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _62061_ (_36904_[4], _16827_, _38997_);
  and _62062_ (_16828_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _62063_ (_16829_, _16828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _62064_ (_36904_[5], _16829_, _38997_);
  and _62065_ (_16830_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or _62066_ (_16831_, _16830_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _62067_ (_36904_[6], _16831_, _38997_);
  nor _62068_ (_16832_, _16056_, _34325_);
  nand _62069_ (_16833_, _16832_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _62070_ (_16834_, _16832_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _62071_ (_16835_, _16834_, _16091_);
  and _62072_ (_36905_[0], _16835_, _16833_);
  or _62073_ (_16836_, _16115_, _16113_);
  and _62074_ (_16837_, _16836_, _16116_);
  or _62075_ (_16838_, _16837_, _34325_);
  or _62076_ (_16839_, _33135_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _62077_ (_16840_, _16839_, _16091_);
  and _62078_ (_36905_[1], _16840_, _16838_);
  and _62079_ (_16841_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and _62080_ (_16842_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and _62081_ (_16843_, _16842_, _36910_);
  or _62082_ (_36909_[0], _16843_, _16841_);
  and _62083_ (_16844_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and _62084_ (_16845_, _16298_, _36910_);
  or _62085_ (_36909_[1], _16845_, _16844_);
  and _62086_ (_16846_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and _62087_ (_16847_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and _62088_ (_16848_, _16847_, _36910_);
  or _62089_ (_36909_[2], _16848_, _16846_);
  and _62090_ (_16849_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and _62091_ (_16850_, _16305_, _36910_);
  or _62092_ (_36909_[3], _16850_, _16849_);
  and _62093_ (_16851_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and _62094_ (_16852_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and _62095_ (_16853_, _16852_, _36910_);
  or _62096_ (_36909_[4], _16853_, _16851_);
  and _62097_ (_16854_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and _62098_ (_16855_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and _62099_ (_16856_, _16855_, _36910_);
  or _62100_ (_36909_[5], _16856_, _16854_);
  and _62101_ (_16857_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and _62102_ (_16858_, _16315_, _36910_);
  or _62103_ (_36909_[6], _16858_, _16857_);
  and _62104_ (_36912_[0], _16144_, _38997_);
  nor _62105_ (_36912_[1], _16154_, rst);
  and _62106_ (_36912_[2], _16150_, _38997_);
  or _62107_ (_16859_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nand _62108_ (_16860_, _16158_, _15469_);
  and _62109_ (_16861_, _16860_, _38997_);
  and _62110_ (_36914_[0], _16861_, _16859_);
  and _62111_ (_16862_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _62112_ (_16863_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or _62113_ (_16864_, _16863_, _16862_);
  and _62114_ (_36914_[1], _16864_, _38997_);
  or _62115_ (_16865_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand _62116_ (_16866_, _16158_, _15501_);
  and _62117_ (_16867_, _16866_, _38997_);
  and _62118_ (_36914_[2], _16867_, _16865_);
  or _62119_ (_16868_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand _62120_ (_16869_, _16158_, _15522_);
  and _62121_ (_16870_, _16869_, _38997_);
  and _62122_ (_36914_[3], _16870_, _16868_);
  or _62123_ (_16871_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nand _62124_ (_16872_, _16158_, _15540_);
  and _62125_ (_16873_, _16872_, _38997_);
  and _62126_ (_36914_[4], _16873_, _16871_);
  or _62127_ (_16874_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand _62128_ (_16875_, _16158_, _15555_);
  and _62129_ (_16876_, _16875_, _38997_);
  and _62130_ (_36914_[5], _16876_, _16874_);
  or _62131_ (_16877_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand _62132_ (_16878_, _16158_, _15576_);
  and _62133_ (_16879_, _16878_, _38997_);
  and _62134_ (_36914_[6], _16879_, _16877_);
  or _62135_ (_16880_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand _62136_ (_16881_, _16158_, _15451_);
  and _62137_ (_16882_, _16881_, _38997_);
  and _62138_ (_36914_[7], _16882_, _16880_);
  and _62139_ (_16883_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _62140_ (_16884_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or _62141_ (_16885_, _16884_, _16883_);
  and _62142_ (_36914_[8], _16885_, _38997_);
  and _62143_ (_16886_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _62144_ (_16887_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or _62145_ (_16888_, _16887_, _16886_);
  and _62146_ (_36914_[9], _16888_, _38997_);
  and _62147_ (_16889_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _62148_ (_16890_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or _62149_ (_16891_, _16890_, _16889_);
  and _62150_ (_36914_[10], _16891_, _38997_);
  and _62151_ (_16892_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _62152_ (_16893_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or _62153_ (_16894_, _16893_, _16892_);
  and _62154_ (_36914_[11], _16894_, _38997_);
  and _62155_ (_16895_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _62156_ (_16896_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _62157_ (_16897_, _16896_, _16895_);
  and _62158_ (_36914_[12], _16897_, _38997_);
  and _62159_ (_16898_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _62160_ (_16899_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or _62161_ (_16900_, _16899_, _16898_);
  and _62162_ (_36914_[13], _16900_, _38997_);
  and _62163_ (_16901_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _62164_ (_16902_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or _62165_ (_16903_, _16902_, _16901_);
  and _62166_ (_36914_[14], _16903_, _38997_);
  and _62167_ (_16904_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _62168_ (_16905_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or _62169_ (_16906_, _16905_, _16904_);
  and _62170_ (_36914_[15], _16906_, _38997_);
  and _62171_ (_16907_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor _62172_ (_16908_, _16158_, _33206_);
  or _62173_ (_16909_, _16908_, _16907_);
  and _62174_ (_36914_[16], _16909_, _38997_);
  and _62175_ (_16910_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _62176_ (_16911_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _62177_ (_16912_, _16911_, _16910_);
  and _62178_ (_36914_[17], _16912_, _38997_);
  and _62179_ (_16913_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor _62180_ (_16914_, _16158_, _33142_);
  or _62181_ (_16915_, _16914_, _16913_);
  and _62182_ (_36914_[18], _16915_, _38997_);
  and _62183_ (_16916_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor _62184_ (_16917_, _16158_, _33184_);
  or _62185_ (_16918_, _16917_, _16916_);
  and _62186_ (_36914_[19], _16918_, _38997_);
  and _62187_ (_16919_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor _62188_ (_16920_, _16158_, _33256_);
  or _62189_ (_16921_, _16920_, _16919_);
  and _62190_ (_36914_[20], _16921_, _38997_);
  and _62191_ (_16922_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor _62192_ (_16923_, _16158_, _33285_);
  or _62193_ (_16924_, _16923_, _16922_);
  and _62194_ (_36914_[21], _16924_, _38997_);
  and _62195_ (_16925_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor _62196_ (_16926_, _16158_, _33331_);
  or _62197_ (_16927_, _16926_, _16925_);
  and _62198_ (_36914_[22], _16927_, _38997_);
  and _62199_ (_16928_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor _62200_ (_16929_, _16158_, _33303_);
  or _62201_ (_16930_, _16929_, _16928_);
  and _62202_ (_36914_[23], _16930_, _38997_);
  and _62203_ (_16931_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor _62204_ (_16932_, _16158_, _34445_);
  or _62205_ (_16933_, _16932_, _16931_);
  and _62206_ (_36914_[24], _16933_, _38997_);
  and _62207_ (_16934_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _62208_ (_16935_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _62209_ (_16936_, _16935_, _16934_);
  and _62210_ (_36914_[25], _16936_, _38997_);
  and _62211_ (_16937_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nor _62212_ (_16938_, _16158_, _34747_);
  or _62213_ (_16939_, _16938_, _16937_);
  and _62214_ (_36914_[26], _16939_, _38997_);
  and _62215_ (_16940_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor _62216_ (_16941_, _16158_, _34405_);
  or _62217_ (_16942_, _16941_, _16940_);
  and _62218_ (_36914_[27], _16942_, _38997_);
  and _62219_ (_16943_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor _62220_ (_16944_, _16158_, _34483_);
  or _62221_ (_16945_, _16944_, _16943_);
  and _62222_ (_36914_[28], _16945_, _38997_);
  and _62223_ (_16946_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor _62224_ (_16947_, _16158_, _34591_);
  or _62225_ (_16948_, _16947_, _16946_);
  and _62226_ (_36914_[29], _16948_, _38997_);
  and _62227_ (_16949_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor _62228_ (_16950_, _16158_, _34673_);
  or _62229_ (_16951_, _16950_, _16949_);
  and _62230_ (_36914_[30], _16951_, _38997_);
  and _62231_ (_16952_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _62232_ (_16953_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _62233_ (_16954_, _16953_, _16952_);
  and _62234_ (_36915_[0], _16954_, _38997_);
  and _62235_ (_16955_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _62236_ (_16956_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _62237_ (_16957_, _16956_, _16955_);
  and _62238_ (_36915_[1], _16957_, _38997_);
  and _62239_ (_16958_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _62240_ (_16959_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _62241_ (_16960_, _16959_, _16958_);
  and _62242_ (_36915_[2], _16960_, _38997_);
  and _62243_ (_16961_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _62244_ (_16962_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _62245_ (_16963_, _16962_, _16961_);
  and _62246_ (_36915_[3], _16963_, _38997_);
  and _62247_ (_16964_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _62248_ (_16965_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _62249_ (_16966_, _16965_, _16964_);
  and _62250_ (_36915_[4], _16966_, _38997_);
  and _62251_ (_16967_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _62252_ (_16968_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _62253_ (_16969_, _16968_, _16967_);
  and _62254_ (_36915_[5], _16969_, _38997_);
  and _62255_ (_16970_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _62256_ (_16971_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _62257_ (_16972_, _16971_, _16970_);
  and _62258_ (_36915_[6], _16972_, _38997_);
  and _62259_ (_16973_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _62260_ (_16974_, _34441_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _62261_ (_16975_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _62262_ (_16976_, _16975_, _16167_);
  and _62263_ (_16977_, _16976_, _16974_);
  or _62264_ (_16978_, _16977_, _16973_);
  and _62265_ (_36918_[0], _16978_, _38997_);
  and _62266_ (_16979_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _62267_ (_16980_, _34548_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _62268_ (_16981_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _62269_ (_16982_, _16981_, _16167_);
  and _62270_ (_16983_, _16982_, _16980_);
  or _62271_ (_16984_, _16983_, _16979_);
  and _62272_ (_36918_[1], _16984_, _38997_);
  and _62273_ (_16985_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _62274_ (_16986_, _34741_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _62275_ (_16987_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _62276_ (_16988_, _16987_, _16167_);
  and _62277_ (_16989_, _16988_, _16986_);
  or _62278_ (_16990_, _16989_, _16985_);
  and _62279_ (_36918_[2], _16990_, _38997_);
  and _62280_ (_16991_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _62281_ (_16992_, _34391_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _62282_ (_16993_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _62283_ (_16994_, _16993_, _16167_);
  and _62284_ (_16995_, _16994_, _16992_);
  or _62285_ (_16996_, _16995_, _16991_);
  and _62286_ (_36918_[3], _16996_, _38997_);
  and _62287_ (_16997_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _62288_ (_16998_, _34517_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _62289_ (_16999_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _62290_ (_17000_, _16999_, _16167_);
  and _62291_ (_17001_, _17000_, _16998_);
  or _62292_ (_17002_, _17001_, _16997_);
  and _62293_ (_36918_[4], _17002_, _38997_);
  and _62294_ (_17003_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _62295_ (_17004_, _34634_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _62296_ (_17005_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _62297_ (_17006_, _17005_, _16167_);
  and _62298_ (_17007_, _17006_, _17004_);
  or _62299_ (_17008_, _17007_, _17003_);
  and _62300_ (_36918_[5], _17008_, _38997_);
  and _62301_ (_17009_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _62302_ (_17010_, _34669_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _62303_ (_17011_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _62304_ (_17012_, _17011_, _16167_);
  and _62305_ (_17013_, _17012_, _17010_);
  or _62306_ (_17014_, _17013_, _17009_);
  and _62307_ (_36918_[6], _17014_, _38997_);
  and _62308_ (_17015_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _62309_ (_17016_, _34320_, _16174_);
  or _62310_ (_17017_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _62311_ (_17018_, _17017_, _16167_);
  and _62312_ (_17019_, _17018_, _17016_);
  or _62313_ (_17020_, _17019_, _17015_);
  and _62314_ (_36918_[7], _17020_, _38997_);
  and _62315_ (_17021_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _62316_ (_17022_, _17021_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _62317_ (_17023_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _16167_);
  and _62318_ (_17024_, _17023_, _38997_);
  and _62319_ (_36918_[8], _17024_, _17022_);
  and _62320_ (_17025_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _62321_ (_17026_, _17025_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _62322_ (_17027_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _16167_);
  and _62323_ (_17028_, _17027_, _38997_);
  and _62324_ (_36918_[9], _17028_, _17026_);
  and _62325_ (_17029_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _62326_ (_17030_, _17029_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _62327_ (_17031_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _16167_);
  and _62328_ (_17032_, _17031_, _38997_);
  and _62329_ (_36918_[10], _17032_, _17030_);
  and _62330_ (_17033_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _62331_ (_17034_, _17033_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _62332_ (_17035_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _16167_);
  and _62333_ (_17036_, _17035_, _38997_);
  and _62334_ (_36918_[11], _17036_, _17034_);
  and _62335_ (_17037_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _62336_ (_17038_, _17037_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _62337_ (_17039_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _16167_);
  and _62338_ (_17040_, _17039_, _38997_);
  and _62339_ (_36918_[12], _17040_, _17038_);
  and _62340_ (_17041_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _62341_ (_17042_, _17041_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _62342_ (_17043_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _16167_);
  and _62343_ (_17044_, _17043_, _38997_);
  and _62344_ (_36918_[13], _17044_, _17042_);
  and _62345_ (_17045_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _62346_ (_17046_, _17045_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _62347_ (_17047_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _16167_);
  and _62348_ (_17048_, _17047_, _38997_);
  and _62349_ (_36918_[14], _17048_, _17046_);
  not _62350_ (_17049_, _16181_);
  or _62351_ (_17050_, _17049_, _14223_);
  or _62352_ (_17051_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _62353_ (_17052_, _17051_, _38997_);
  and _62354_ (_36922_[0], _17052_, _17050_);
  or _62355_ (_17053_, _17049_, _14289_);
  or _62356_ (_17054_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _62357_ (_17055_, _17054_, _38997_);
  and _62358_ (_36922_[1], _17055_, _17053_);
  nand _62359_ (_17056_, _16181_, _14356_);
  or _62360_ (_17057_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _62361_ (_17058_, _17057_, _38997_);
  and _62362_ (_36922_[2], _17058_, _17056_);
  nand _62363_ (_17059_, _16181_, _14423_);
  or _62364_ (_17060_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _62365_ (_17061_, _17060_, _38997_);
  and _62366_ (_36922_[3], _17061_, _17059_);
  or _62367_ (_17062_, _17049_, _14494_);
  or _62368_ (_17063_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and _62369_ (_17064_, _17063_, _38997_);
  and _62370_ (_36922_[4], _17064_, _17062_);
  nand _62371_ (_17065_, _16181_, _14570_);
  or _62372_ (_17066_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and _62373_ (_17067_, _17066_, _38997_);
  and _62374_ (_36922_[5], _17067_, _17065_);
  or _62375_ (_17068_, _17049_, _14632_);
  or _62376_ (_17069_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and _62377_ (_17070_, _17069_, _38997_);
  and _62378_ (_36922_[6], _17070_, _17068_);
  nand _62379_ (_17071_, _16181_, _14098_);
  or _62380_ (_17072_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and _62381_ (_17073_, _17072_, _38997_);
  and _62382_ (_36922_[7], _17073_, _17071_);
  or _62383_ (_17074_, _17049_, _14250_);
  or _62384_ (_17075_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and _62385_ (_17076_, _17075_, _38997_);
  and _62386_ (_36922_[8], _17076_, _17074_);
  nand _62387_ (_17077_, _16181_, _14323_);
  or _62388_ (_17078_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and _62389_ (_17079_, _17078_, _38997_);
  and _62390_ (_36922_[9], _17079_, _17077_);
  nand _62391_ (_17080_, _16181_, _14387_);
  or _62392_ (_17081_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and _62393_ (_17082_, _17081_, _38997_);
  and _62394_ (_36922_[10], _17082_, _17080_);
  nand _62395_ (_17083_, _16181_, _14456_);
  or _62396_ (_17084_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and _62397_ (_17085_, _17084_, _38997_);
  and _62398_ (_36922_[11], _17085_, _17083_);
  nand _62399_ (_17086_, _16181_, _14529_);
  or _62400_ (_17087_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and _62401_ (_17088_, _17087_, _38997_);
  and _62402_ (_36922_[12], _17088_, _17086_);
  nand _62403_ (_17089_, _16181_, _14602_);
  or _62404_ (_17090_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and _62405_ (_17091_, _17090_, _38997_);
  and _62406_ (_36922_[13], _17091_, _17089_);
  or _62407_ (_17092_, _17049_, _14659_);
  or _62408_ (_17093_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and _62409_ (_17094_, _17093_, _38997_);
  and _62410_ (_36922_[14], _17094_, _17092_);
  nor _62411_ (_36880_, _34369_, rst);
  and _62412_ (_17095_, _34258_, _34247_);
  nand _62413_ (_17096_, _17095_, _34221_);
  or _62414_ (_17097_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _62415_ (_17098_, _17097_, _38997_);
  and _62416_ (_36881_[7], _17098_, _17096_);
  not _62417_ (_17099_, _34260_);
  nor _62418_ (_17100_, _17099_, _34221_);
  and _62419_ (_17101_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _62420_ (_17102_, _17101_, _34248_);
  or _62421_ (_17103_, _17102_, _17100_);
  or _62422_ (_17104_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _62423_ (_17105_, _17104_, _38997_);
  and _62424_ (_36882_[7], _17105_, _17103_);
  and _62425_ (_17106_, _34263_, _34247_);
  not _62426_ (_17107_, _17106_);
  nor _62427_ (_17108_, _17107_, _34221_);
  and _62428_ (_17109_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or _62429_ (_17110_, _17109_, _17108_);
  and _62430_ (_36883_[7], _17110_, _38997_);
  and _62431_ (_17111_, _34255_, _34247_);
  not _62432_ (_17112_, _17111_);
  nor _62433_ (_17113_, _17112_, _34221_);
  and _62434_ (_17114_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or _62435_ (_17115_, _17114_, _17113_);
  and _62436_ (_36884_[7], _17115_, _38997_);
  and _62437_ (_17116_, _34268_, _34247_);
  not _62438_ (_17117_, _17116_);
  nor _62439_ (_17118_, _17117_, _34221_);
  and _62440_ (_17119_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or _62441_ (_17120_, _17119_, _17118_);
  and _62442_ (_36885_[7], _17120_, _38997_);
  and _62443_ (_17121_, _34269_, _34247_);
  and _62444_ (_17122_, _17121_, _34318_);
  and _62445_ (_17123_, _34270_, _34266_);
  nand _62446_ (_17124_, _34261_, _34247_);
  or _62447_ (_17125_, _17124_, _17123_);
  or _62448_ (_17126_, _34255_, _34263_);
  or _62449_ (_17127_, _34268_, _17126_);
  and _62450_ (_17128_, _17127_, _34247_);
  or _62451_ (_17129_, _17128_, _17125_);
  and _62452_ (_17130_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  or _62453_ (_17131_, _17130_, _17122_);
  and _62454_ (_36886_[7], _17131_, _38997_);
  and _62455_ (_17132_, _34271_, _34247_);
  not _62456_ (_17133_, _17132_);
  nor _62457_ (_17134_, _17133_, _34221_);
  and _62458_ (_17135_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or _62459_ (_17136_, _17135_, _17134_);
  and _62460_ (_36887_[7], _17136_, _38997_);
  not _62461_ (_17137_, _34266_);
  or _62462_ (_17138_, _34279_, _17137_);
  and _62463_ (_17139_, _17138_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nand _62464_ (_17140_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor _62465_ (_17141_, _17140_, _34273_);
  nor _62466_ (_17142_, _34278_, _34221_);
  or _62467_ (_17143_, _17142_, _17141_);
  or _62468_ (_17144_, _17143_, _17139_);
  and _62469_ (_36888_[7], _17144_, _38997_);
  nand _62470_ (_17145_, _17095_, _34148_);
  or _62471_ (_17146_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _62472_ (_17147_, _17146_, _38997_);
  and _62473_ (_36881_[0], _17147_, _17145_);
  not _62474_ (_17148_, _17095_);
  or _62475_ (_17149_, _17148_, _34122_);
  or _62476_ (_17150_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _62477_ (_17151_, _17150_, _38997_);
  and _62478_ (_36881_[1], _17151_, _17149_);
  or _62479_ (_17152_, _17148_, _34089_);
  or _62480_ (_17153_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _62481_ (_17154_, _17153_, _38997_);
  and _62482_ (_36881_[2], _17154_, _17152_);
  nand _62483_ (_17155_, _17095_, _34052_);
  or _62484_ (_17156_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _62485_ (_17157_, _17156_, _38997_);
  and _62486_ (_36881_[3], _17157_, _17155_);
  nand _62487_ (_17158_, _17095_, _34017_);
  or _62488_ (_17159_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _62489_ (_17160_, _17159_, _38997_);
  and _62490_ (_36881_[4], _17160_, _17158_);
  or _62491_ (_17161_, _17148_, _33978_);
  or _62492_ (_17162_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _62493_ (_17163_, _17162_, _38997_);
  and _62494_ (_36881_[5], _17163_, _17161_);
  or _62495_ (_17164_, _17148_, _33942_);
  or _62496_ (_17165_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _62497_ (_17166_, _17165_, _38997_);
  and _62498_ (_36881_[6], _17166_, _17164_);
  and _62499_ (_17167_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _62500_ (_17168_, _34260_, _34149_);
  or _62501_ (_17169_, _17168_, _34248_);
  or _62502_ (_17170_, _17169_, _17167_);
  or _62503_ (_17171_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _62504_ (_17172_, _17171_, _38997_);
  and _62505_ (_36882_[0], _17172_, _17170_);
  and _62506_ (_17173_, _34260_, _34122_);
  and _62507_ (_17174_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or _62508_ (_17175_, _17174_, _34248_);
  or _62509_ (_17176_, _17175_, _17173_);
  or _62510_ (_17177_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _62511_ (_17178_, _17177_, _38997_);
  and _62512_ (_36882_[1], _17178_, _17176_);
  and _62513_ (_17179_, _34260_, _34089_);
  and _62514_ (_17180_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _62515_ (_17181_, _17180_, _34248_);
  or _62516_ (_17182_, _17181_, _17179_);
  or _62517_ (_17183_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _62518_ (_17184_, _17183_, _38997_);
  and _62519_ (_36882_[2], _17184_, _17182_);
  nor _62520_ (_17185_, _17099_, _34052_);
  and _62521_ (_17186_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _62522_ (_17187_, _17186_, _34248_);
  or _62523_ (_17188_, _17187_, _17185_);
  or _62524_ (_17189_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _62525_ (_17190_, _17189_, _38997_);
  and _62526_ (_36882_[3], _17190_, _17188_);
  nor _62527_ (_17191_, _17099_, _34017_);
  and _62528_ (_17192_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _62529_ (_17193_, _17192_, _34248_);
  or _62530_ (_17194_, _17193_, _17191_);
  or _62531_ (_17195_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _62532_ (_17196_, _17195_, _38997_);
  and _62533_ (_36882_[4], _17196_, _17194_);
  and _62534_ (_17197_, _34260_, _33978_);
  and _62535_ (_17198_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _62536_ (_17199_, _17198_, _34248_);
  or _62537_ (_17200_, _17199_, _17197_);
  or _62538_ (_17201_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _62539_ (_17202_, _17201_, _38997_);
  and _62540_ (_36882_[5], _17202_, _17200_);
  and _62541_ (_17203_, _34260_, _33942_);
  and _62542_ (_17204_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _62543_ (_17205_, _17204_, _34248_);
  or _62544_ (_17206_, _17205_, _17203_);
  or _62545_ (_17207_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _62546_ (_17208_, _17207_, _38997_);
  and _62547_ (_36882_[6], _17208_, _17206_);
  or _62548_ (_17209_, _34265_, _34248_);
  and _62549_ (_17210_, _17209_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nand _62550_ (_17211_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _62551_ (_17212_, _17211_, _34261_);
  and _62552_ (_17213_, _17106_, _34149_);
  or _62553_ (_17214_, _17213_, _17212_);
  or _62554_ (_17215_, _17214_, _17210_);
  and _62555_ (_36883_[0], _17215_, _38997_);
  and _62556_ (_17216_, _17106_, _34122_);
  and _62557_ (_17217_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or _62558_ (_17218_, _17217_, _17216_);
  and _62559_ (_36883_[1], _17218_, _38997_);
  and _62560_ (_17219_, _17106_, _34089_);
  and _62561_ (_17220_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or _62562_ (_17221_, _17220_, _17219_);
  and _62563_ (_36883_[2], _17221_, _38997_);
  nor _62564_ (_17222_, _17107_, _34052_);
  and _62565_ (_17223_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or _62566_ (_17224_, _17223_, _17222_);
  and _62567_ (_36883_[3], _17224_, _38997_);
  and _62568_ (_17225_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _62569_ (_17226_, _17107_, _34017_);
  or _62570_ (_17227_, _17226_, _17225_);
  and _62571_ (_36883_[4], _17227_, _38997_);
  and _62572_ (_17228_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _62573_ (_17229_, _17106_, _33978_);
  or _62574_ (_17230_, _17229_, _17228_);
  and _62575_ (_36883_[5], _17230_, _38997_);
  and _62576_ (_17231_, _17106_, _33942_);
  and _62577_ (_17232_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or _62578_ (_17233_, _17232_, _17231_);
  and _62579_ (_36883_[6], _17233_, _38997_);
  and _62580_ (_17234_, _17111_, _34149_);
  and _62581_ (_17235_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or _62582_ (_17236_, _17235_, _17234_);
  and _62583_ (_36884_[0], _17236_, _38997_);
  and _62584_ (_17237_, _17111_, _34122_);
  and _62585_ (_17238_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or _62586_ (_17239_, _17238_, _17237_);
  and _62587_ (_36884_[1], _17239_, _38997_);
  and _62588_ (_17240_, _17111_, _34089_);
  and _62589_ (_17241_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or _62590_ (_17242_, _17241_, _17240_);
  and _62591_ (_36884_[2], _17242_, _38997_);
  and _62592_ (_17243_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor _62593_ (_17244_, _17112_, _34052_);
  or _62594_ (_17245_, _17244_, _17243_);
  and _62595_ (_36884_[3], _17245_, _38997_);
  nor _62596_ (_17246_, _17112_, _34017_);
  and _62597_ (_17247_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or _62598_ (_17248_, _17247_, _17246_);
  and _62599_ (_36884_[4], _17248_, _38997_);
  and _62600_ (_17249_, _17111_, _33978_);
  and _62601_ (_17250_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or _62602_ (_17251_, _17250_, _17249_);
  and _62603_ (_36884_[5], _17251_, _38997_);
  and _62604_ (_17252_, _17111_, _33942_);
  and _62605_ (_17253_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or _62606_ (_17254_, _17253_, _17252_);
  and _62607_ (_36884_[6], _17254_, _38997_);
  and _62608_ (_17255_, _17116_, _34149_);
  and _62609_ (_17256_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  or _62610_ (_17257_, _17256_, _17255_);
  and _62611_ (_36885_[0], _17257_, _38997_);
  and _62612_ (_17258_, _17116_, _34122_);
  and _62613_ (_17259_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  or _62614_ (_17260_, _17259_, _17258_);
  and _62615_ (_36885_[1], _17260_, _38997_);
  and _62616_ (_17261_, _17116_, _34089_);
  and _62617_ (_17262_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or _62618_ (_17263_, _17262_, _17261_);
  and _62619_ (_36885_[2], _17263_, _38997_);
  nor _62620_ (_17264_, _17117_, _34052_);
  and _62621_ (_17265_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or _62622_ (_17266_, _17265_, _17264_);
  and _62623_ (_36885_[3], _17266_, _38997_);
  nor _62624_ (_17267_, _17117_, _34017_);
  and _62625_ (_17268_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or _62626_ (_17269_, _17268_, _17267_);
  and _62627_ (_36885_[4], _17269_, _38997_);
  and _62628_ (_17270_, _34268_, _33978_);
  and _62629_ (_17271_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or _62630_ (_17272_, _17271_, _17270_);
  or _62631_ (_17273_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _62632_ (_17274_, _17273_, _38997_);
  and _62633_ (_36885_[5], _17274_, _17272_);
  and _62634_ (_17275_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _62635_ (_17276_, _17116_, _33942_);
  or _62636_ (_17277_, _17276_, _17275_);
  and _62637_ (_36885_[6], _17277_, _38997_);
  and _62638_ (_17278_, _17121_, _34149_);
  and _62639_ (_17279_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  or _62640_ (_17280_, _17279_, _17278_);
  and _62641_ (_36886_[0], _17280_, _38997_);
  or _62642_ (_17281_, _17127_, _17125_);
  and _62643_ (_17282_, _17281_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _62644_ (_17283_, _17121_, _34122_);
  or _62645_ (_17284_, _17283_, _17282_);
  and _62646_ (_36886_[1], _17284_, _38997_);
  and _62647_ (_17285_, _17121_, _34089_);
  and _62648_ (_17286_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  or _62649_ (_17287_, _17286_, _17285_);
  and _62650_ (_36886_[2], _17287_, _38997_);
  and _62651_ (_17288_, _17121_, _34389_);
  and _62652_ (_17289_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or _62653_ (_17290_, _17289_, _17288_);
  and _62654_ (_36886_[3], _17290_, _38997_);
  and _62655_ (_17291_, _17121_, _34515_);
  and _62656_ (_17292_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  or _62657_ (_17293_, _17292_, _17291_);
  and _62658_ (_36886_[4], _17293_, _38997_);
  and _62659_ (_17294_, _17121_, _33978_);
  and _62660_ (_17295_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  or _62661_ (_17296_, _17295_, _17294_);
  and _62662_ (_36886_[5], _17296_, _38997_);
  and _62663_ (_17297_, _17121_, _33942_);
  and _62664_ (_17298_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or _62665_ (_17299_, _17298_, _17297_);
  and _62666_ (_36886_[6], _17299_, _38997_);
  and _62667_ (_17300_, _17132_, _34149_);
  and _62668_ (_17301_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  or _62669_ (_17302_, _17301_, _17300_);
  and _62670_ (_36887_[0], _17302_, _38997_);
  not _62671_ (_17303_, _34265_);
  or _62672_ (_17304_, _34275_, _17303_);
  and _62673_ (_17305_, _17304_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nand _62674_ (_17306_, _34270_, _34256_);
  and _62675_ (_17307_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _62676_ (_17308_, _17307_, _17306_);
  and _62677_ (_17309_, _17132_, _34122_);
  or _62678_ (_17310_, _17309_, _17308_);
  or _62679_ (_17311_, _17310_, _17305_);
  and _62680_ (_36887_[1], _17311_, _38997_);
  and _62681_ (_17312_, _17132_, _34089_);
  and _62682_ (_17313_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or _62683_ (_17314_, _17313_, _17312_);
  and _62684_ (_36887_[2], _17314_, _38997_);
  nor _62685_ (_17315_, _17133_, _34052_);
  and _62686_ (_17316_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or _62687_ (_17317_, _17316_, _17315_);
  and _62688_ (_36887_[3], _17317_, _38997_);
  nor _62689_ (_17318_, _17133_, _34017_);
  and _62690_ (_17319_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  or _62691_ (_17320_, _17319_, _17318_);
  and _62692_ (_36887_[4], _17320_, _38997_);
  and _62693_ (_17321_, _17132_, _33978_);
  and _62694_ (_17322_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or _62695_ (_17323_, _17322_, _17321_);
  and _62696_ (_36887_[5], _17323_, _38997_);
  and _62697_ (_17324_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and _62698_ (_17325_, _17132_, _33942_);
  or _62699_ (_17326_, _17325_, _17324_);
  and _62700_ (_36887_[6], _17326_, _38997_);
  and _62701_ (_17327_, _17138_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _62702_ (_17328_, _34267_, _34254_);
  and _62703_ (_17329_, _17328_, _34149_);
  not _62704_ (_17330_, _34273_);
  and _62705_ (_17331_, _17330_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or _62706_ (_17332_, _17331_, _17329_);
  and _62707_ (_17333_, _17332_, _34247_);
  or _62708_ (_17334_, _17333_, _17327_);
  and _62709_ (_36888_[0], _17334_, _38997_);
  and _62710_ (_17335_, _17138_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _62711_ (_17336_, _17328_, _34122_);
  and _62712_ (_17337_, _17330_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  or _62713_ (_17338_, _17337_, _17336_);
  and _62714_ (_17339_, _17338_, _34247_);
  or _62715_ (_17340_, _17339_, _17335_);
  and _62716_ (_36888_[1], _17340_, _38997_);
  and _62717_ (_17341_, _17138_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nand _62718_ (_17342_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _62719_ (_17343_, _17342_, _34273_);
  and _62720_ (_17344_, _34277_, _34089_);
  or _62721_ (_17345_, _17344_, _17343_);
  or _62722_ (_17346_, _17345_, _17341_);
  and _62723_ (_36888_[2], _17346_, _38997_);
  and _62724_ (_17347_, _17138_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nand _62725_ (_17348_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _62726_ (_17349_, _17348_, _34273_);
  nor _62727_ (_17350_, _34278_, _34052_);
  or _62728_ (_17351_, _17350_, _17349_);
  or _62729_ (_17352_, _17351_, _17347_);
  and _62730_ (_36888_[3], _17352_, _38997_);
  and _62731_ (_17353_, _17138_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nand _62732_ (_17354_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor _62733_ (_17355_, _17354_, _34273_);
  nor _62734_ (_17356_, _34278_, _34017_);
  or _62735_ (_17357_, _17356_, _17355_);
  or _62736_ (_17358_, _17357_, _17353_);
  and _62737_ (_36888_[4], _17358_, _38997_);
  and _62738_ (_17359_, _34279_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _62739_ (_17360_, _34277_, _33978_);
  nand _62740_ (_17361_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _62741_ (_17362_, _17361_, _34274_);
  or _62742_ (_17363_, _17362_, _17360_);
  or _62743_ (_17364_, _17363_, _17359_);
  and _62744_ (_36888_[5], _17364_, _38997_);
  and _62745_ (_17365_, _34277_, _33942_);
  and _62746_ (_17366_, _34278_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or _62747_ (_17367_, _17366_, _17365_);
  and _62748_ (_36888_[6], _17367_, _38997_);
  not _62749_ (_17368_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _62750_ (_17369_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and _62751_ (_17370_, _17369_, _17368_);
  and _62752_ (_17371_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _38997_);
  and _62753_ (_38985_, _17371_, _17370_);
  nor _62754_ (_17372_, _17370_, rst);
  nand _62755_ (_17373_, _17369_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or _62756_ (_17374_, _17369_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _62757_ (_17375_, _17374_, _17373_);
  and _62758_ (_38986_[3], _17375_, _17372_);
  not _62759_ (_17376_, _34691_);
  and _62760_ (_17377_, _34637_, _17376_);
  and _62761_ (_17378_, _34421_, _34346_);
  and _62762_ (_17379_, _17378_, _34699_);
  and _62763_ (_17380_, _17379_, _17377_);
  not _62764_ (_17381_, _34770_);
  nand _62765_ (_17382_, _14846_, _14832_);
  or _62766_ (_17383_, _14846_, _14832_);
  nand _62767_ (_17384_, _17383_, _17382_);
  or _62768_ (_17385_, _14869_, _14858_);
  nand _62769_ (_17386_, _14869_, _14858_);
  nand _62770_ (_17387_, _17386_, _17385_);
  nand _62771_ (_17388_, _17387_, _17384_);
  or _62772_ (_17389_, _17387_, _17384_);
  nand _62773_ (_17390_, _17389_, _17388_);
  or _62774_ (_17391_, _14894_, _14882_);
  nand _62775_ (_17392_, _14894_, _14882_);
  nand _62776_ (_17393_, _17392_, _17391_);
  or _62777_ (_17394_, _14904_, _14815_);
  nand _62778_ (_17395_, _14904_, _14815_);
  and _62779_ (_17396_, _17395_, _17394_);
  nand _62780_ (_17397_, _17396_, _17393_);
  or _62781_ (_17398_, _17396_, _17393_);
  nand _62782_ (_17399_, _17398_, _17397_);
  nand _62783_ (_17400_, _17399_, _17390_);
  or _62784_ (_17401_, _17399_, _17390_);
  and _62785_ (_17402_, _17401_, _17400_);
  or _62786_ (_17403_, _17402_, _17381_);
  and _62787_ (_17404_, _34579_, _34471_);
  or _62788_ (_17405_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _62789_ (_17406_, _17405_, _17404_);
  and _62790_ (_17407_, _17406_, _17403_);
  not _62791_ (_17408_, _34579_);
  nor _62792_ (_17409_, _17408_, _34471_);
  and _62793_ (_17410_, _17409_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _62794_ (_17411_, _17408_, _34471_);
  and _62795_ (_17412_, _17411_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _62796_ (_17413_, _17412_, _17410_);
  and _62797_ (_17414_, _17413_, _17381_);
  nor _62798_ (_17415_, _34579_, _34471_);
  nor _62799_ (_17416_, _34770_, _13513_);
  and _62800_ (_17417_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _62801_ (_17418_, _17417_, _17416_);
  and _62802_ (_17419_, _17418_, _17415_);
  and _62803_ (_17420_, _17409_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _62804_ (_17421_, _17411_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _62805_ (_17422_, _17421_, _17420_);
  and _62806_ (_17423_, _17422_, _34770_);
  or _62807_ (_17424_, _17423_, _17419_);
  or _62808_ (_17425_, _17424_, _17414_);
  or _62809_ (_17426_, _17425_, _17407_);
  and _62810_ (_17427_, _17426_, _17380_);
  not _62811_ (_17428_, _34421_);
  nor _62812_ (_17429_, _34637_, _17376_);
  nor _62813_ (_17430_, _34770_, _12205_);
  and _62814_ (_17431_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _62815_ (_17432_, _17431_, _17430_);
  and _62816_ (_17433_, _17432_, _17409_);
  and _62817_ (_17434_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _62818_ (_17435_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _62819_ (_17436_, _17435_, _17434_);
  and _62820_ (_17437_, _17436_, _17411_);
  nor _62821_ (_17438_, _34770_, _12203_);
  and _62822_ (_17439_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _62823_ (_17440_, _17439_, _17438_);
  and _62824_ (_17441_, _17440_, _17404_);
  or _62825_ (_17442_, _17441_, _17437_);
  and _62826_ (_17443_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _62827_ (_17444_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _62828_ (_17445_, _17444_, _17443_);
  and _62829_ (_17446_, _17445_, _17415_);
  or _62830_ (_17447_, _17446_, _17442_);
  or _62831_ (_17448_, _17447_, _17433_);
  and _62832_ (_17449_, _34699_, _34346_);
  and _62833_ (_17450_, _17449_, _17448_);
  and _62834_ (_17451_, _34529_, _34346_);
  and _62835_ (_17452_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _62836_ (_17453_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _62837_ (_17454_, _17453_, _17452_);
  and _62838_ (_17455_, _17454_, _17415_);
  and _62839_ (_17456_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _62840_ (_17457_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _62841_ (_17458_, _17457_, _17456_);
  and _62842_ (_17459_, _17458_, _17411_);
  nor _62843_ (_17460_, _34770_, _12174_);
  and _62844_ (_17461_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or _62845_ (_17462_, _17461_, _17460_);
  and _62846_ (_17463_, _17462_, _17404_);
  or _62847_ (_17464_, _17463_, _17459_);
  nor _62848_ (_17465_, _34770_, _12178_);
  and _62849_ (_17466_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _62850_ (_17467_, _17466_, _17465_);
  and _62851_ (_17468_, _17467_, _17409_);
  or _62852_ (_17469_, _17468_, _17464_);
  or _62853_ (_17470_, _17469_, _17455_);
  and _62854_ (_17471_, _17470_, _17451_);
  or _62855_ (_17472_, _17471_, _17450_);
  and _62856_ (_17473_, _17472_, _17429_);
  and _62857_ (_17474_, _34637_, _34691_);
  nor _62858_ (_17475_, _34770_, _11307_);
  and _62859_ (_17476_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _62860_ (_17477_, _17476_, _17475_);
  and _62861_ (_17478_, _17477_, _17409_);
  nor _62862_ (_17479_, _34770_, _10903_);
  and _62863_ (_17480_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _62864_ (_17481_, _17480_, _17479_);
  and _62865_ (_17482_, _17481_, _17411_);
  nor _62866_ (_17483_, _34770_, _10920_);
  and _62867_ (_17484_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _62868_ (_17485_, _17484_, _17483_);
  and _62869_ (_17486_, _17485_, _17404_);
  or _62870_ (_17487_, _17486_, _17482_);
  nor _62871_ (_17488_, _34770_, _11281_);
  and _62872_ (_17489_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _62873_ (_17490_, _17489_, _17488_);
  and _62874_ (_17491_, _17490_, _17415_);
  or _62875_ (_17492_, _17491_, _17487_);
  or _62876_ (_17493_, _17492_, _17478_);
  and _62877_ (_17494_, _17493_, _17449_);
  nor _62878_ (_17495_, _34770_, _11404_);
  and _62879_ (_17496_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _62880_ (_17497_, _17496_, _17495_);
  and _62881_ (_17498_, _17497_, _17411_);
  nor _62882_ (_17499_, _34770_, _11494_);
  and _62883_ (_17500_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _62884_ (_17501_, _17500_, _17499_);
  and _62885_ (_17502_, _17501_, _17404_);
  or _62886_ (_17503_, _17502_, _17498_);
  and _62887_ (_17504_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _62888_ (_17505_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _62889_ (_17506_, _17505_, _17504_);
  and _62890_ (_17507_, _17506_, _17415_);
  and _62891_ (_17508_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _62892_ (_17509_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _62893_ (_17510_, _17509_, _17508_);
  and _62894_ (_17511_, _17510_, _17409_);
  or _62895_ (_17512_, _17511_, _17507_);
  or _62896_ (_17513_, _17512_, _17503_);
  and _62897_ (_17514_, _17513_, _17451_);
  or _62898_ (_17515_, _17514_, _17494_);
  and _62899_ (_17516_, _17515_, _17474_);
  or _62900_ (_17517_, _17516_, _17473_);
  and _62901_ (_17518_, _17517_, _17428_);
  and _62902_ (_17519_, _17451_, _34421_);
  not _62903_ (_17520_, _34355_);
  not _62904_ (_17521_, _33433_);
  and _62905_ (_17522_, _33201_, _33381_);
  nor _62906_ (_17523_, _17522_, _33396_);
  and _62907_ (_17524_, _17523_, _17521_);
  and _62908_ (_17525_, _17524_, _17520_);
  and _62909_ (_17526_, _17525_, _15407_);
  nor _62910_ (_17527_, _33348_, _33323_);
  and _62911_ (_17528_, _33515_, _17527_);
  or _62912_ (_17529_, _15124_, _33430_);
  or _62913_ (_17530_, _17529_, _17528_);
  nor _62914_ (_17531_, _17530_, _15061_);
  and _62915_ (_17532_, _17531_, _15400_);
  and _62916_ (_17533_, _17532_, _17526_);
  and _62917_ (_17534_, _17533_, _33428_);
  nor _62918_ (_17535_, _17534_, _33477_);
  or _62919_ (_17536_, _17535_, p0_in[4]);
  not _62920_ (_17537_, _17535_);
  or _62921_ (_17538_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _62922_ (_17539_, _17538_, _17536_);
  and _62923_ (_17540_, _17539_, _17381_);
  or _62924_ (_17541_, _17535_, p0_in[0]);
  or _62925_ (_17542_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _62926_ (_17543_, _17542_, _17541_);
  and _62927_ (_17544_, _17543_, _34770_);
  or _62928_ (_17545_, _17544_, _17540_);
  and _62929_ (_17546_, _17545_, _17404_);
  or _62930_ (_17547_, _17535_, p0_in[7]);
  or _62931_ (_17548_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _62932_ (_17549_, _17548_, _17547_);
  and _62933_ (_17550_, _17549_, _17381_);
  or _62934_ (_17551_, _17535_, p0_in[3]);
  or _62935_ (_17552_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _62936_ (_17553_, _17552_, _17551_);
  and _62937_ (_17554_, _17553_, _34770_);
  or _62938_ (_17555_, _17554_, _17550_);
  and _62939_ (_17556_, _17555_, _17415_);
  or _62940_ (_17557_, _17556_, _17546_);
  or _62941_ (_17558_, _17535_, p0_in[5]);
  or _62942_ (_17559_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _62943_ (_17560_, _17559_, _17558_);
  and _62944_ (_17561_, _17560_, _17381_);
  or _62945_ (_17562_, _17535_, p0_in[1]);
  or _62946_ (_17563_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _62947_ (_17564_, _17563_, _17562_);
  and _62948_ (_17565_, _17564_, _34770_);
  or _62949_ (_17566_, _17565_, _17561_);
  and _62950_ (_17567_, _17566_, _17409_);
  nor _62951_ (_17568_, _17535_, p0_in[6]);
  and _62952_ (_17569_, _17535_, _13246_);
  nor _62953_ (_17570_, _17569_, _17568_);
  and _62954_ (_17571_, _17570_, _17381_);
  or _62955_ (_17572_, _17535_, p0_in[2]);
  nand _62956_ (_17573_, _17535_, _13190_);
  and _62957_ (_17574_, _17573_, _17572_);
  and _62958_ (_17575_, _17574_, _34770_);
  or _62959_ (_17576_, _17575_, _17571_);
  and _62960_ (_17577_, _17576_, _17411_);
  or _62961_ (_17578_, _17577_, _17567_);
  or _62962_ (_17579_, _17578_, _17557_);
  and _62963_ (_17580_, _17579_, _17519_);
  or _62964_ (_17581_, _17535_, p1_in[4]);
  or _62965_ (_17582_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _62966_ (_17583_, _17582_, _17581_);
  and _62967_ (_17584_, _17583_, _17381_);
  or _62968_ (_17585_, _17535_, p1_in[0]);
  or _62969_ (_17586_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _62970_ (_17587_, _17586_, _17585_);
  and _62971_ (_17588_, _17587_, _34770_);
  or _62972_ (_17589_, _17588_, _17584_);
  and _62973_ (_17590_, _17589_, _17404_);
  or _62974_ (_17591_, _17535_, p1_in[7]);
  or _62975_ (_17592_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _62976_ (_17593_, _17592_, _17591_);
  and _62977_ (_17594_, _17593_, _17381_);
  or _62978_ (_17595_, _17535_, p1_in[3]);
  or _62979_ (_17596_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _62980_ (_17597_, _17596_, _17595_);
  and _62981_ (_17598_, _17597_, _34770_);
  or _62982_ (_17599_, _17598_, _17594_);
  and _62983_ (_17600_, _17599_, _17415_);
  or _62984_ (_17601_, _17600_, _17590_);
  or _62985_ (_17602_, _17535_, p1_in[5]);
  or _62986_ (_17603_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _62987_ (_17604_, _17603_, _17602_);
  and _62988_ (_17605_, _17604_, _17381_);
  or _62989_ (_17606_, _17535_, p1_in[1]);
  or _62990_ (_17607_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _62991_ (_17608_, _17607_, _17606_);
  and _62992_ (_17609_, _17608_, _34770_);
  or _62993_ (_17610_, _17609_, _17605_);
  and _62994_ (_17611_, _17610_, _17409_);
  nor _62995_ (_17612_, _17535_, p1_in[6]);
  and _62996_ (_17613_, _17535_, _13330_);
  nor _62997_ (_17614_, _17613_, _17612_);
  and _62998_ (_17615_, _17614_, _17381_);
  or _62999_ (_17616_, _17535_, p1_in[2]);
  or _63000_ (_17617_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _63001_ (_17618_, _17617_, _17616_);
  and _63002_ (_17619_, _17618_, _34770_);
  or _63003_ (_17620_, _17619_, _17615_);
  and _63004_ (_17621_, _17620_, _17411_);
  or _63005_ (_17622_, _17621_, _17611_);
  or _63006_ (_17623_, _17622_, _17601_);
  and _63007_ (_17624_, _17623_, _17379_);
  or _63008_ (_17625_, _17624_, _17580_);
  and _63009_ (_17626_, _17625_, _17474_);
  nor _63010_ (_17627_, _34637_, _34691_);
  nor _63011_ (_17628_, _34770_, _14686_);
  and _63012_ (_17629_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _63013_ (_17630_, _17629_, _17628_);
  and _63014_ (_17631_, _17630_, _17415_);
  nor _63015_ (_17632_, _34770_, _14782_);
  and _63016_ (_17633_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _63017_ (_17634_, _17633_, _17632_);
  and _63018_ (_17635_, _17634_, _17411_);
  nor _63019_ (_17636_, _34770_, _14755_);
  and _63020_ (_17637_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or _63021_ (_17638_, _17637_, _17636_);
  and _63022_ (_17639_, _17638_, _17404_);
  or _63023_ (_17640_, _17639_, _17635_);
  nor _63024_ (_17641_, _34770_, _14769_);
  and _63025_ (_17642_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _63026_ (_17643_, _17642_, _17641_);
  and _63027_ (_17644_, _17643_, _17409_);
  or _63028_ (_17645_, _17644_, _17640_);
  or _63029_ (_17646_, _17645_, _17631_);
  and _63030_ (_17647_, _17646_, _17627_);
  or _63031_ (_17648_, _17535_, p3_in[7]);
  or _63032_ (_17649_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _63033_ (_17650_, _17649_, _17648_);
  and _63034_ (_17651_, _17650_, _17381_);
  or _63035_ (_17652_, _17535_, p3_in[3]);
  or _63036_ (_17653_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _63037_ (_17654_, _17653_, _17652_);
  and _63038_ (_17655_, _17654_, _34770_);
  or _63039_ (_17656_, _17655_, _17651_);
  and _63040_ (_17657_, _17656_, _17415_);
  nor _63041_ (_17658_, _17535_, p3_in[6]);
  and _63042_ (_17659_, _17535_, _13500_);
  nor _63043_ (_17660_, _17659_, _17658_);
  and _63044_ (_17661_, _17660_, _17381_);
  or _63045_ (_17662_, _17535_, p3_in[2]);
  or _63046_ (_17663_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _63047_ (_17664_, _17663_, _17662_);
  and _63048_ (_17665_, _17664_, _34770_);
  or _63049_ (_17666_, _17665_, _17661_);
  and _63050_ (_17667_, _17666_, _17411_);
  or _63051_ (_17668_, _17667_, _17657_);
  or _63052_ (_17669_, _17535_, p3_in[4]);
  or _63053_ (_17670_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _63054_ (_17671_, _17670_, _17669_);
  and _63055_ (_17672_, _17671_, _17381_);
  or _63056_ (_17673_, _17535_, p3_in[0]);
  or _63057_ (_17674_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _63058_ (_17675_, _17674_, _17673_);
  and _63059_ (_17676_, _17675_, _34770_);
  or _63060_ (_17677_, _17676_, _17672_);
  and _63061_ (_17678_, _17677_, _17404_);
  or _63062_ (_17679_, _17535_, p3_in[5]);
  or _63063_ (_17680_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _63064_ (_17681_, _17680_, _17679_);
  and _63065_ (_17682_, _17681_, _17381_);
  or _63066_ (_17683_, _17535_, p3_in[1]);
  or _63067_ (_17684_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _63068_ (_17685_, _17684_, _17683_);
  and _63069_ (_17686_, _17685_, _34770_);
  or _63070_ (_17687_, _17686_, _17682_);
  and _63071_ (_17688_, _17687_, _17409_);
  or _63072_ (_17689_, _17688_, _17678_);
  or _63073_ (_17690_, _17689_, _17668_);
  and _63074_ (_17691_, _17690_, _17429_);
  or _63075_ (_17692_, _17691_, _17647_);
  and _63076_ (_17693_, _17692_, _17379_);
  and _63077_ (_17694_, _15621_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _63078_ (_17695_, _17451_, _17377_);
  and _63079_ (_17696_, _17695_, _17428_);
  nand _63080_ (_17697_, _34691_, _34346_);
  or _63081_ (_17698_, _17697_, _34421_);
  nand _63082_ (_17699_, _17698_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nand _63083_ (_17700_, _34529_, _34637_);
  or _63084_ (_17701_, _17700_, _34691_);
  and _63085_ (_17702_, _17701_, _17378_);
  or _63086_ (_17703_, _17702_, _17699_);
  nor _63087_ (_17704_, _17703_, _17696_);
  and _63088_ (_17705_, _17627_, _17519_);
  nor _63089_ (_17706_, _34770_, _33984_);
  and _63090_ (_17707_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _63091_ (_17708_, _17707_, _17706_);
  and _63092_ (_17709_, _17708_, _17404_);
  nor _63093_ (_17710_, _34770_, _34193_);
  and _63094_ (_17711_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _63095_ (_17712_, _17711_, _17710_);
  and _63096_ (_17713_, _17712_, _17415_);
  or _63097_ (_17714_, _17713_, _17709_);
  nor _63098_ (_17715_, _34770_, _33773_);
  and _63099_ (_17716_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _63100_ (_17717_, _17716_, _17715_);
  and _63101_ (_17718_, _17717_, _17411_);
  nor _63102_ (_17719_, _34770_, _33948_);
  and _63103_ (_17720_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _63104_ (_17721_, _17720_, _17719_);
  and _63105_ (_17722_, _17721_, _17409_);
  or _63106_ (_17723_, _17722_, _17718_);
  or _63107_ (_17724_, _17723_, _17714_);
  and _63108_ (_17725_, _17724_, _17705_);
  or _63109_ (_17726_, _17725_, _17704_);
  nor _63110_ (_17727_, _34770_, _13097_);
  and _63111_ (_17728_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _63112_ (_17729_, _17728_, _17727_);
  and _63113_ (_17730_, _17729_, _17411_);
  nor _63114_ (_17731_, _34770_, _11000_);
  and _63115_ (_17732_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or _63116_ (_17733_, _17732_, _17731_);
  and _63117_ (_17734_, _17733_, _17404_);
  or _63118_ (_17735_, _17734_, _17730_);
  and _63119_ (_17736_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _63120_ (_17737_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _63121_ (_17738_, _17737_, _17736_);
  and _63122_ (_17739_, _17738_, _17415_);
  nor _63123_ (_17740_, _34770_, _10900_);
  and _63124_ (_17741_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _63125_ (_17742_, _17741_, _17740_);
  and _63126_ (_17743_, _17742_, _17409_);
  or _63127_ (_17744_, _17743_, _17739_);
  or _63128_ (_17745_, _17744_, _17735_);
  and _63129_ (_17746_, _17745_, _17696_);
  and _63130_ (_17747_, _17519_, _17429_);
  or _63131_ (_17748_, _17535_, p2_in[7]);
  or _63132_ (_17749_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _63133_ (_17750_, _17749_, _17748_);
  and _63134_ (_17751_, _17750_, _17381_);
  or _63135_ (_17752_, _17535_, p2_in[3]);
  or _63136_ (_17753_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _63137_ (_17754_, _17753_, _17752_);
  and _63138_ (_17755_, _17754_, _34770_);
  or _63139_ (_17756_, _17755_, _17751_);
  and _63140_ (_17757_, _17756_, _17415_);
  or _63141_ (_17758_, _17535_, p2_in[5]);
  or _63142_ (_17759_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _63143_ (_17760_, _17759_, _17758_);
  and _63144_ (_17761_, _17760_, _17381_);
  or _63145_ (_17762_, _17535_, p2_in[1]);
  or _63146_ (_17763_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _63147_ (_17764_, _17763_, _17762_);
  and _63148_ (_17765_, _17764_, _34770_);
  or _63149_ (_17766_, _17765_, _17761_);
  and _63150_ (_17767_, _17766_, _17409_);
  or _63151_ (_17768_, _17767_, _17757_);
  or _63152_ (_17769_, _17535_, p2_in[4]);
  or _63153_ (_17770_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _63154_ (_17771_, _17770_, _17769_);
  and _63155_ (_17772_, _17771_, _17381_);
  or _63156_ (_17773_, _17535_, p2_in[0]);
  or _63157_ (_17774_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _63158_ (_17775_, _17774_, _17773_);
  and _63159_ (_17776_, _17775_, _34770_);
  or _63160_ (_17777_, _17776_, _17772_);
  and _63161_ (_17778_, _17777_, _17404_);
  nor _63162_ (_17779_, _17535_, p2_in[6]);
  and _63163_ (_17780_, _17535_, _13415_);
  nor _63164_ (_17781_, _17780_, _17779_);
  and _63165_ (_17782_, _17781_, _17381_);
  or _63166_ (_17783_, _17535_, p2_in[2]);
  or _63167_ (_17784_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _63168_ (_17785_, _17784_, _17783_);
  and _63169_ (_17786_, _17785_, _34770_);
  or _63170_ (_17787_, _17786_, _17782_);
  and _63171_ (_17788_, _17787_, _17411_);
  or _63172_ (_17789_, _17788_, _17778_);
  or _63173_ (_17790_, _17789_, _17768_);
  and _63174_ (_17791_, _17790_, _17747_);
  or _63175_ (_17792_, _17791_, _17746_);
  or _63176_ (_17793_, _17792_, _17726_);
  or _63177_ (_17794_, _17793_, _17694_);
  or _63178_ (_17795_, _17794_, _17693_);
  or _63179_ (_17796_, _17795_, _17626_);
  or _63180_ (_17797_, _17796_, _17518_);
  or _63181_ (_17798_, _17797_, _17427_);
  and _63182_ (_17799_, _17705_, _14795_);
  nor _63183_ (_17800_, _17799_, _15630_);
  nand _63184_ (_17801_, _17694_, _35722_);
  and _63185_ (_17802_, _17801_, _17800_);
  and _63186_ (_17803_, _17802_, _17798_);
  nor _63187_ (_17804_, _34770_, _34221_);
  and _63188_ (_17805_, _34770_, _34389_);
  or _63189_ (_17806_, _17805_, _17804_);
  and _63190_ (_17807_, _17806_, _17415_);
  and _63191_ (_17808_, _17381_, _33942_);
  and _63192_ (_17809_, _34770_, _34089_);
  or _63193_ (_17810_, _17809_, _17808_);
  and _63194_ (_17811_, _17810_, _17411_);
  nor _63195_ (_17812_, _34770_, _34017_);
  and _63196_ (_17813_, _34770_, _34149_);
  or _63197_ (_17814_, _17813_, _17812_);
  and _63198_ (_17815_, _17814_, _17404_);
  or _63199_ (_17816_, _17815_, _17811_);
  and _63200_ (_17817_, _17381_, _33978_);
  and _63201_ (_17818_, _34770_, _34122_);
  or _63202_ (_17819_, _17818_, _17817_);
  and _63203_ (_17820_, _17819_, _17409_);
  or _63204_ (_17821_, _17820_, _17816_);
  nor _63205_ (_17822_, _17821_, _17807_);
  nor _63206_ (_17823_, _17822_, _17800_);
  or _63207_ (_17824_, _17823_, _17803_);
  and _63208_ (_38987_, _17824_, _38997_);
  and _63209_ (_17825_, _34770_, _34421_);
  and _63210_ (_17826_, _17474_, _17451_);
  and _63211_ (_17827_, _17826_, _17415_);
  and _63212_ (_17828_, _17827_, _17825_);
  and _63213_ (_17829_, _17828_, _14101_);
  and _63214_ (_17830_, _34699_, _34637_);
  nor _63215_ (_17831_, _34691_, _35178_);
  and _63216_ (_17832_, _17825_, _17404_);
  and _63217_ (_17833_, _17832_, _17831_);
  and _63218_ (_17834_, _17833_, _17830_);
  and _63219_ (_17835_, _17834_, _13518_);
  nor _63220_ (_17836_, _17835_, _17829_);
  nor _63221_ (_17837_, _17836_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _63222_ (_17838_, _17837_);
  not _63223_ (_17839_, _11084_);
  and _63224_ (_17840_, _17415_, _17381_);
  nor _63225_ (_17841_, _17840_, _17839_);
  and _63226_ (_17842_, _17841_, _15608_);
  nor _63227_ (_17843_, _34699_, _34637_);
  and _63228_ (_17844_, _17843_, _17833_);
  and _63229_ (_17845_, _17844_, _14819_);
  nor _63230_ (_17846_, _17845_, _17842_);
  and _63231_ (_17847_, _17846_, _15624_);
  and _63232_ (_17848_, _17847_, _17838_);
  and _63233_ (_17849_, _17825_, _17411_);
  and _63234_ (_17850_, _17849_, _17826_);
  and _63235_ (_17851_, _17850_, _14101_);
  or _63236_ (_17852_, _17851_, rst);
  nor _63237_ (_38988_, _17852_, _17848_);
  and _63238_ (_17853_, _34770_, _17428_);
  and _63239_ (_17854_, _17853_, _17404_);
  and _63240_ (_17855_, _17854_, _17826_);
  and _63241_ (_17856_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _63242_ (_17857_, _17853_, _17415_);
  and _63243_ (_17858_, _17857_, _17695_);
  and _63244_ (_17859_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or _63245_ (_17860_, _17859_, _17856_);
  and _63246_ (_17861_, _17840_, _34421_);
  and _63247_ (_17862_, _17449_, _17429_);
  and _63248_ (_17863_, _17862_, _17861_);
  and _63249_ (_17864_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _63250_ (_17865_, _17451_, _17429_);
  and _63251_ (_17866_, _17865_, _17854_);
  and _63252_ (_17867_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _63253_ (_17868_, _17867_, _17864_);
  or _63254_ (_17869_, _17868_, _17860_);
  and _63255_ (_17870_, _17854_, _17695_);
  and _63256_ (_17871_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor _63257_ (_17872_, _34770_, _34421_);
  and _63258_ (_17873_, _17872_, _17404_);
  and _63259_ (_17874_, _17873_, _17695_);
  and _63260_ (_17875_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _63261_ (_17876_, _17875_, _17871_);
  and _63262_ (_17877_, _17872_, _17409_);
  and _63263_ (_17878_, _17877_, _17695_);
  and _63264_ (_17879_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _63265_ (_17880_, _17853_, _17411_);
  and _63266_ (_17881_, _17880_, _17695_);
  and _63267_ (_17882_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _63268_ (_17883_, _17882_, _17879_);
  or _63269_ (_17884_, _17883_, _17876_);
  or _63270_ (_17885_, _17884_, _17869_);
  and _63271_ (_17886_, _17857_, _17826_);
  and _63272_ (_17887_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _63273_ (_17888_, _17853_, _17409_);
  and _63274_ (_17889_, _17888_, _17826_);
  and _63275_ (_17890_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or _63276_ (_17891_, _17890_, _17887_);
  and _63277_ (_17892_, _17877_, _17826_);
  and _63278_ (_17893_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _63279_ (_17894_, _17880_, _17826_);
  and _63280_ (_17895_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _63281_ (_17896_, _17895_, _17893_);
  or _63282_ (_17897_, _17896_, _17891_);
  and _63283_ (_17898_, _17474_, _17449_);
  and _63284_ (_17899_, _17898_, _17854_);
  and _63285_ (_17900_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _63286_ (_17901_, _17888_, _17898_);
  and _63287_ (_17902_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or _63288_ (_17903_, _17902_, _17900_);
  and _63289_ (_17904_, _17873_, _17826_);
  and _63290_ (_17905_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _63291_ (_17906_, _17861_, _17826_);
  and _63292_ (_17907_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _63293_ (_17908_, _17907_, _17905_);
  or _63294_ (_17909_, _17908_, _17903_);
  or _63295_ (_17910_, _17909_, _17897_);
  or _63296_ (_17911_, _17910_, _17885_);
  and _63297_ (_17912_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _63298_ (_17913_, _17825_, _17415_);
  and _63299_ (_17914_, _17913_, _17826_);
  and _63300_ (_17915_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _63301_ (_17916_, _17915_, _17912_);
  and _63302_ (_17917_, _17627_, _17449_);
  and _63303_ (_17918_, _17917_, _17832_);
  and _63304_ (_17919_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _63305_ (_17920_, _17825_, _17409_);
  and _63306_ (_17921_, _17920_, _17826_);
  and _63307_ (_17922_, _17921_, _34223_);
  or _63308_ (_17923_, _17922_, _17919_);
  or _63309_ (_17924_, _17923_, _17916_);
  and _63310_ (_17925_, _17865_, _17832_);
  and _63311_ (_17926_, _17925_, _17750_);
  and _63312_ (_17927_, _17862_, _17832_);
  and _63313_ (_17928_, _17927_, _17650_);
  or _63314_ (_17929_, _17928_, _17926_);
  and _63315_ (_17930_, _17832_, _17826_);
  and _63316_ (_17931_, _17930_, _17549_);
  and _63317_ (_17932_, _17898_, _17832_);
  and _63318_ (_17933_, _17932_, _17593_);
  or _63319_ (_17934_, _17933_, _17931_);
  or _63320_ (_17935_, _17934_, _17929_);
  or _63321_ (_17936_, _17935_, _17924_);
  and _63322_ (_17937_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _63323_ (_17938_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _63324_ (_17939_, _17938_, _17937_);
  or _63325_ (_17940_, _17939_, _17936_);
  or _63326_ (_17941_, _17940_, _17911_);
  and _63327_ (_17942_, _17941_, _17848_);
  nor _63328_ (_17943_, _17881_, _17878_);
  nand _63329_ (_17944_, _17696_, _17404_);
  and _63330_ (_17945_, _17944_, _17943_);
  nor _63331_ (_17946_, _17858_, _17855_);
  nor _63332_ (_17947_, _17866_, _17863_);
  and _63333_ (_17948_, _17947_, _17946_);
  and _63334_ (_17949_, _17948_, _17945_);
  nor _63335_ (_17950_, _17889_, _17886_);
  nor _63336_ (_17951_, _17894_, _17892_);
  and _63337_ (_17952_, _17951_, _17950_);
  nor _63338_ (_17953_, _17906_, _17904_);
  nor _63339_ (_17954_, _17901_, _17899_);
  and _63340_ (_17955_, _17954_, _17953_);
  and _63341_ (_17956_, _17955_, _17952_);
  and _63342_ (_17957_, _17956_, _17949_);
  not _63343_ (_17958_, _17832_);
  or _63344_ (_17959_, _17958_, _17697_);
  nor _63345_ (_17960_, _17914_, _17850_);
  nor _63346_ (_17961_, _17921_, _17918_);
  and _63347_ (_17962_, _17961_, _17960_);
  and _63348_ (_17963_, _17962_, _17959_);
  nor _63349_ (_17964_, _17844_, _17834_);
  and _63350_ (_17965_, _17964_, _17963_);
  nand _63351_ (_17966_, _17965_, _17957_);
  nand _63352_ (_17967_, _17966_, _17848_);
  and _63353_ (_17968_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or _63354_ (_17969_, _17968_, _17942_);
  or _63355_ (_17970_, _17969_, _17851_);
  nand _63356_ (_17971_, _17851_, _14098_);
  and _63357_ (_17972_, _17971_, _38997_);
  and _63358_ (_38989_[7], _17972_, _17970_);
  nor _63359_ (_38986_[0], \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or _63360_ (_17973_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor _63361_ (_17974_, _17369_, rst);
  and _63362_ (_38986_[1], _17974_, _17973_);
  nor _63363_ (_17975_, _17369_, _17368_);
  or _63364_ (_17976_, _17975_, _17370_);
  and _63365_ (_17977_, _17373_, _38997_);
  and _63366_ (_38986_[2], _17977_, _17976_);
  and _63367_ (_17978_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _63368_ (_17979_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or _63369_ (_17980_, _17979_, _17978_);
  and _63370_ (_17981_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _63371_ (_17982_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _63372_ (_17983_, _17982_, _17981_);
  or _63373_ (_17984_, _17983_, _17980_);
  and _63374_ (_17985_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _63375_ (_17986_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or _63376_ (_17987_, _17986_, _17985_);
  and _63377_ (_17988_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _63378_ (_17989_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _63379_ (_17990_, _17989_, _17988_);
  or _63380_ (_17991_, _17990_, _17987_);
  or _63381_ (_17992_, _17991_, _17984_);
  and _63382_ (_17993_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _63383_ (_17994_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _63384_ (_17995_, _17994_, _17993_);
  and _63385_ (_17996_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _63386_ (_17997_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or _63387_ (_17998_, _17997_, _17996_);
  or _63388_ (_17999_, _17998_, _17995_);
  and _63389_ (_18000_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _63390_ (_18001_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _63391_ (_18002_, _18001_, _18000_);
  and _63392_ (_18003_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and _63393_ (_18004_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _63394_ (_18005_, _18004_, _18003_);
  or _63395_ (_18006_, _18005_, _18002_);
  or _63396_ (_18007_, _18006_, _17999_);
  or _63397_ (_18008_, _18007_, _17992_);
  and _63398_ (_18009_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _63399_ (_18010_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _63400_ (_18011_, _18010_, _18009_);
  and _63401_ (_18012_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not _63402_ (_18013_, _17921_);
  nor _63403_ (_18014_, _18013_, _34466_);
  or _63404_ (_18015_, _18014_, _18012_);
  or _63405_ (_18016_, _18015_, _18011_);
  and _63406_ (_18017_, _17927_, _17675_);
  and _63407_ (_18018_, _17925_, _17775_);
  or _63408_ (_18019_, _18018_, _18017_);
  and _63409_ (_18020_, _17930_, _17543_);
  and _63410_ (_18021_, _17932_, _17587_);
  or _63411_ (_18022_, _18021_, _18020_);
  or _63412_ (_18023_, _18022_, _18019_);
  or _63413_ (_18024_, _18023_, _18016_);
  and _63414_ (_18025_, _17834_, _17402_);
  and _63415_ (_18026_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _63416_ (_18027_, _18026_, _18025_);
  or _63417_ (_18028_, _18027_, _18024_);
  or _63418_ (_18029_, _18028_, _18008_);
  and _63419_ (_18030_, _18029_, _17848_);
  and _63420_ (_18031_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or _63421_ (_18032_, _18031_, _17851_);
  or _63422_ (_18033_, _18032_, _18030_);
  nand _63423_ (_18034_, _17851_, _14224_);
  and _63424_ (_18035_, _18034_, _38997_);
  and _63425_ (_38989_[0], _18035_, _18033_);
  and _63426_ (_18036_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  not _63427_ (_18037_, _17851_);
  and _63428_ (_18038_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and _63429_ (_18039_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _63430_ (_18040_, _18039_, _18038_);
  and _63431_ (_18041_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _63432_ (_18042_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _63433_ (_18043_, _18042_, _18041_);
  or _63434_ (_18044_, _18043_, _18040_);
  and _63435_ (_18045_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _63436_ (_18046_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _63437_ (_18047_, _18046_, _18045_);
  and _63438_ (_18048_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _63439_ (_18049_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _63440_ (_18050_, _18049_, _18048_);
  or _63441_ (_18051_, _18050_, _18047_);
  or _63442_ (_18052_, _18051_, _18044_);
  and _63443_ (_18053_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _63444_ (_18054_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _63445_ (_18055_, _18054_, _18053_);
  and _63446_ (_18056_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _63447_ (_18057_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _63448_ (_18058_, _18057_, _18056_);
  or _63449_ (_18059_, _18058_, _18055_);
  and _63450_ (_18060_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _63451_ (_18061_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _63452_ (_18062_, _18061_, _18060_);
  and _63453_ (_18063_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _63454_ (_18064_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _63455_ (_18065_, _18064_, _18063_);
  or _63456_ (_18066_, _18065_, _18062_);
  or _63457_ (_18067_, _18066_, _18059_);
  or _63458_ (_18068_, _18067_, _18052_);
  and _63459_ (_18069_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _63460_ (_18070_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _63461_ (_18071_, _18070_, _18069_);
  and _63462_ (_18072_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _63463_ (_18073_, _17921_, _34558_);
  or _63464_ (_18074_, _18073_, _18072_);
  or _63465_ (_18075_, _18074_, _18071_);
  and _63466_ (_18076_, _17932_, _17608_);
  and _63467_ (_18077_, _17930_, _17564_);
  or _63468_ (_18078_, _18077_, _18076_);
  and _63469_ (_18079_, _17927_, _17685_);
  and _63470_ (_18080_, _17925_, _17764_);
  or _63471_ (_18081_, _18080_, _18079_);
  or _63472_ (_18082_, _18081_, _18078_);
  or _63473_ (_18083_, _18082_, _18075_);
  and _63474_ (_18084_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _63475_ (_18085_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _63476_ (_18086_, _18085_, _18084_);
  or _63477_ (_18087_, _18086_, _18083_);
  or _63478_ (_18088_, _18087_, _18068_);
  nand _63479_ (_18089_, _18088_, _17848_);
  nand _63480_ (_18090_, _18089_, _18037_);
  or _63481_ (_18091_, _18090_, _18036_);
  nand _63482_ (_18092_, _17851_, _14290_);
  and _63483_ (_18093_, _18092_, _38997_);
  and _63484_ (_38989_[1], _18093_, _18091_);
  and _63485_ (_18094_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _63486_ (_18095_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _63487_ (_18096_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _63488_ (_18097_, _18096_, _18095_);
  and _63489_ (_18098_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _63490_ (_18099_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _63491_ (_18100_, _18099_, _18098_);
  or _63492_ (_18101_, _18100_, _18097_);
  and _63493_ (_18102_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _63494_ (_18103_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _63495_ (_18104_, _18103_, _18102_);
  and _63496_ (_18105_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _63497_ (_18106_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _63498_ (_18107_, _18106_, _18105_);
  or _63499_ (_18108_, _18107_, _18104_);
  or _63500_ (_18109_, _18108_, _18101_);
  and _63501_ (_18110_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _63502_ (_18111_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or _63503_ (_18112_, _18111_, _18110_);
  and _63504_ (_18113_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _63505_ (_18114_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _63506_ (_18115_, _18114_, _18113_);
  or _63507_ (_18116_, _18115_, _18112_);
  and _63508_ (_18117_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and _63509_ (_18118_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _63510_ (_18119_, _18118_, _18117_);
  and _63511_ (_18120_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _63512_ (_18121_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _63513_ (_18122_, _18121_, _18120_);
  or _63514_ (_18123_, _18122_, _18119_);
  or _63515_ (_18124_, _18123_, _18116_);
  or _63516_ (_18125_, _18124_, _18109_);
  and _63517_ (_18126_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _63518_ (_18127_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _63519_ (_18128_, _18127_, _18126_);
  and _63520_ (_18129_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _63521_ (_18130_, _17921_, _34767_);
  or _63522_ (_18131_, _18130_, _18129_);
  or _63523_ (_18132_, _18131_, _18128_);
  and _63524_ (_18133_, _17925_, _17785_);
  and _63525_ (_18134_, _17927_, _17664_);
  or _63526_ (_18135_, _18134_, _18133_);
  and _63527_ (_18136_, _17930_, _17574_);
  and _63528_ (_18137_, _17932_, _17618_);
  or _63529_ (_18138_, _18137_, _18136_);
  or _63530_ (_18139_, _18138_, _18135_);
  or _63531_ (_18140_, _18139_, _18132_);
  and _63532_ (_18141_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _63533_ (_18142_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _63534_ (_18143_, _18142_, _18141_);
  or _63535_ (_18144_, _18143_, _18140_);
  or _63536_ (_18145_, _18144_, _18125_);
  and _63537_ (_18146_, _18145_, _17848_);
  or _63538_ (_18147_, _18146_, _17851_);
  or _63539_ (_18148_, _18147_, _18094_);
  nand _63540_ (_18149_, _17851_, _14356_);
  and _63541_ (_18150_, _18149_, _38997_);
  and _63542_ (_38989_[2], _18150_, _18148_);
  and _63543_ (_18151_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _63544_ (_18152_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _63545_ (_18153_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _63546_ (_18154_, _18153_, _18152_);
  and _63547_ (_18155_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _63548_ (_18156_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _63549_ (_18157_, _18156_, _18155_);
  or _63550_ (_18158_, _18157_, _18154_);
  and _63551_ (_18159_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _63552_ (_18160_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or _63553_ (_18161_, _18160_, _18159_);
  and _63554_ (_18162_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _63555_ (_18163_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _63556_ (_18164_, _18163_, _18162_);
  or _63557_ (_18165_, _18164_, _18161_);
  or _63558_ (_18166_, _18165_, _18158_);
  and _63559_ (_18167_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _63560_ (_18168_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or _63561_ (_18169_, _18168_, _18167_);
  and _63562_ (_18170_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _63563_ (_18171_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _63564_ (_18172_, _18171_, _18170_);
  or _63565_ (_18173_, _18172_, _18169_);
  and _63566_ (_18174_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and _63567_ (_18175_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _63568_ (_18176_, _18175_, _18174_);
  and _63569_ (_18177_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _63570_ (_18178_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or _63571_ (_18179_, _18178_, _18177_);
  or _63572_ (_18180_, _18179_, _18176_);
  or _63573_ (_18181_, _18180_, _18173_);
  or _63574_ (_18182_, _18181_, _18166_);
  and _63575_ (_18183_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _63576_ (_18184_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _63577_ (_18185_, _18184_, _18183_);
  and _63578_ (_18186_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _63579_ (_18187_, _17921_, _34401_);
  or _63580_ (_18188_, _18187_, _18186_);
  or _63581_ (_18189_, _18188_, _18185_);
  and _63582_ (_18190_, _17925_, _17754_);
  and _63583_ (_18191_, _17927_, _17654_);
  or _63584_ (_18192_, _18191_, _18190_);
  and _63585_ (_18193_, _17930_, _17553_);
  and _63586_ (_18194_, _17932_, _17597_);
  or _63587_ (_18195_, _18194_, _18193_);
  or _63588_ (_18196_, _18195_, _18192_);
  or _63589_ (_18197_, _18196_, _18189_);
  and _63590_ (_18198_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _63591_ (_18199_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _63592_ (_18200_, _18199_, _18198_);
  or _63593_ (_18201_, _18200_, _18197_);
  or _63594_ (_18202_, _18201_, _18182_);
  nand _63595_ (_18203_, _18202_, _17848_);
  nand _63596_ (_18204_, _18203_, _18037_);
  or _63597_ (_18205_, _18204_, _18151_);
  nand _63598_ (_18206_, _17851_, _14423_);
  and _63599_ (_18207_, _18206_, _38997_);
  and _63600_ (_38989_[3], _18207_, _18205_);
  and _63601_ (_18208_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _63602_ (_18209_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _63603_ (_18210_, _18209_, _18208_);
  and _63604_ (_18211_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _63605_ (_18212_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or _63606_ (_18213_, _18212_, _18211_);
  or _63607_ (_18214_, _18213_, _18210_);
  and _63608_ (_18215_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _63609_ (_18216_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _63610_ (_18217_, _18216_, _18215_);
  and _63611_ (_18218_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _63612_ (_18219_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _63613_ (_18220_, _18219_, _18218_);
  or _63614_ (_18221_, _18220_, _18217_);
  or _63615_ (_18222_, _18221_, _18214_);
  and _63616_ (_18223_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _63617_ (_18224_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _63618_ (_18225_, _18224_, _18223_);
  and _63619_ (_18226_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _63620_ (_18227_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  or _63621_ (_18228_, _18227_, _18226_);
  or _63622_ (_18229_, _18228_, _18225_);
  and _63623_ (_18230_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and _63624_ (_18231_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _63625_ (_18232_, _18231_, _18230_);
  and _63626_ (_18233_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _63627_ (_18234_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or _63628_ (_18235_, _18234_, _18233_);
  or _63629_ (_18236_, _18235_, _18232_);
  or _63630_ (_18237_, _18236_, _18229_);
  or _63631_ (_18238_, _18237_, _18222_);
  and _63632_ (_18239_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _63633_ (_18240_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _63634_ (_18241_, _18240_, _18239_);
  and _63635_ (_18242_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _63636_ (_18243_, _17921_, _34525_);
  or _63637_ (_18244_, _18243_, _18242_);
  or _63638_ (_18245_, _18244_, _18241_);
  and _63639_ (_18246_, _17930_, _17539_);
  and _63640_ (_18247_, _17932_, _17583_);
  or _63641_ (_18248_, _18247_, _18246_);
  and _63642_ (_18249_, _17927_, _17671_);
  and _63643_ (_18250_, _17925_, _17771_);
  or _63644_ (_18251_, _18250_, _18249_);
  or _63645_ (_18252_, _18251_, _18248_);
  or _63646_ (_18253_, _18252_, _18245_);
  and _63647_ (_18254_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _63648_ (_18255_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _63649_ (_18256_, _18255_, _18254_);
  or _63650_ (_18257_, _18256_, _18253_);
  or _63651_ (_18258_, _18257_, _18238_);
  and _63652_ (_18259_, _18258_, _17848_);
  and _63653_ (_18260_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or _63654_ (_18261_, _18260_, _18259_);
  or _63655_ (_18262_, _18261_, _17851_);
  nand _63656_ (_18263_, _17851_, _14495_);
  and _63657_ (_18264_, _18263_, _38997_);
  and _63658_ (_38989_[4], _18264_, _18262_);
  and _63659_ (_18265_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _63660_ (_18266_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _63661_ (_18267_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _63662_ (_18268_, _18267_, _18266_);
  and _63663_ (_18269_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _63664_ (_18270_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _63665_ (_18271_, _18270_, _18269_);
  or _63666_ (_18272_, _18271_, _18268_);
  and _63667_ (_18273_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _63668_ (_18274_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _63669_ (_18275_, _18274_, _18273_);
  and _63670_ (_18276_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _63671_ (_18277_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _63672_ (_18278_, _18277_, _18276_);
  or _63673_ (_18279_, _18278_, _18275_);
  or _63674_ (_18280_, _18279_, _18272_);
  and _63675_ (_18281_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _63676_ (_18282_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _63677_ (_18283_, _18282_, _18281_);
  and _63678_ (_18284_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _63679_ (_18285_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _63680_ (_18286_, _18285_, _18284_);
  or _63681_ (_18287_, _18286_, _18283_);
  and _63682_ (_18288_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _63683_ (_18289_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _63684_ (_18290_, _18289_, _18288_);
  and _63685_ (_18291_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _63686_ (_18292_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _63687_ (_18293_, _18292_, _18291_);
  or _63688_ (_18294_, _18293_, _18290_);
  or _63689_ (_18295_, _18294_, _18287_);
  or _63690_ (_18296_, _18295_, _18280_);
  and _63691_ (_18297_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _63692_ (_18298_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _63693_ (_18299_, _18298_, _18297_);
  and _63694_ (_18300_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor _63695_ (_18301_, _18013_, _34615_);
  or _63696_ (_18302_, _18301_, _18300_);
  or _63697_ (_18303_, _18302_, _18299_);
  and _63698_ (_18304_, _17932_, _17604_);
  and _63699_ (_18305_, _17930_, _17560_);
  or _63700_ (_18306_, _18305_, _18304_);
  and _63701_ (_18307_, _17927_, _17681_);
  and _63702_ (_18308_, _17925_, _17760_);
  or _63703_ (_18309_, _18308_, _18307_);
  or _63704_ (_18310_, _18309_, _18306_);
  or _63705_ (_18311_, _18310_, _18303_);
  and _63706_ (_18312_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _63707_ (_18313_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _63708_ (_18314_, _18313_, _18312_);
  or _63709_ (_18315_, _18314_, _18311_);
  or _63710_ (_18316_, _18315_, _18296_);
  nand _63711_ (_18317_, _18316_, _17848_);
  nand _63712_ (_18318_, _18317_, _18037_);
  or _63713_ (_18319_, _18318_, _18265_);
  nand _63714_ (_18320_, _17851_, _14570_);
  and _63715_ (_18321_, _18320_, _38997_);
  and _63716_ (_38989_[5], _18321_, _18319_);
  and _63717_ (_18322_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _63718_ (_18323_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nand _63719_ (_18324_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _63720_ (_18325_, _18324_, _18323_);
  nand _63721_ (_18326_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nand _63722_ (_18327_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _63723_ (_18328_, _18327_, _18326_);
  and _63724_ (_18329_, _18328_, _18325_);
  nand _63725_ (_18330_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _63726_ (_18331_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _63727_ (_18332_, _18331_, _18330_);
  nand _63728_ (_18333_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nand _63729_ (_18334_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _63730_ (_18335_, _18334_, _18333_);
  and _63731_ (_18336_, _18335_, _18332_);
  and _63732_ (_18337_, _18336_, _18329_);
  nand _63733_ (_18338_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand _63734_ (_18339_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _63735_ (_18340_, _18339_, _18338_);
  nand _63736_ (_18341_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _63737_ (_18342_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _63738_ (_18343_, _18342_, _18341_);
  and _63739_ (_18344_, _18343_, _18340_);
  nand _63740_ (_18345_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand _63741_ (_18346_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and _63742_ (_18347_, _18346_, _18345_);
  nand _63743_ (_18348_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  nand _63744_ (_18349_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _63745_ (_18350_, _18349_, _18348_);
  and _63746_ (_18351_, _18350_, _18347_);
  and _63747_ (_18352_, _18351_, _18344_);
  and _63748_ (_18353_, _18352_, _18337_);
  nand _63749_ (_18354_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nand _63750_ (_18355_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and _63751_ (_18356_, _18355_, _18354_);
  nand _63752_ (_18357_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or _63753_ (_18358_, _18013_, _34649_);
  and _63754_ (_18359_, _18358_, _18357_);
  and _63755_ (_18360_, _18359_, _18356_);
  nand _63756_ (_18361_, _17927_, _17660_);
  nand _63757_ (_18362_, _17925_, _17781_);
  and _63758_ (_18363_, _18362_, _18361_);
  nand _63759_ (_18364_, _17932_, _17614_);
  nand _63760_ (_18365_, _17930_, _17570_);
  and _63761_ (_18366_, _18365_, _18364_);
  and _63762_ (_18367_, _18366_, _18363_);
  and _63763_ (_18368_, _18367_, _18360_);
  nand _63764_ (_18369_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand _63765_ (_18370_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _63766_ (_18371_, _18370_, _18369_);
  and _63767_ (_18372_, _18371_, _18368_);
  nand _63768_ (_18373_, _18372_, _18353_);
  nand _63769_ (_18374_, _18373_, _17848_);
  nand _63770_ (_18375_, _18374_, _18037_);
  or _63771_ (_18376_, _18375_, _18322_);
  or _63772_ (_18377_, _18037_, _14632_);
  and _63773_ (_18378_, _18377_, _38997_);
  and _63774_ (_38989_[6], _18378_, _18376_);
  and _63775_ (_36924_, _34788_, _38997_);
  and _63776_ (_36925_[7], _35813_, _38997_);
  nor _63777_ (_36927_[2], _34770_, rst);
  and _63778_ (_36925_[0], _35732_, _38997_);
  and _63779_ (_36925_[1], _35748_, _38997_);
  and _63780_ (_36925_[2], _35757_, _38997_);
  and _63781_ (_36925_[3], _35767_, _38997_);
  and _63782_ (_36925_[4], _35778_, _38997_);
  and _63783_ (_36925_[5], _35791_, _38997_);
  and _63784_ (_36925_[6], _35802_, _38997_);
  nor _63785_ (_36927_[0], _34471_, rst);
  nor _63786_ (_36927_[1], _34579_, rst);
  nor _63787_ (_18379_, _16449_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _63788_ (_18380_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _63789_ (_18381_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _18380_);
  nor _63790_ (_18382_, _18381_, _18379_);
  nor _63791_ (_18383_, _16471_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _63792_ (_18384_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _18380_);
  nor _63793_ (_18385_, _18384_, _18383_);
  nor _63794_ (_18386_, _18385_, _18382_);
  and _63795_ (_18387_, _18386_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _63796_ (_18388_, _18385_, _18382_);
  and _63797_ (_18389_, _18388_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _63798_ (_18390_, _18389_, _18387_);
  not _63799_ (_18391_, _18382_);
  and _63800_ (_18392_, _18385_, _18391_);
  and _63801_ (_18393_, _18392_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _63802_ (_18394_, _18385_, _18391_);
  and _63803_ (_18395_, _18394_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _63804_ (_18396_, _18395_, _18393_);
  and _63805_ (_18397_, _18396_, _18390_);
  nor _63806_ (_18398_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _63807_ (_18399_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _18380_);
  nor _63808_ (_18400_, _18399_, _18398_);
  nor _63809_ (_18401_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _63810_ (_18402_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _18380_);
  nor _63811_ (_18403_, _18402_, _18401_);
  and _63812_ (_18404_, _18403_, _18400_);
  not _63813_ (_18405_, _18404_);
  nor _63814_ (_18406_, _18405_, _18397_);
  and _63815_ (_18407_, _18394_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _63816_ (_18408_, _18386_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _63817_ (_18409_, _18408_, _18407_);
  and _63818_ (_18410_, _18392_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _63819_ (_18411_, _18388_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _63820_ (_18412_, _18411_, _18410_);
  and _63821_ (_18413_, _18412_, _18409_);
  nor _63822_ (_18414_, _18403_, _18400_);
  not _63823_ (_18415_, _18414_);
  nor _63824_ (_18416_, _18415_, _18413_);
  nor _63825_ (_18417_, _18416_, _18406_);
  and _63826_ (_18418_, _18392_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _63827_ (_18419_, _18386_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _63828_ (_18420_, _18419_, _18418_);
  and _63829_ (_18421_, _18394_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _63830_ (_18422_, _18388_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _63831_ (_18423_, _18422_, _18421_);
  and _63832_ (_18424_, _18423_, _18420_);
  not _63833_ (_18425_, _18403_);
  and _63834_ (_18426_, _18425_, _18400_);
  not _63835_ (_18427_, _18426_);
  nor _63836_ (_18428_, _18427_, _18424_);
  and _63837_ (_18429_, _18388_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _63838_ (_18430_, _18386_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _63839_ (_18431_, _18430_, _18429_);
  and _63840_ (_18432_, _18392_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _63841_ (_18433_, _18394_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _63842_ (_18434_, _18433_, _18432_);
  and _63843_ (_18435_, _18434_, _18431_);
  not _63844_ (_18436_, _18400_);
  and _63845_ (_18437_, _18403_, _18436_);
  not _63846_ (_18438_, _18437_);
  nor _63847_ (_18439_, _18438_, _18435_);
  nor _63848_ (_18440_, _18439_, _18428_);
  and _63849_ (_18441_, _18440_, _18417_);
  and _63850_ (_18442_, _18441_, word_in[7]);
  not _63851_ (_18443_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand _63852_ (_18444_, _18400_, _18443_);
  or _63853_ (_18445_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _63854_ (_18446_, _18445_, _18444_);
  nor _63855_ (_18447_, _18403_, _18382_);
  and _63856_ (_18448_, _18447_, _18446_);
  or _63857_ (_18449_, _18448_, _18385_);
  and _63858_ (_18450_, _18403_, _18382_);
  not _63859_ (_18451_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _63860_ (_18452_, _18400_, _18451_);
  or _63861_ (_18453_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _63862_ (_18454_, _18453_, _18452_);
  and _63863_ (_18455_, _18454_, _18450_);
  and _63864_ (_18456_, _18425_, _18382_);
  not _63865_ (_18457_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand _63866_ (_18458_, _18400_, _18457_);
  or _63867_ (_18459_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _63868_ (_18460_, _18459_, _18458_);
  and _63869_ (_18461_, _18460_, _18456_);
  not _63870_ (_18462_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _63871_ (_18463_, _18400_, _18462_);
  or _63872_ (_18464_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _63873_ (_18465_, _18464_, _18463_);
  nor _63874_ (_18466_, _18425_, _18382_);
  and _63875_ (_18467_, _18466_, _18465_);
  or _63876_ (_18468_, _18467_, _18461_);
  or _63877_ (_18469_, _18468_, _18455_);
  or _63878_ (_18470_, _18469_, _18449_);
  not _63879_ (_18471_, _18385_);
  not _63880_ (_18472_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _63881_ (_18473_, _18400_, _18472_);
  or _63882_ (_18474_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _63883_ (_18475_, _18474_, _18473_);
  and _63884_ (_18476_, _18475_, _18447_);
  or _63885_ (_18477_, _18476_, _18471_);
  not _63886_ (_18478_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _63887_ (_18479_, _18400_, _18478_);
  or _63888_ (_18480_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _63889_ (_18481_, _18480_, _18479_);
  and _63890_ (_18482_, _18481_, _18456_);
  not _63891_ (_18483_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _63892_ (_18484_, _18400_, _18483_);
  or _63893_ (_18485_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _63894_ (_18486_, _18485_, _18484_);
  and _63895_ (_18487_, _18486_, _18450_);
  or _63896_ (_18488_, _18487_, _18482_);
  not _63897_ (_18489_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _63898_ (_18490_, _18400_, _18489_);
  or _63899_ (_18491_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _63900_ (_18492_, _18491_, _18490_);
  and _63901_ (_18493_, _18492_, _18466_);
  or _63902_ (_18494_, _18493_, _18488_);
  or _63903_ (_18495_, _18494_, _18477_);
  nand _63904_ (_18496_, _18495_, _18470_);
  nor _63905_ (_18497_, _18496_, _18441_);
  or _63906_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _18497_, _18442_);
  nor _63907_ (_18498_, _18404_, _18382_);
  and _63908_ (_18499_, _18404_, _18382_);
  nor _63909_ (_18500_, _18499_, _18498_);
  not _63910_ (_18501_, _18500_);
  nor _63911_ (_18502_, _18499_, _18471_);
  and _63912_ (_18503_, _18404_, _18394_);
  nor _63913_ (_18504_, _18503_, _18502_);
  and _63914_ (_18505_, _18504_, _18501_);
  and _63915_ (_18506_, _18505_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not _63916_ (_18507_, _18506_);
  not _63917_ (_18508_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nand _63918_ (_18509_, _18504_, _18508_);
  nor _63919_ (_18510_, _18504_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _63920_ (_18511_, _18510_, _18501_);
  and _63921_ (_18512_, _18511_, _18509_);
  nor _63922_ (_18513_, _18504_, _18500_);
  and _63923_ (_18514_, _18513_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _63924_ (_18515_, _18514_, _18512_);
  and _63925_ (_18516_, _18515_, _18507_);
  nor _63926_ (_18517_, _18516_, _18415_);
  and _63927_ (_18518_, _18505_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not _63928_ (_18519_, _18518_);
  not _63929_ (_18520_, _18504_);
  or _63930_ (_18521_, _18520_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _63931_ (_18522_, _18504_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _63932_ (_18523_, _18522_, _18501_);
  and _63933_ (_18524_, _18523_, _18521_);
  and _63934_ (_18525_, _18513_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _63935_ (_18526_, _18525_, _18524_);
  and _63936_ (_18527_, _18526_, _18519_);
  nor _63937_ (_18528_, _18527_, _18438_);
  nor _63938_ (_18529_, _18528_, _18517_);
  and _63939_ (_18530_, _18505_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not _63940_ (_18531_, _18530_);
  not _63941_ (_18532_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nand _63942_ (_18533_, _18504_, _18532_);
  nor _63943_ (_18534_, _18504_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _63944_ (_18535_, _18534_, _18501_);
  and _63945_ (_18536_, _18535_, _18533_);
  and _63946_ (_18537_, _18513_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _63947_ (_18538_, _18537_, _18536_);
  and _63948_ (_18539_, _18538_, _18531_);
  nor _63949_ (_18540_, _18539_, _18405_);
  and _63950_ (_18541_, _18505_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not _63951_ (_18542_, _18541_);
  not _63952_ (_18543_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nand _63953_ (_18544_, _18504_, _18543_);
  nor _63954_ (_18545_, _18504_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _63955_ (_18546_, _18545_, _18501_);
  and _63956_ (_18547_, _18546_, _18544_);
  and _63957_ (_18548_, _18513_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _63958_ (_18549_, _18548_, _18547_);
  and _63959_ (_18550_, _18549_, _18542_);
  nor _63960_ (_18551_, _18550_, _18427_);
  nor _63961_ (_18552_, _18551_, _18540_);
  and _63962_ (_18553_, _18552_, _18529_);
  and _63963_ (_18554_, _18553_, word_in[15]);
  or _63964_ (_18555_, _18414_, _18404_);
  not _63965_ (_18556_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand _63966_ (_18557_, _18400_, _18556_);
  or _63967_ (_18558_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _63968_ (_18559_, _18558_, _18557_);
  and _63969_ (_18560_, _18559_, _18555_);
  not _63970_ (_18561_, _18555_);
  and _63971_ (_18562_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nor _63972_ (_18563_, _18400_, _18462_);
  or _63973_ (_18564_, _18563_, _18562_);
  and _63974_ (_18565_, _18564_, _18561_);
  nor _63975_ (_18566_, _18565_, _18560_);
  nor _63976_ (_18567_, _18566_, _18500_);
  and _63977_ (_18568_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _63978_ (_18569_, _18400_, _18457_);
  or _63979_ (_18570_, _18569_, _18568_);
  and _63980_ (_18571_, _18570_, _18555_);
  not _63981_ (_18572_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand _63982_ (_18573_, _18400_, _18572_);
  or _63983_ (_18574_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _63984_ (_18575_, _18574_, _18573_);
  and _63985_ (_18576_, _18575_, _18561_);
  or _63986_ (_18577_, _18576_, _18571_);
  and _63987_ (_18578_, _18577_, _18500_);
  nor _63988_ (_18579_, _18578_, _18567_);
  nand _63989_ (_18580_, _18579_, _18504_);
  not _63990_ (_18581_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _63991_ (_18582_, _18400_, _18581_);
  or _63992_ (_18583_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _63993_ (_18584_, _18583_, _18582_);
  and _63994_ (_18585_, _18584_, _18555_);
  not _63995_ (_18586_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _63996_ (_18587_, _18400_, _18586_);
  or _63997_ (_18588_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _63998_ (_18589_, _18588_, _18587_);
  and _63999_ (_18590_, _18589_, _18561_);
  nor _64000_ (_18591_, _18590_, _18585_);
  nor _64001_ (_18592_, _18591_, _18500_);
  not _64002_ (_18593_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _64003_ (_18594_, _18400_, _18593_);
  or _64004_ (_18595_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _64005_ (_18596_, _18595_, _18594_);
  and _64006_ (_18597_, _18596_, _18555_);
  not _64007_ (_18598_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _64008_ (_18599_, _18400_, _18598_);
  or _64009_ (_18600_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _64010_ (_18601_, _18600_, _18599_);
  and _64011_ (_18602_, _18601_, _18561_);
  or _64012_ (_18603_, _18602_, _18597_);
  and _64013_ (_18604_, _18603_, _18500_);
  or _64014_ (_18605_, _18604_, _18592_);
  or _64015_ (_18606_, _18605_, _18504_);
  nand _64016_ (_18607_, _18606_, _18580_);
  nor _64017_ (_18608_, _18607_, _18553_);
  or _64018_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _18608_, _18554_);
  not _64019_ (_18609_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _64020_ (_18610_, _18450_, _18471_);
  not _64021_ (_18611_, _18610_);
  or _64022_ (_18612_, _18450_, _18471_);
  and _64023_ (_18613_, _18612_, _18611_);
  and _64024_ (_18614_, _18613_, _18609_);
  nor _64025_ (_18615_, _18450_, _18447_);
  not _64026_ (_18616_, _18615_);
  and _64027_ (_18617_, _18616_, _18613_);
  and _64028_ (_18618_, _18616_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _64029_ (_18619_, _18618_, _18617_);
  nor _64030_ (_18620_, _18619_, _18614_);
  and _64031_ (_18621_, _18613_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not _64032_ (_18622_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _64033_ (_18623_, _18613_, _18622_);
  nor _64034_ (_18624_, _18623_, _18621_);
  nor _64035_ (_18625_, _18624_, _18391_);
  nor _64036_ (_18626_, _18625_, _18620_);
  nor _64037_ (_18627_, _18626_, _18403_);
  and _64038_ (_18628_, _18613_, _18508_);
  not _64039_ (_18629_, _18466_);
  not _64040_ (_18630_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _64041_ (_18631_, _18385_, _18630_);
  nor _64042_ (_18632_, _18631_, _18629_);
  not _64043_ (_18633_, _18632_);
  nor _64044_ (_18634_, _18633_, _18628_);
  not _64045_ (_18635_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _64046_ (_18636_, _18613_, _18635_);
  and _64047_ (_18637_, _18450_, _18385_);
  and _64048_ (_18638_, _18450_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _64049_ (_18639_, _18638_, _18637_);
  nor _64050_ (_18640_, _18639_, _18636_);
  or _64051_ (_18641_, _18640_, _18436_);
  or _64052_ (_18642_, _18641_, _18634_);
  nor _64053_ (_18643_, _18642_, _18627_);
  not _64054_ (_18644_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _64055_ (_18645_, _18613_, _18644_);
  not _64056_ (_18646_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _64057_ (_18647_, _18615_, _18646_);
  nor _64058_ (_18648_, _18647_, _18617_);
  nor _64059_ (_18649_, _18648_, _18645_);
  and _64060_ (_18650_, _18613_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not _64061_ (_18651_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _64062_ (_18652_, _18613_, _18651_);
  nor _64063_ (_18653_, _18652_, _18650_);
  nor _64064_ (_18654_, _18653_, _18391_);
  nor _64065_ (_18655_, _18654_, _18649_);
  nor _64066_ (_18656_, _18655_, _18403_);
  not _64067_ (_18657_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _64068_ (_18658_, _18613_, _18657_);
  and _64069_ (_18659_, _18450_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _64070_ (_18660_, _18659_, _18637_);
  nor _64071_ (_18661_, _18660_, _18658_);
  and _64072_ (_18662_, _18613_, _18532_);
  not _64073_ (_18663_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _64074_ (_18664_, _18385_, _18663_);
  nor _64075_ (_18665_, _18664_, _18629_);
  not _64076_ (_18666_, _18665_);
  nor _64077_ (_18667_, _18666_, _18662_);
  or _64078_ (_18668_, _18667_, _18400_);
  or _64079_ (_18669_, _18668_, _18661_);
  nor _64080_ (_18670_, _18669_, _18656_);
  nor _64081_ (_18671_, _18670_, _18643_);
  not _64082_ (_18672_, _18671_);
  and _64083_ (_18673_, _18672_, word_in[23]);
  and _64084_ (_18674_, _18466_, _18460_);
  and _64085_ (_18675_, _18465_, _18447_);
  or _64086_ (_18676_, _18675_, _18674_);
  and _64087_ (_18677_, _18456_, _18454_);
  and _64088_ (_18678_, _18450_, _18446_);
  or _64089_ (_18679_, _18678_, _18677_);
  nor _64090_ (_18680_, _18679_, _18676_);
  nand _64091_ (_18681_, _18680_, _18613_);
  and _64092_ (_18682_, _18481_, _18466_);
  and _64093_ (_18683_, _18492_, _18447_);
  or _64094_ (_18684_, _18683_, _18682_);
  and _64095_ (_18685_, _18486_, _18456_);
  and _64096_ (_18686_, _18475_, _18450_);
  or _64097_ (_18687_, _18686_, _18685_);
  or _64098_ (_18688_, _18687_, _18684_);
  or _64099_ (_18689_, _18688_, _18613_);
  and _64100_ (_18690_, _18689_, _18681_);
  and _64101_ (_18691_, _18690_, _18671_);
  or _64102_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _18691_, _18673_);
  and _64103_ (_18692_, _18415_, _18382_);
  and _64104_ (_18693_, _18692_, _18385_);
  nor _64105_ (_18694_, _18692_, _18385_);
  nor _64106_ (_18695_, _18694_, _18693_);
  nor _64107_ (_18696_, _18695_, \oc8051_symbolic_cxrom1.regvalid [5]);
  not _64108_ (_18697_, _18696_);
  nor _64109_ (_18698_, _18415_, _18382_);
  nor _64110_ (_18699_, _18692_, _18698_);
  not _64111_ (_18700_, _18699_);
  nor _64112_ (_18701_, _18700_, _18631_);
  and _64113_ (_18702_, _18701_, _18697_);
  nor _64114_ (_18703_, _18695_, _18635_);
  and _64115_ (_18704_, _18695_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _64116_ (_18705_, _18704_, _18703_);
  nor _64117_ (_18706_, _18705_, _18699_);
  nor _64118_ (_18707_, _18706_, _18702_);
  nor _64119_ (_18708_, _18707_, _18438_);
  nor _64120_ (_18709_, _18695_, _18657_);
  and _64121_ (_18710_, _18695_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _64122_ (_18711_, _18710_, _18709_);
  nor _64123_ (_18712_, _18711_, _18699_);
  nor _64124_ (_18713_, _18695_, \oc8051_symbolic_cxrom1.regvalid [4]);
  not _64125_ (_18714_, _18713_);
  nor _64126_ (_18715_, _18700_, _18664_);
  and _64127_ (_18716_, _18715_, _18714_);
  nor _64128_ (_18717_, _18716_, _18712_);
  nor _64129_ (_18718_, _18717_, _18427_);
  nor _64130_ (_18719_, _18718_, _18708_);
  nor _64131_ (_18720_, _18695_, _18609_);
  and _64132_ (_18721_, _18695_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _64133_ (_18722_, _18721_, _18720_);
  nor _64134_ (_18723_, _18722_, _18699_);
  nand _64135_ (_18724_, _18695_, _18622_);
  nor _64136_ (_18725_, _18695_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _64137_ (_18726_, _18725_, _18700_);
  and _64138_ (_18727_, _18726_, _18724_);
  nor _64139_ (_18728_, _18727_, _18723_);
  nor _64140_ (_18729_, _18728_, _18415_);
  nor _64141_ (_18730_, _18695_, _18644_);
  and _64142_ (_18731_, _18695_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _64143_ (_18732_, _18731_, _18730_);
  nor _64144_ (_18733_, _18732_, _18699_);
  nand _64145_ (_18734_, _18695_, _18651_);
  nor _64146_ (_18735_, _18695_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _64147_ (_18736_, _18735_, _18700_);
  and _64148_ (_18737_, _18736_, _18734_);
  nor _64149_ (_18738_, _18737_, _18733_);
  nor _64150_ (_18739_, _18738_, _18405_);
  nor _64151_ (_18740_, _18739_, _18729_);
  and _64152_ (_18741_, _18740_, _18719_);
  and _64153_ (_18742_, _18601_, _18555_);
  and _64154_ (_18743_, _18596_, _18561_);
  or _64155_ (_18744_, _18743_, _18742_);
  and _64156_ (_18745_, _18744_, _18699_);
  and _64157_ (_18746_, _18589_, _18555_);
  and _64158_ (_18747_, _18584_, _18561_);
  nor _64159_ (_18748_, _18747_, _18746_);
  nor _64160_ (_18749_, _18748_, _18699_);
  or _64161_ (_18750_, _18749_, _18745_);
  and _64162_ (_18751_, _18750_, _18695_);
  not _64163_ (_18752_, _18695_);
  and _64164_ (_18753_, _18575_, _18555_);
  and _64165_ (_18754_, _18570_, _18561_);
  or _64166_ (_18755_, _18754_, _18753_);
  and _64167_ (_18756_, _18755_, _18699_);
  and _64168_ (_18757_, _18564_, _18555_);
  and _64169_ (_18758_, _18559_, _18561_);
  nor _64170_ (_18759_, _18758_, _18757_);
  nor _64171_ (_18760_, _18759_, _18699_);
  or _64172_ (_18761_, _18760_, _18756_);
  and _64173_ (_18762_, _18761_, _18752_);
  nor _64174_ (_18763_, _18762_, _18751_);
  nor _64175_ (_18764_, _18763_, _18741_);
  and _64176_ (_18765_, _18741_, word_in[31]);
  or _64177_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _18765_, _18764_);
  or _64178_ (_18766_, _18388_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _64179_ (_36729_[15], _18766_, _38997_);
  and _64180_ (_18767_, _18741_, _38997_);
  and _64181_ (_18768_, _18767_, word_in[31]);
  and _64182_ (_18769_, _18414_, _18388_);
  and _64183_ (_18770_, _18767_, _18769_);
  and _64184_ (_18771_, _18770_, _18768_);
  not _64185_ (_18772_, _18770_);
  and _64186_ (_18773_, _18643_, _38997_);
  and _64187_ (_18774_, _18773_, _18425_);
  not _64188_ (_18775_, _18613_);
  nor _64189_ (_18776_, _18671_, rst);
  and _64190_ (_18777_, _18776_, _18775_);
  and _64191_ (_18778_, _18777_, _18615_);
  and _64192_ (_18779_, _18778_, _18774_);
  and _64193_ (_18780_, _18553_, _38997_);
  and _64194_ (_18781_, _18780_, _18500_);
  and _64195_ (_18782_, _18781_, _18520_);
  and _64196_ (_18783_, _18782_, _18437_);
  and _64197_ (_18784_, _18499_, _18385_);
  and _64198_ (_18785_, _18441_, _38997_);
  and _64199_ (_18786_, _18785_, _18784_);
  and _64200_ (_18787_, _18786_, word_in[7]);
  nor _64201_ (_18788_, _18786_, _18483_);
  nor _64202_ (_18789_, _18788_, _18787_);
  nor _64203_ (_18790_, _18789_, _18783_);
  and _64204_ (_18791_, _18780_, word_in[15]);
  and _64205_ (_18792_, _18791_, _18783_);
  nor _64206_ (_18793_, _18792_, _18790_);
  nor _64207_ (_18794_, _18793_, _18779_);
  and _64208_ (_18795_, _18776_, word_in[23]);
  and _64209_ (_18796_, _18795_, _18779_);
  or _64210_ (_18797_, _18796_, _18794_);
  and _64211_ (_18798_, _18797_, _18772_);
  or _64212_ (_36785_, _18798_, _18771_);
  and _64213_ (_18799_, _18414_, _18386_);
  or _64214_ (_18800_, _18693_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _64215_ (_18801_, _18800_, _18799_);
  and _64216_ (_36858_, _18801_, _38997_);
  and _64217_ (_18802_, _18425_, _18386_);
  or _64218_ (_18803_, _18784_, _18802_);
  and _64219_ (_18804_, _18437_, _18388_);
  or _64220_ (_18805_, _18804_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _64221_ (_18806_, _18805_, _18803_);
  and _64222_ (_36729_[1], _18806_, _38997_);
  and _64223_ (_18807_, _18437_, _18386_);
  or _64224_ (_18808_, _18807_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _64225_ (_18809_, _18808_, _18803_);
  and _64226_ (_36729_[2], _18809_, _38997_);
  or _64227_ (_18810_, _18386_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _64228_ (_36729_[3], _18810_, _38997_);
  and _64229_ (_18811_, _18414_, _18394_);
  nand _64230_ (_18812_, _18694_, _18405_);
  and _64231_ (_18813_, _18812_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _64232_ (_18814_, _18813_, _18811_);
  nor _64233_ (_18815_, _18814_, _18386_);
  and _64234_ (_18816_, _18404_, _18386_);
  and _64235_ (_18817_, _18426_, _18386_);
  and _64236_ (_18818_, _18799_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _64237_ (_18819_, _18818_, _18817_);
  or _64238_ (_18820_, _18819_, _18816_);
  or _64239_ (_18821_, _18820_, _18807_);
  or _64240_ (_18822_, _18821_, _18815_);
  and _64241_ (_36729_[4], _18822_, _38997_);
  nor _64242_ (_18823_, _18784_, _18386_);
  and _64243_ (_18824_, _18426_, _18394_);
  or _64244_ (_18825_, _18824_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor _64245_ (_18826_, _18694_, _18784_);
  and _64246_ (_18827_, _18826_, _18825_);
  nor _64247_ (_18828_, _18385_, _18508_);
  and _64248_ (_18829_, _18466_, _18828_);
  or _64249_ (_18830_, _18829_, _18811_);
  or _64250_ (_18831_, _18830_, _18827_);
  and _64251_ (_18832_, _18831_, _18823_);
  and _64252_ (_18833_, _18817_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _64253_ (_18834_, _18833_, _18807_);
  and _64254_ (_18835_, _18698_, _18828_);
  and _64255_ (_18836_, _18825_, _18784_);
  or _64256_ (_18837_, _18836_, _18835_);
  or _64257_ (_18838_, _18837_, _18834_);
  or _64258_ (_18839_, _18838_, _18816_);
  or _64259_ (_18840_, _18839_, _18832_);
  and _64260_ (_36729_[5], _18840_, _38997_);
  not _64261_ (_18841_, _18824_);
  nor _64262_ (_18842_, _18816_, _18811_);
  nand _64263_ (_18843_, _18842_, _18841_);
  and _64264_ (_18844_, _18405_, _18386_);
  and _64265_ (_18845_, _18844_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _64266_ (_18846_, _18450_, _18385_);
  and _64267_ (_18847_, _18437_, _18394_);
  or _64268_ (_18848_, _18400_, _18385_);
  nor _64269_ (_18849_, _18386_, _18543_);
  and _64270_ (_18850_, _18849_, _18848_);
  or _64271_ (_18851_, _18850_, _18847_);
  and _64272_ (_18852_, _18851_, _18846_);
  or _64273_ (_18853_, _18852_, _18845_);
  or _64274_ (_18854_, _18853_, _18843_);
  and _64275_ (_36729_[6], _18854_, _38997_);
  or _64276_ (_18855_, _18502_, _18610_);
  and _64277_ (_18856_, _18425_, _18395_);
  nand _64278_ (_18857_, _18438_, _18394_);
  and _64279_ (_18858_, _18857_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _64280_ (_18859_, _18858_, _18856_);
  and _64281_ (_18860_, _18859_, _18502_);
  or _64282_ (_18861_, _18856_, _18610_);
  or _64283_ (_18862_, _18861_, _18860_);
  and _64284_ (_18863_, _18862_, _18855_);
  and _64285_ (_18864_, _18859_, _18784_);
  and _64286_ (_18865_, _18807_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _64287_ (_18866_, _18816_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _64288_ (_18867_, _18802_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _64289_ (_18868_, _18867_, _18811_);
  or _64290_ (_18869_, _18868_, _18866_);
  or _64291_ (_18870_, _18869_, _18865_);
  or _64292_ (_18871_, _18870_, _18864_);
  or _64293_ (_18872_, _18871_, _18824_);
  or _64294_ (_18873_, _18872_, _18863_);
  and _64295_ (_36729_[7], _18873_, _38997_);
  and _64296_ (_18874_, _18561_, _18386_);
  not _64297_ (_18875_, _18698_);
  nand _64298_ (_18876_, _18842_, _18875_);
  or _64299_ (_18877_, _18876_, _18874_);
  and _64300_ (_18878_, _18877_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _64301_ (_18879_, _18400_, _18394_);
  or _64302_ (_18880_, _18698_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _64303_ (_18881_, _18880_, _18385_);
  or _64304_ (_18882_, _18881_, _18879_);
  or _64305_ (_18883_, _18882_, _18847_);
  or _64306_ (_18884_, _18883_, _18878_);
  and _64307_ (_36729_[8], _18884_, _38997_);
  not _64308_ (_18885_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _64309_ (_18886_, _18846_, _18885_);
  and _64310_ (_18887_, _18846_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _64311_ (_18888_, _18426_, _18392_);
  or _64312_ (_18889_, _18888_, _18698_);
  or _64313_ (_18890_, _18889_, _18887_);
  and _64314_ (_18891_, _18890_, _18385_);
  or _64315_ (_18892_, _18891_, _18610_);
  or _64316_ (_18893_, _18892_, _18886_);
  and _64317_ (_36729_[9], _18893_, _38997_);
  and _64318_ (_18894_, _18615_, _18385_);
  or _64319_ (_18895_, _18894_, _18804_);
  or _64320_ (_18896_, _18895_, _18784_);
  nand _64321_ (_18897_, _18561_, _18394_);
  nand _64322_ (_18898_, _18842_, _18897_);
  and _64323_ (_18899_, _18898_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _64324_ (_18900_, _18437_, _18392_);
  and _64325_ (_18901_, _18799_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _64326_ (_18902_, _18874_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _64327_ (_18903_, _18902_, _18901_);
  or _64328_ (_18904_, _18903_, _18900_);
  and _64329_ (_18905_, _18698_, _18385_);
  or _64330_ (_18906_, _18905_, _18503_);
  and _64331_ (_18907_, _18906_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _64332_ (_18908_, _18498_, _18471_);
  or _64333_ (_18909_, _18908_, _18888_);
  and _64334_ (_18910_, _18909_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _64335_ (_18911_, _18910_, _18907_);
  or _64336_ (_18912_, _18911_, _18904_);
  or _64337_ (_18913_, _18912_, _18899_);
  and _64338_ (_18914_, _18913_, _18896_);
  nor _64339_ (_18915_, _18824_, _18807_);
  and _64340_ (_18916_, _18915_, _18842_);
  nor _64341_ (_18917_, _18916_, _18646_);
  and _64342_ (_18918_, _18847_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _64343_ (_18919_, _18802_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _64344_ (_18920_, _18919_, _18503_);
  or _64345_ (_18921_, _18920_, _18918_);
  or _64346_ (_18922_, _18921_, _18917_);
  or _64347_ (_18923_, _18922_, _18888_);
  or _64348_ (_18924_, _18923_, _18905_);
  or _64349_ (_18925_, _18924_, _18914_);
  and _64350_ (_36729_[10], _18925_, _38997_);
  and _64351_ (_18926_, _18404_, _18392_);
  or _64352_ (_18927_, _18926_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _64353_ (_18928_, _18500_, _18385_);
  and _64354_ (_18929_, _18928_, _18927_);
  or _64355_ (_18930_, _18811_, _18824_);
  and _64356_ (_18931_, _18930_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _64357_ (_18932_, _18847_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _64358_ (_18933_, _18932_, _18931_);
  and _64359_ (_18934_, _18816_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _64360_ (_18935_, _18934_, _18933_);
  and _64361_ (_18936_, _18905_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _64362_ (_18937_, _18874_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _64363_ (_18938_, _18937_, _18936_);
  and _64364_ (_18939_, _18888_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _64365_ (_18940_, _18503_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _64366_ (_18941_, _18940_, _18900_);
  or _64367_ (_18942_, _18941_, _18939_);
  or _64368_ (_18943_, _18942_, _18938_);
  or _64369_ (_18944_, _18943_, _18935_);
  or _64370_ (_18945_, _18944_, _18929_);
  and _64371_ (_18946_, _18945_, _18895_);
  or _64372_ (_18947_, _18937_, _18940_);
  or _64373_ (_18948_, _18947_, _18935_);
  and _64374_ (_18949_, _18799_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _64375_ (_18950_, _18784_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _64376_ (_18951_, _18950_, _18949_);
  or _64377_ (_18952_, _18951_, _18905_);
  or _64378_ (_18953_, _18952_, _18948_);
  or _64379_ (_18954_, _18953_, _18888_);
  or _64380_ (_18955_, _18954_, _18946_);
  and _64381_ (_36729_[11], _18955_, _38997_);
  and _64382_ (_18956_, _18693_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _64383_ (_18957_, _18415_, _18394_);
  and _64384_ (_18958_, _18957_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _64385_ (_18959_, _18816_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _64386_ (_18960_, _18811_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _64387_ (_18961_, _18698_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _64388_ (_18962_, _18961_, _18888_);
  or _64389_ (_18963_, _18962_, _18960_);
  or _64390_ (_18964_, _18963_, _18959_);
  and _64391_ (_18965_, _18874_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _64392_ (_18966_, _18426_, _18388_);
  not _64393_ (_18967_, _18966_);
  and _64394_ (_18968_, _18894_, _18967_);
  or _64395_ (_18969_, _18968_, _18965_);
  or _64396_ (_18970_, _18969_, _18964_);
  or _64397_ (_18971_, _18970_, _18958_);
  or _64398_ (_18972_, _18971_, _18956_);
  and _64399_ (_36729_[12], _18972_, _38997_);
  or _64400_ (_18973_, _18894_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _64401_ (_36729_[13], _18973_, _38997_);
  or _64402_ (_18974_, _18928_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _64403_ (_36729_[14], _18974_, _38997_);
  and _64404_ (_18975_, _18767_, _18699_);
  and _64405_ (_18976_, _18767_, _18695_);
  nor _64406_ (_18977_, _18976_, _18975_);
  and _64407_ (_18978_, _18977_, _18426_);
  and _64408_ (_18979_, _18978_, _18767_);
  and _64409_ (_18980_, _18776_, _18425_);
  nor _64410_ (_18981_, _18980_, _18773_);
  and _64411_ (_18982_, _18981_, _18776_);
  and _64412_ (_18983_, _18982_, _18617_);
  and _64413_ (_18984_, _18780_, _18784_);
  not _64414_ (_18985_, _18984_);
  or _64415_ (_18986_, _18985_, word_in[8]);
  not _64416_ (_18987_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _64417_ (_18988_, _18785_, _18799_);
  nor _64418_ (_18989_, _18988_, _18987_);
  and _64419_ (_18990_, _18988_, word_in[0]);
  or _64420_ (_18991_, _18990_, _18989_);
  or _64421_ (_18992_, _18991_, _18984_);
  and _64422_ (_18993_, _18992_, _18986_);
  or _64423_ (_18994_, _18993_, _18983_);
  not _64424_ (_18995_, _18983_);
  or _64425_ (_18996_, _18995_, word_in[16]);
  and _64426_ (_18997_, _18996_, _18994_);
  or _64427_ (_18998_, _18997_, _18979_);
  not _64428_ (_18999_, _18979_);
  or _64429_ (_19000_, _18999_, word_in[24]);
  and _64430_ (_36730_, _19000_, _18998_);
  and _64431_ (_19001_, _18780_, word_in[9]);
  and _64432_ (_19002_, _19001_, _18984_);
  not _64433_ (_19003_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _64434_ (_19004_, _18988_, _19003_);
  and _64435_ (_19005_, _18988_, word_in[1]);
  nor _64436_ (_19006_, _19005_, _19004_);
  nor _64437_ (_19007_, _19006_, _18984_);
  or _64438_ (_19008_, _19007_, _19002_);
  or _64439_ (_19009_, _19008_, _18983_);
  or _64440_ (_19010_, _18995_, word_in[17]);
  and _64441_ (_19011_, _19010_, _19009_);
  or _64442_ (_19012_, _19011_, _18979_);
  or _64443_ (_19013_, _18999_, word_in[25]);
  and _64444_ (_36731_, _19013_, _19012_);
  or _64445_ (_19014_, _18985_, word_in[10]);
  and _64446_ (_19015_, _18988_, word_in[2]);
  not _64447_ (_19016_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _64448_ (_19017_, _18988_, _19016_);
  or _64449_ (_19018_, _19017_, _19015_);
  or _64450_ (_19019_, _19018_, _18984_);
  and _64451_ (_19020_, _19019_, _19014_);
  or _64452_ (_19021_, _19020_, _18983_);
  or _64453_ (_19022_, _18995_, word_in[18]);
  and _64454_ (_19023_, _19022_, _19021_);
  or _64455_ (_19024_, _19023_, _18979_);
  or _64456_ (_19025_, _18999_, word_in[26]);
  and _64457_ (_36732_, _19025_, _19024_);
  or _64458_ (_19026_, _18985_, word_in[11]);
  not _64459_ (_19027_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _64460_ (_19028_, _18988_, _19027_);
  and _64461_ (_19029_, _18988_, word_in[3]);
  or _64462_ (_19030_, _19029_, _19028_);
  or _64463_ (_19031_, _19030_, _18984_);
  and _64464_ (_19032_, _19031_, _19026_);
  or _64465_ (_19033_, _19032_, _18983_);
  or _64466_ (_19034_, _18995_, word_in[19]);
  and _64467_ (_19035_, _19034_, _19033_);
  or _64468_ (_19036_, _19035_, _18979_);
  or _64469_ (_19037_, _18999_, word_in[27]);
  and _64470_ (_36733_, _19037_, _19036_);
  and _64471_ (_19038_, _18767_, word_in[28]);
  and _64472_ (_19039_, _19038_, _18978_);
  or _64473_ (_19040_, _18995_, word_in[20]);
  or _64474_ (_19041_, _18985_, word_in[12]);
  not _64475_ (_19042_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _64476_ (_19043_, _18988_, _19042_);
  and _64477_ (_19044_, _18988_, word_in[4]);
  or _64478_ (_19045_, _19044_, _19043_);
  or _64479_ (_19046_, _19045_, _18984_);
  and _64480_ (_19047_, _19046_, _19041_);
  or _64481_ (_19048_, _19047_, _18983_);
  and _64482_ (_19049_, _19048_, _18999_);
  and _64483_ (_19050_, _19049_, _19040_);
  or _64484_ (_36734_, _19050_, _19039_);
  or _64485_ (_19051_, _18995_, word_in[21]);
  or _64486_ (_19052_, _18985_, word_in[13]);
  and _64487_ (_19053_, _18988_, word_in[5]);
  not _64488_ (_19054_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _64489_ (_19055_, _18988_, _19054_);
  or _64490_ (_19056_, _19055_, _19053_);
  or _64491_ (_19057_, _19056_, _18984_);
  and _64492_ (_19058_, _19057_, _19052_);
  or _64493_ (_19059_, _19058_, _18983_);
  and _64494_ (_19060_, _19059_, _18999_);
  and _64495_ (_19061_, _19060_, _19051_);
  and _64496_ (_19062_, _18979_, word_in[29]);
  or _64497_ (_36735_, _19062_, _19061_);
  or _64498_ (_19063_, _18985_, word_in[14]);
  and _64499_ (_19064_, _18988_, word_in[6]);
  not _64500_ (_19065_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _64501_ (_19066_, _18988_, _19065_);
  or _64502_ (_19067_, _19066_, _19064_);
  or _64503_ (_19068_, _19067_, _18984_);
  and _64504_ (_19069_, _19068_, _19063_);
  or _64505_ (_19070_, _19069_, _18983_);
  or _64506_ (_19071_, _18995_, word_in[22]);
  and _64507_ (_19072_, _19071_, _19070_);
  or _64508_ (_19073_, _19072_, _18979_);
  or _64509_ (_19074_, _18999_, word_in[30]);
  and _64510_ (_36736_, _19074_, _19073_);
  or _64511_ (_19075_, _18985_, word_in[15]);
  and _64512_ (_19076_, _18988_, word_in[7]);
  nor _64513_ (_19077_, _18988_, _18556_);
  or _64514_ (_19078_, _19077_, _19076_);
  or _64515_ (_19079_, _19078_, _18984_);
  and _64516_ (_19080_, _19079_, _19075_);
  or _64517_ (_19081_, _19080_, _18983_);
  or _64518_ (_19082_, _18995_, word_in[23]);
  and _64519_ (_19083_, _19082_, _19081_);
  or _64520_ (_19084_, _19083_, _18979_);
  or _64521_ (_19085_, _18999_, word_in[31]);
  and _64522_ (_36737_, _19085_, _19084_);
  and _64523_ (_19086_, _18767_, _18437_);
  and _64524_ (_19087_, _19086_, _18977_);
  not _64525_ (_19088_, _18617_);
  and _64526_ (_19089_, _18776_, _19088_);
  and _64527_ (_19090_, _18773_, _18403_);
  not _64528_ (_19091_, _19090_);
  nor _64529_ (_19092_, _19091_, _19089_);
  and _64530_ (_19093_, _18780_, _18799_);
  nand _64531_ (_19094_, _18785_, _18817_);
  and _64532_ (_19095_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _64533_ (_19096_, _18785_, word_in[0]);
  and _64534_ (_19097_, _19096_, _18817_);
  or _64535_ (_19098_, _19097_, _19095_);
  or _64536_ (_19099_, _19098_, _19093_);
  not _64537_ (_19100_, _19093_);
  or _64538_ (_19101_, _19100_, word_in[8]);
  and _64539_ (_19102_, _19101_, _19099_);
  or _64540_ (_19103_, _19102_, _19092_);
  and _64541_ (_19104_, _18776_, word_in[16]);
  not _64542_ (_19105_, _19092_);
  or _64543_ (_19106_, _19105_, _19104_);
  and _64544_ (_19107_, _19106_, _19103_);
  or _64545_ (_19108_, _19107_, _19087_);
  not _64546_ (_19109_, _19087_);
  or _64547_ (_19110_, _19109_, word_in[24]);
  and _64548_ (_36786_, _19110_, _19108_);
  and _64549_ (_19111_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _64550_ (_19112_, _18785_, word_in[1]);
  and _64551_ (_19113_, _19112_, _18817_);
  nor _64552_ (_19114_, _19113_, _19111_);
  nor _64553_ (_19115_, _19114_, _19093_);
  and _64554_ (_19116_, _19093_, word_in[9]);
  nor _64555_ (_19117_, _19116_, _19115_);
  nor _64556_ (_19118_, _19117_, _19092_);
  and _64557_ (_19119_, _18776_, word_in[17]);
  and _64558_ (_19120_, _19092_, _19119_);
  or _64559_ (_19121_, _19120_, _19087_);
  or _64560_ (_19122_, _19121_, _19118_);
  or _64561_ (_19123_, _19109_, word_in[25]);
  and _64562_ (_36787_, _19123_, _19122_);
  and _64563_ (_19124_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _64564_ (_19125_, _18785_, word_in[2]);
  and _64565_ (_19126_, _19125_, _18817_);
  nor _64566_ (_19127_, _19126_, _19124_);
  nor _64567_ (_19128_, _19127_, _19093_);
  and _64568_ (_19129_, _19093_, word_in[10]);
  nor _64569_ (_19130_, _19129_, _19128_);
  nor _64570_ (_19131_, _19130_, _19092_);
  and _64571_ (_19132_, _18776_, word_in[18]);
  and _64572_ (_19133_, _19092_, _19132_);
  or _64573_ (_19134_, _19133_, _19087_);
  or _64574_ (_19135_, _19134_, _19131_);
  or _64575_ (_19136_, _19109_, word_in[26]);
  and _64576_ (_36788_, _19136_, _19135_);
  and _64577_ (_19137_, _18785_, word_in[3]);
  and _64578_ (_19138_, _19137_, _18817_);
  and _64579_ (_19139_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _64580_ (_19140_, _19139_, _19138_);
  nor _64581_ (_19141_, _19140_, _19093_);
  and _64582_ (_19142_, _19093_, word_in[11]);
  nor _64583_ (_19143_, _19142_, _19141_);
  nor _64584_ (_19144_, _19143_, _19092_);
  and _64585_ (_19145_, _18776_, word_in[19]);
  and _64586_ (_19146_, _19092_, _19145_);
  or _64587_ (_19147_, _19146_, _19087_);
  or _64588_ (_19148_, _19147_, _19144_);
  or _64589_ (_19149_, _19109_, word_in[27]);
  and _64590_ (_36789_, _19149_, _19148_);
  and _64591_ (_19150_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _64592_ (_19151_, _18785_, word_in[4]);
  and _64593_ (_19152_, _19151_, _18817_);
  or _64594_ (_19153_, _19152_, _19150_);
  or _64595_ (_19154_, _19153_, _19093_);
  or _64596_ (_19155_, _19100_, word_in[12]);
  and _64597_ (_19156_, _19155_, _19154_);
  or _64598_ (_19157_, _19156_, _19092_);
  and _64599_ (_19158_, _18776_, word_in[20]);
  or _64600_ (_19159_, _19105_, _19158_);
  and _64601_ (_19160_, _19159_, _19157_);
  or _64602_ (_19161_, _19160_, _19087_);
  or _64603_ (_19162_, _19109_, word_in[28]);
  and _64604_ (_36790_, _19162_, _19161_);
  and _64605_ (_19163_, _18785_, word_in[5]);
  and _64606_ (_19164_, _19163_, _18817_);
  and _64607_ (_19165_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _64608_ (_19166_, _19165_, _19164_);
  nor _64609_ (_19167_, _19166_, _19093_);
  and _64610_ (_19168_, _19093_, word_in[13]);
  nor _64611_ (_19169_, _19168_, _19167_);
  nor _64612_ (_19170_, _19169_, _19092_);
  and _64613_ (_19171_, _18776_, word_in[21]);
  and _64614_ (_19172_, _19092_, _19171_);
  or _64615_ (_19173_, _19172_, _19087_);
  or _64616_ (_19174_, _19173_, _19170_);
  or _64617_ (_19175_, _19109_, word_in[29]);
  and _64618_ (_36791_, _19175_, _19174_);
  and _64619_ (_19176_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _64620_ (_19177_, _18785_, word_in[6]);
  and _64621_ (_19178_, _19177_, _18817_);
  nor _64622_ (_19179_, _19178_, _19176_);
  nor _64623_ (_19180_, _19179_, _19093_);
  and _64624_ (_19181_, _19093_, word_in[14]);
  nor _64625_ (_19182_, _19181_, _19180_);
  nor _64626_ (_19183_, _19182_, _19092_);
  and _64627_ (_19184_, _18776_, word_in[22]);
  and _64628_ (_19185_, _19092_, _19184_);
  or _64629_ (_19186_, _19185_, _19087_);
  or _64630_ (_19187_, _19186_, _19183_);
  or _64631_ (_19188_, _19109_, word_in[30]);
  and _64632_ (_36792_, _19188_, _19187_);
  and _64633_ (_19189_, _18785_, word_in[7]);
  and _64634_ (_19190_, _19189_, _18817_);
  and _64635_ (_19191_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _64636_ (_19192_, _19191_, _19190_);
  nor _64637_ (_19193_, _19192_, _19093_);
  and _64638_ (_19194_, _19093_, word_in[15]);
  nor _64639_ (_19195_, _19194_, _19193_);
  nor _64640_ (_19196_, _19195_, _19092_);
  and _64641_ (_19197_, _19092_, _18795_);
  or _64642_ (_19198_, _19197_, _19087_);
  or _64643_ (_19199_, _19198_, _19196_);
  or _64644_ (_19200_, _19109_, word_in[31]);
  and _64645_ (_36793_, _19200_, _19199_);
  and _64646_ (_19201_, _18767_, _18404_);
  and _64647_ (_19202_, _19201_, _18977_);
  not _64648_ (_19203_, _19202_);
  not _64649_ (_19204_, _18773_);
  and _64650_ (_19205_, _18980_, _19204_);
  and _64651_ (_19206_, _19205_, _18617_);
  and _64652_ (_19207_, _18780_, _18817_);
  and _64653_ (_19208_, _19096_, _18807_);
  nand _64654_ (_19209_, _18785_, _18807_);
  and _64655_ (_19210_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor _64656_ (_19211_, _19210_, _19208_);
  nor _64657_ (_19212_, _19211_, _19207_);
  and _64658_ (_19213_, _19207_, word_in[8]);
  nor _64659_ (_19214_, _19213_, _19212_);
  nor _64660_ (_19215_, _19214_, _19206_);
  and _64661_ (_19216_, _19206_, _19104_);
  or _64662_ (_19217_, _19216_, _19215_);
  and _64663_ (_19218_, _19217_, _19203_);
  and _64664_ (_19219_, _19202_, word_in[24]);
  or _64665_ (_36794_, _19219_, _19218_);
  and _64666_ (_19220_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _64667_ (_19221_, _19112_, _18807_);
  nor _64668_ (_19222_, _19221_, _19220_);
  nor _64669_ (_19223_, _19222_, _19207_);
  and _64670_ (_19224_, _19207_, word_in[9]);
  nor _64671_ (_19225_, _19224_, _19223_);
  nor _64672_ (_19226_, _19225_, _19206_);
  and _64673_ (_19227_, _19206_, _19119_);
  or _64674_ (_19228_, _19227_, _19226_);
  and _64675_ (_19229_, _19228_, _19203_);
  and _64676_ (_19230_, _19202_, word_in[25]);
  or _64677_ (_36795_, _19230_, _19229_);
  and _64678_ (_19231_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _64679_ (_19232_, _19125_, _18807_);
  nor _64680_ (_19233_, _19232_, _19231_);
  nor _64681_ (_19234_, _19233_, _19207_);
  and _64682_ (_19235_, _19207_, word_in[10]);
  nor _64683_ (_19236_, _19235_, _19234_);
  nor _64684_ (_19237_, _19236_, _19206_);
  and _64685_ (_19238_, _19206_, _19132_);
  or _64686_ (_19239_, _19238_, _19237_);
  and _64687_ (_19240_, _19239_, _19203_);
  and _64688_ (_19241_, _19202_, word_in[26]);
  or _64689_ (_36796_, _19241_, _19240_);
  and _64690_ (_19242_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _64691_ (_19243_, _19137_, _18807_);
  nor _64692_ (_19244_, _19243_, _19242_);
  nor _64693_ (_19245_, _19244_, _19207_);
  and _64694_ (_19246_, _19207_, word_in[11]);
  nor _64695_ (_19247_, _19246_, _19245_);
  nor _64696_ (_19248_, _19247_, _19206_);
  and _64697_ (_19249_, _19206_, _19145_);
  or _64698_ (_19250_, _19249_, _19248_);
  and _64699_ (_19251_, _19250_, _19203_);
  and _64700_ (_19252_, _19202_, word_in[27]);
  or _64701_ (_36797_, _19252_, _19251_);
  and _64702_ (_19253_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _64703_ (_19254_, _19151_, _18807_);
  or _64704_ (_19255_, _19254_, _19253_);
  or _64705_ (_19256_, _19255_, _19207_);
  not _64706_ (_19257_, word_in[12]);
  nand _64707_ (_19258_, _19207_, _19257_);
  nand _64708_ (_19259_, _19258_, _19256_);
  nor _64709_ (_19260_, _19259_, _19206_);
  and _64710_ (_19261_, _19206_, _19158_);
  or _64711_ (_19262_, _19261_, _19260_);
  or _64712_ (_19263_, _19262_, _19202_);
  or _64713_ (_19264_, _19203_, word_in[28]);
  and _64714_ (_36798_, _19264_, _19263_);
  and _64715_ (_19265_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _64716_ (_19266_, _19163_, _18807_);
  nor _64717_ (_19267_, _19266_, _19265_);
  nor _64718_ (_19268_, _19267_, _19207_);
  and _64719_ (_19269_, _19207_, word_in[13]);
  nor _64720_ (_19270_, _19269_, _19268_);
  nor _64721_ (_19271_, _19270_, _19206_);
  and _64722_ (_19272_, _19206_, _19171_);
  or _64723_ (_19273_, _19272_, _19271_);
  and _64724_ (_19274_, _19273_, _19203_);
  and _64725_ (_19275_, _19202_, word_in[29]);
  or _64726_ (_36799_, _19275_, _19274_);
  and _64727_ (_19276_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _64728_ (_19277_, _19177_, _18807_);
  nor _64729_ (_19278_, _19277_, _19276_);
  nor _64730_ (_19279_, _19278_, _19207_);
  and _64731_ (_19280_, _19207_, word_in[14]);
  nor _64732_ (_19281_, _19280_, _19279_);
  nor _64733_ (_19282_, _19281_, _19206_);
  and _64734_ (_19283_, _19206_, _19184_);
  or _64735_ (_19284_, _19283_, _19282_);
  and _64736_ (_19285_, _19284_, _19203_);
  and _64737_ (_19286_, _19202_, word_in[30]);
  or _64738_ (_36800_, _19286_, _19285_);
  and _64739_ (_19287_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _64740_ (_19288_, _19189_, _18807_);
  nor _64741_ (_19289_, _19288_, _19287_);
  nor _64742_ (_19290_, _19289_, _19207_);
  and _64743_ (_19291_, _19207_, word_in[15]);
  nor _64744_ (_19292_, _19291_, _19290_);
  nor _64745_ (_19293_, _19292_, _19206_);
  and _64746_ (_19294_, _19206_, _18795_);
  or _64747_ (_19295_, _19294_, _19293_);
  and _64748_ (_19296_, _19295_, _19203_);
  and _64749_ (_19297_, _19202_, word_in[31]);
  or _64750_ (_36801_, _19297_, _19296_);
  and _64751_ (_19298_, _18767_, _18799_);
  not _64752_ (_19299_, _19298_);
  not _64753_ (_19300_, _18774_);
  nor _64754_ (_19301_, _19089_, _19300_);
  and _64755_ (_19302_, _18780_, _18807_);
  nand _64756_ (_19303_, _18785_, _18816_);
  and _64757_ (_19304_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _64758_ (_19305_, _19096_, _18816_);
  nor _64759_ (_19306_, _19305_, _19304_);
  nor _64760_ (_19307_, _19306_, _19302_);
  and _64761_ (_19308_, _19302_, word_in[8]);
  nor _64762_ (_19309_, _19308_, _19307_);
  nor _64763_ (_19310_, _19309_, _19301_);
  and _64764_ (_19311_, _19301_, _19104_);
  or _64765_ (_19312_, _19311_, _19310_);
  and _64766_ (_19313_, _19312_, _19299_);
  and _64767_ (_19314_, _19298_, word_in[24]);
  or _64768_ (_36802_, _19314_, _19313_);
  and _64769_ (_19315_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _64770_ (_19316_, _19112_, _18816_);
  nor _64771_ (_19317_, _19316_, _19315_);
  nor _64772_ (_19318_, _19317_, _19302_);
  and _64773_ (_19319_, _19302_, word_in[9]);
  nor _64774_ (_19320_, _19319_, _19318_);
  nor _64775_ (_19321_, _19320_, _19301_);
  and _64776_ (_19322_, _19301_, _19119_);
  or _64777_ (_19323_, _19322_, _19321_);
  and _64778_ (_19324_, _19323_, _19299_);
  and _64779_ (_19325_, _19298_, word_in[25]);
  or _64780_ (_36803_, _19325_, _19324_);
  and _64781_ (_19326_, _19125_, _18816_);
  and _64782_ (_19327_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor _64783_ (_19328_, _19327_, _19326_);
  nor _64784_ (_19329_, _19328_, _19302_);
  and _64785_ (_19330_, _19302_, word_in[10]);
  nor _64786_ (_19331_, _19330_, _19329_);
  nor _64787_ (_19332_, _19331_, _19301_);
  and _64788_ (_19333_, _19301_, _19132_);
  or _64789_ (_19334_, _19333_, _19332_);
  and _64790_ (_19335_, _19334_, _19299_);
  and _64791_ (_19336_, _19298_, word_in[26]);
  or _64792_ (_36804_, _19336_, _19335_);
  and _64793_ (_19337_, _19137_, _18816_);
  and _64794_ (_19338_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _64795_ (_19339_, _19338_, _19337_);
  nor _64796_ (_19340_, _19339_, _19302_);
  and _64797_ (_19341_, _19302_, word_in[11]);
  nor _64798_ (_19342_, _19341_, _19340_);
  nor _64799_ (_19343_, _19342_, _19301_);
  and _64800_ (_19344_, _19301_, _19145_);
  or _64801_ (_19345_, _19344_, _19343_);
  and _64802_ (_19346_, _19345_, _19299_);
  and _64803_ (_19347_, _19298_, word_in[27]);
  or _64804_ (_36805_, _19347_, _19346_);
  and _64805_ (_19348_, _19298_, _19038_);
  and _64806_ (_19349_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _64807_ (_19350_, _19151_, _18816_);
  or _64808_ (_19351_, _19350_, _19349_);
  or _64809_ (_19352_, _19351_, _19302_);
  nand _64810_ (_19353_, _19302_, _19257_);
  and _64811_ (_19354_, _19353_, _19352_);
  or _64812_ (_19355_, _19354_, _19301_);
  not _64813_ (_19356_, _19301_);
  or _64814_ (_19357_, _19356_, _19158_);
  and _64815_ (_19358_, _19357_, _19299_);
  and _64816_ (_19359_, _19358_, _19355_);
  or _64817_ (_36806_, _19359_, _19348_);
  and _64818_ (_19360_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _64819_ (_19361_, _19163_, _18816_);
  nor _64820_ (_19362_, _19361_, _19360_);
  nor _64821_ (_19363_, _19362_, _19302_);
  and _64822_ (_19364_, _19302_, word_in[13]);
  nor _64823_ (_19365_, _19364_, _19363_);
  nor _64824_ (_19366_, _19365_, _19301_);
  and _64825_ (_19367_, _19301_, _19171_);
  or _64826_ (_19368_, _19367_, _19366_);
  and _64827_ (_19369_, _19368_, _19299_);
  and _64828_ (_19370_, _19298_, word_in[29]);
  or _64829_ (_36807_, _19370_, _19369_);
  and _64830_ (_19371_, _19177_, _18816_);
  and _64831_ (_19372_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _64832_ (_19373_, _19372_, _19371_);
  nor _64833_ (_19374_, _19373_, _19302_);
  and _64834_ (_19375_, _19302_, word_in[14]);
  nor _64835_ (_19376_, _19375_, _19374_);
  nor _64836_ (_19377_, _19376_, _19301_);
  and _64837_ (_19378_, _19301_, _19184_);
  or _64838_ (_19379_, _19378_, _19377_);
  and _64839_ (_19380_, _19379_, _19299_);
  and _64840_ (_19381_, _19298_, word_in[30]);
  or _64841_ (_36808_, _19381_, _19380_);
  and _64842_ (_19382_, _19189_, _18816_);
  and _64843_ (_19383_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  or _64844_ (_19384_, _19383_, _19382_);
  or _64845_ (_19385_, _19384_, _19302_);
  not _64846_ (_19386_, word_in[15]);
  nand _64847_ (_19387_, _19302_, _19386_);
  and _64848_ (_19388_, _19387_, _19385_);
  or _64849_ (_19389_, _19388_, _19301_);
  or _64850_ (_19390_, _19356_, _18795_);
  and _64851_ (_19391_, _19390_, _19389_);
  or _64852_ (_19392_, _19391_, _19298_);
  or _64853_ (_19393_, _19299_, word_in[31]);
  and _64854_ (_36809_, _19393_, _19392_);
  and _64855_ (_19394_, _18975_, _18752_);
  and _64856_ (_19395_, _19394_, _18426_);
  not _64857_ (_19396_, _19395_);
  not _64858_ (_19397_, _18916_);
  and _64859_ (_19398_, _19397_, _18776_);
  and _64860_ (_19399_, _19398_, _18981_);
  and _64861_ (_19400_, _18781_, _18504_);
  and _64862_ (_19401_, _19400_, _18404_);
  nand _64863_ (_19402_, _18785_, _18811_);
  and _64864_ (_19403_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _64865_ (_19404_, _19096_, _18811_);
  nor _64866_ (_19405_, _19404_, _19403_);
  nor _64867_ (_19406_, _19405_, _19401_);
  and _64868_ (_19407_, _18780_, word_in[8]);
  and _64869_ (_19408_, _19401_, _19407_);
  nor _64870_ (_19409_, _19408_, _19406_);
  nor _64871_ (_19410_, _19409_, _19399_);
  and _64872_ (_19411_, _19399_, _19104_);
  or _64873_ (_19412_, _19411_, _19410_);
  and _64874_ (_19413_, _19412_, _19396_);
  and _64875_ (_19414_, _18767_, word_in[24]);
  and _64876_ (_19415_, _19395_, _19414_);
  or _64877_ (_36810_, _19415_, _19413_);
  and _64878_ (_19416_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _64879_ (_19417_, _19112_, _18811_);
  nor _64880_ (_19418_, _19417_, _19416_);
  nor _64881_ (_19419_, _19418_, _19401_);
  and _64882_ (_19420_, _19401_, _19001_);
  nor _64883_ (_19421_, _19420_, _19419_);
  nor _64884_ (_19422_, _19421_, _19399_);
  and _64885_ (_19423_, _19399_, _19119_);
  or _64886_ (_19424_, _19423_, _19422_);
  and _64887_ (_19425_, _19424_, _19396_);
  and _64888_ (_19426_, _18767_, word_in[25]);
  and _64889_ (_19427_, _19395_, _19426_);
  or _64890_ (_36811_, _19427_, _19425_);
  and _64891_ (_19428_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _64892_ (_19429_, _19125_, _18811_);
  nor _64893_ (_19430_, _19429_, _19428_);
  nor _64894_ (_19431_, _19430_, _19401_);
  and _64895_ (_19432_, _18780_, word_in[10]);
  and _64896_ (_19433_, _19401_, _19432_);
  nor _64897_ (_19434_, _19433_, _19431_);
  nor _64898_ (_19435_, _19434_, _19399_);
  and _64899_ (_19436_, _19399_, _19132_);
  or _64900_ (_19437_, _19436_, _19395_);
  or _64901_ (_19438_, _19437_, _19435_);
  and _64902_ (_19439_, _18767_, word_in[26]);
  or _64903_ (_19440_, _19396_, _19439_);
  and _64904_ (_36812_, _19440_, _19438_);
  and _64905_ (_19441_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _64906_ (_19442_, _19137_, _18811_);
  nor _64907_ (_19443_, _19442_, _19441_);
  nor _64908_ (_19444_, _19443_, _19401_);
  and _64909_ (_19445_, _18780_, word_in[11]);
  and _64910_ (_19446_, _19401_, _19445_);
  nor _64911_ (_19447_, _19446_, _19444_);
  nor _64912_ (_19448_, _19447_, _19399_);
  and _64913_ (_19449_, _19399_, _19145_);
  or _64914_ (_19450_, _19449_, _19448_);
  and _64915_ (_19451_, _19450_, _19396_);
  and _64916_ (_19452_, _18767_, word_in[27]);
  and _64917_ (_19453_, _19395_, _19452_);
  or _64918_ (_36813_, _19453_, _19451_);
  and _64919_ (_19454_, _18780_, word_in[12]);
  not _64920_ (_19455_, _19401_);
  or _64921_ (_19456_, _19455_, _19454_);
  and _64922_ (_19457_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _64923_ (_19458_, _19151_, _18811_);
  or _64924_ (_19459_, _19458_, _19457_);
  or _64925_ (_19460_, _19459_, _19401_);
  and _64926_ (_19461_, _19460_, _19456_);
  or _64927_ (_19462_, _19461_, _19399_);
  not _64928_ (_19463_, _19399_);
  or _64929_ (_19464_, _19463_, _19158_);
  and _64930_ (_19465_, _19464_, _19396_);
  and _64931_ (_19466_, _19465_, _19462_);
  and _64932_ (_19467_, _19395_, _19038_);
  or _64933_ (_36814_, _19467_, _19466_);
  and _64934_ (_19468_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _64935_ (_19469_, _19163_, _18811_);
  nor _64936_ (_19470_, _19469_, _19468_);
  nor _64937_ (_19471_, _19470_, _19401_);
  and _64938_ (_19472_, _18780_, word_in[13]);
  and _64939_ (_19473_, _19401_, _19472_);
  nor _64940_ (_19474_, _19473_, _19471_);
  nor _64941_ (_19475_, _19474_, _19399_);
  and _64942_ (_19476_, _19399_, _19171_);
  or _64943_ (_19477_, _19476_, _19475_);
  and _64944_ (_19478_, _19477_, _19396_);
  and _64945_ (_19479_, _18767_, word_in[29]);
  and _64946_ (_19480_, _19395_, _19479_);
  or _64947_ (_36815_, _19480_, _19478_);
  and _64948_ (_19481_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _64949_ (_19482_, _19177_, _18811_);
  nor _64950_ (_19483_, _19482_, _19481_);
  nor _64951_ (_19484_, _19483_, _19401_);
  and _64952_ (_19485_, _18780_, word_in[14]);
  and _64953_ (_19486_, _19401_, _19485_);
  nor _64954_ (_19487_, _19486_, _19484_);
  nor _64955_ (_19488_, _19487_, _19399_);
  and _64956_ (_19489_, _19399_, _19184_);
  or _64957_ (_19490_, _19489_, _19488_);
  and _64958_ (_19491_, _19490_, _19396_);
  and _64959_ (_19492_, _18767_, word_in[30]);
  and _64960_ (_19493_, _19395_, _19492_);
  or _64961_ (_36816_, _19493_, _19491_);
  or _64962_ (_19494_, _19455_, _18791_);
  and _64963_ (_19495_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _64964_ (_19496_, _19189_, _18811_);
  or _64965_ (_19497_, _19496_, _19495_);
  or _64966_ (_19498_, _19497_, _19401_);
  and _64967_ (_19499_, _19498_, _19494_);
  or _64968_ (_19500_, _19499_, _19399_);
  or _64969_ (_19501_, _19463_, _18795_);
  and _64970_ (_19502_, _19501_, _19396_);
  and _64971_ (_19503_, _19502_, _19500_);
  and _64972_ (_19504_, _19395_, _18768_);
  or _64973_ (_36857_[7], _19504_, _19503_);
  and _64974_ (_19505_, _19398_, _19090_);
  and _64975_ (_19506_, _19400_, _18414_);
  and _64976_ (_19507_, _19096_, _18824_);
  nand _64977_ (_19508_, _18785_, _18824_);
  and _64978_ (_19509_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  or _64979_ (_19510_, _19509_, _19507_);
  or _64980_ (_19511_, _19510_, _19506_);
  not _64981_ (_19512_, _19506_);
  or _64982_ (_19513_, _19512_, _19407_);
  and _64983_ (_19514_, _19513_, _19511_);
  or _64984_ (_19515_, _19514_, _19505_);
  and _64985_ (_19516_, _19394_, _18437_);
  not _64986_ (_19517_, _19516_);
  not _64987_ (_19518_, _19505_);
  or _64988_ (_19519_, _19518_, _19104_);
  and _64989_ (_19520_, _19519_, _19517_);
  and _64990_ (_19521_, _19520_, _19515_);
  and _64991_ (_19522_, _19516_, _19414_);
  or _64992_ (_36817_, _19522_, _19521_);
  and _64993_ (_19523_, _19112_, _18824_);
  and _64994_ (_19524_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  or _64995_ (_19525_, _19524_, _19523_);
  or _64996_ (_19526_, _19525_, _19506_);
  or _64997_ (_19527_, _19512_, _19001_);
  and _64998_ (_19528_, _19527_, _19526_);
  or _64999_ (_19529_, _19528_, _19505_);
  or _65000_ (_19530_, _19518_, _19119_);
  and _65001_ (_19531_, _19530_, _19517_);
  and _65002_ (_19532_, _19531_, _19529_);
  and _65003_ (_19533_, _19516_, _19426_);
  or _65004_ (_36818_, _19533_, _19532_);
  and _65005_ (_19534_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and _65006_ (_19535_, _19125_, _18824_);
  nor _65007_ (_19536_, _19535_, _19534_);
  nor _65008_ (_19537_, _19536_, _19506_);
  and _65009_ (_19538_, _19506_, _19432_);
  or _65010_ (_19539_, _19538_, _19537_);
  and _65011_ (_19540_, _19539_, _19518_);
  and _65012_ (_19541_, _19505_, _19132_);
  or _65013_ (_19542_, _19541_, _19516_);
  or _65014_ (_19543_, _19542_, _19540_);
  or _65015_ (_19544_, _19517_, _19439_);
  and _65016_ (_36819_, _19544_, _19543_);
  and _65017_ (_19545_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and _65018_ (_19546_, _19137_, _18824_);
  nor _65019_ (_19547_, _19546_, _19545_);
  nor _65020_ (_19548_, _19547_, _19506_);
  and _65021_ (_19549_, _19506_, _19445_);
  or _65022_ (_19550_, _19549_, _19548_);
  and _65023_ (_19551_, _19550_, _19518_);
  and _65024_ (_19552_, _19505_, _19145_);
  or _65025_ (_19553_, _19552_, _19516_);
  or _65026_ (_19554_, _19553_, _19551_);
  or _65027_ (_19555_, _19517_, _19452_);
  and _65028_ (_36820_, _19555_, _19554_);
  and _65029_ (_19556_, _19505_, _19158_);
  and _65030_ (_19557_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _65031_ (_19558_, _19151_, _18824_);
  nor _65032_ (_19559_, _19558_, _19557_);
  nor _65033_ (_19560_, _19559_, _19506_);
  and _65034_ (_19561_, _19506_, _19454_);
  or _65035_ (_19562_, _19561_, _19560_);
  and _65036_ (_19563_, _19562_, _19518_);
  or _65037_ (_19564_, _19563_, _19556_);
  and _65038_ (_19565_, _19564_, _19517_);
  and _65039_ (_19566_, _19516_, _19038_);
  or _65040_ (_36821_, _19566_, _19565_);
  and _65041_ (_19567_, _19505_, _19171_);
  and _65042_ (_19568_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and _65043_ (_19569_, _19163_, _18824_);
  nor _65044_ (_19570_, _19569_, _19568_);
  nor _65045_ (_19571_, _19570_, _19506_);
  and _65046_ (_19572_, _19506_, _19472_);
  or _65047_ (_19573_, _19572_, _19571_);
  and _65048_ (_19574_, _19573_, _19518_);
  or _65049_ (_19575_, _19574_, _19567_);
  and _65050_ (_19576_, _19575_, _19517_);
  and _65051_ (_19577_, _19516_, _19479_);
  or _65052_ (_36822_, _19577_, _19576_);
  and _65053_ (_19578_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _65054_ (_19579_, _19177_, _18824_);
  nor _65055_ (_19580_, _19579_, _19578_);
  nor _65056_ (_19581_, _19580_, _19506_);
  and _65057_ (_19582_, _19506_, _19485_);
  or _65058_ (_19583_, _19582_, _19581_);
  and _65059_ (_19584_, _19583_, _19518_);
  and _65060_ (_19585_, _19505_, _19184_);
  or _65061_ (_19586_, _19585_, _19516_);
  or _65062_ (_19587_, _19586_, _19584_);
  or _65063_ (_19588_, _19517_, _19492_);
  and _65064_ (_36823_, _19588_, _19587_);
  and _65065_ (_19589_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _65066_ (_19590_, _19189_, _18824_);
  nor _65067_ (_19591_, _19590_, _19589_);
  nor _65068_ (_19592_, _19591_, _19506_);
  and _65069_ (_19593_, _19506_, _18791_);
  or _65070_ (_19594_, _19593_, _19592_);
  and _65071_ (_19595_, _19594_, _19518_);
  and _65072_ (_19596_, _19505_, _18795_);
  or _65073_ (_19597_, _19596_, _19516_);
  or _65074_ (_19598_, _19597_, _19595_);
  or _65075_ (_19599_, _19517_, _18768_);
  and _65076_ (_36824_, _19599_, _19598_);
  and _65077_ (_19600_, _19205_, _19397_);
  and _65078_ (_19601_, _19400_, _18426_);
  and _65079_ (_19602_, _18785_, _18847_);
  and _65080_ (_19603_, _19602_, word_in[0]);
  not _65081_ (_19604_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor _65082_ (_19605_, _19602_, _19604_);
  nor _65083_ (_19606_, _19605_, _19603_);
  nor _65084_ (_19607_, _19606_, _19601_);
  and _65085_ (_19608_, _19601_, _19407_);
  or _65086_ (_19609_, _19608_, _19607_);
  or _65087_ (_19610_, _19609_, _19600_);
  and _65088_ (_19611_, _19394_, _18404_);
  not _65089_ (_19612_, _19611_);
  not _65090_ (_19613_, _19600_);
  or _65091_ (_19614_, _19613_, _19104_);
  and _65092_ (_19615_, _19614_, _19612_);
  and _65093_ (_19616_, _19615_, _19610_);
  and _65094_ (_19617_, _19611_, _19414_);
  or _65095_ (_36825_, _19617_, _19616_);
  not _65096_ (_19618_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _65097_ (_19619_, _19602_, _19618_);
  and _65098_ (_19620_, _19602_, _19112_);
  or _65099_ (_19621_, _19620_, _19619_);
  or _65100_ (_19622_, _19621_, _19601_);
  not _65101_ (_19623_, _19601_);
  or _65102_ (_19624_, _19623_, _19001_);
  and _65103_ (_19625_, _19624_, _19622_);
  or _65104_ (_19626_, _19625_, _19600_);
  or _65105_ (_19627_, _19613_, _19119_);
  and _65106_ (_19628_, _19627_, _19612_);
  and _65107_ (_19629_, _19628_, _19626_);
  and _65108_ (_19630_, _19611_, _19426_);
  or _65109_ (_36826_, _19630_, _19629_);
  and _65110_ (_19631_, _19602_, word_in[2]);
  not _65111_ (_19632_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor _65112_ (_19633_, _19602_, _19632_);
  nor _65113_ (_19634_, _19633_, _19631_);
  nor _65114_ (_19635_, _19634_, _19601_);
  and _65115_ (_19636_, _19601_, _19432_);
  nor _65116_ (_19637_, _19636_, _19635_);
  nor _65117_ (_19638_, _19637_, _19600_);
  and _65118_ (_19639_, _19600_, _19132_);
  or _65119_ (_19640_, _19639_, _19611_);
  or _65120_ (_19641_, _19640_, _19638_);
  or _65121_ (_19642_, _19612_, _19439_);
  and _65122_ (_36827_, _19642_, _19641_);
  and _65123_ (_19643_, _19600_, _19145_);
  and _65124_ (_19644_, _19602_, word_in[3]);
  not _65125_ (_19645_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _65126_ (_19646_, _19602_, _19645_);
  nor _65127_ (_19647_, _19646_, _19644_);
  nor _65128_ (_19648_, _19647_, _19601_);
  and _65129_ (_19649_, _19601_, _19445_);
  nor _65130_ (_19650_, _19649_, _19648_);
  nor _65131_ (_19651_, _19650_, _19600_);
  or _65132_ (_19652_, _19651_, _19643_);
  and _65133_ (_19653_, _19652_, _19612_);
  and _65134_ (_19654_, _19611_, _19452_);
  or _65135_ (_36828_, _19654_, _19653_);
  and _65136_ (_19655_, _19600_, _19158_);
  and _65137_ (_19656_, _19602_, word_in[4]);
  not _65138_ (_19657_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor _65139_ (_19658_, _19602_, _19657_);
  nor _65140_ (_19659_, _19658_, _19656_);
  nor _65141_ (_19660_, _19659_, _19601_);
  and _65142_ (_19661_, _19601_, _19454_);
  nor _65143_ (_19662_, _19661_, _19660_);
  nor _65144_ (_19663_, _19662_, _19600_);
  or _65145_ (_19664_, _19663_, _19655_);
  and _65146_ (_19665_, _19664_, _19612_);
  and _65147_ (_19666_, _19611_, _19038_);
  or _65148_ (_36829_, _19666_, _19665_);
  not _65149_ (_19667_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _65150_ (_19668_, _19602_, _19667_);
  and _65151_ (_19669_, _19602_, _19163_);
  or _65152_ (_19670_, _19669_, _19668_);
  or _65153_ (_19671_, _19670_, _19601_);
  or _65154_ (_19672_, _19623_, _19472_);
  and _65155_ (_19673_, _19672_, _19671_);
  or _65156_ (_19674_, _19673_, _19600_);
  or _65157_ (_19675_, _19613_, _19171_);
  and _65158_ (_19676_, _19675_, _19612_);
  and _65159_ (_19677_, _19676_, _19674_);
  and _65160_ (_19678_, _19611_, _19479_);
  or _65161_ (_36830_, _19678_, _19677_);
  not _65162_ (_19679_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _65163_ (_19680_, _19602_, _19679_);
  and _65164_ (_19681_, _19602_, _19177_);
  or _65165_ (_19682_, _19681_, _19680_);
  or _65166_ (_19683_, _19682_, _19601_);
  or _65167_ (_19684_, _19623_, _19485_);
  and _65168_ (_19685_, _19684_, _19683_);
  or _65169_ (_19686_, _19685_, _19600_);
  or _65170_ (_19687_, _19613_, _19184_);
  and _65171_ (_19688_, _19687_, _19612_);
  and _65172_ (_19689_, _19688_, _19686_);
  and _65173_ (_19690_, _19611_, _19492_);
  or _65174_ (_36831_, _19690_, _19689_);
  and _65175_ (_19691_, _19602_, word_in[7]);
  nor _65176_ (_19692_, _19602_, _18572_);
  nor _65177_ (_19693_, _19692_, _19691_);
  nor _65178_ (_19694_, _19693_, _19601_);
  and _65179_ (_19695_, _19601_, _18791_);
  nor _65180_ (_19696_, _19695_, _19694_);
  nor _65181_ (_19697_, _19696_, _19600_);
  and _65182_ (_19698_, _19600_, _18795_);
  or _65183_ (_19699_, _19698_, _19697_);
  and _65184_ (_19700_, _19699_, _19612_);
  and _65185_ (_19701_, _19611_, _18768_);
  or _65186_ (_36832_, _19701_, _19700_);
  and _65187_ (_19702_, _18767_, _18811_);
  and _65188_ (_19703_, _19398_, _18774_);
  and _65189_ (_19704_, _19400_, _18437_);
  not _65190_ (_19705_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _65191_ (_19706_, _18785_, _18503_);
  nor _65192_ (_19707_, _19706_, _19705_);
  and _65193_ (_19708_, _19706_, _19096_);
  or _65194_ (_19709_, _19708_, _19707_);
  or _65195_ (_19710_, _19709_, _19704_);
  not _65196_ (_19711_, _19704_);
  or _65197_ (_19712_, _19711_, _19407_);
  and _65198_ (_19713_, _19712_, _19710_);
  or _65199_ (_19714_, _19713_, _19703_);
  not _65200_ (_19715_, _19703_);
  or _65201_ (_19716_, _19715_, word_in[16]);
  and _65202_ (_19717_, _19716_, _19714_);
  or _65203_ (_19718_, _19717_, _19702_);
  not _65204_ (_19719_, _19702_);
  or _65205_ (_19720_, _19719_, word_in[24]);
  and _65206_ (_36833_, _19720_, _19718_);
  not _65207_ (_19721_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor _65208_ (_19722_, _19706_, _19721_);
  and _65209_ (_19723_, _19706_, word_in[1]);
  nor _65210_ (_19724_, _19723_, _19722_);
  nor _65211_ (_19725_, _19724_, _19704_);
  and _65212_ (_19726_, _19704_, _19001_);
  or _65213_ (_19727_, _19726_, _19725_);
  and _65214_ (_19728_, _19727_, _19715_);
  and _65215_ (_19729_, _19703_, word_in[17]);
  or _65216_ (_19730_, _19729_, _19728_);
  and _65217_ (_19731_, _19730_, _19719_);
  and _65218_ (_19732_, _19702_, word_in[25]);
  or _65219_ (_36834_, _19732_, _19731_);
  and _65220_ (_19733_, _19702_, word_in[26]);
  and _65221_ (_19734_, _19706_, word_in[2]);
  not _65222_ (_19735_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _65223_ (_19736_, _19706_, _19735_);
  nor _65224_ (_19737_, _19736_, _19734_);
  nor _65225_ (_19738_, _19737_, _19704_);
  and _65226_ (_19739_, _19704_, _19432_);
  or _65227_ (_19740_, _19739_, _19738_);
  and _65228_ (_19741_, _19740_, _19715_);
  and _65229_ (_19742_, _19703_, word_in[18]);
  or _65230_ (_19743_, _19742_, _19741_);
  and _65231_ (_19744_, _19743_, _19719_);
  or _65232_ (_36835_, _19744_, _19733_);
  not _65233_ (_19745_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _65234_ (_19746_, _19706_, _19745_);
  and _65235_ (_19747_, _19706_, _19137_);
  or _65236_ (_19748_, _19747_, _19746_);
  or _65237_ (_19749_, _19748_, _19704_);
  or _65238_ (_19750_, _19711_, _19445_);
  and _65239_ (_19751_, _19750_, _19749_);
  or _65240_ (_19752_, _19751_, _19703_);
  or _65241_ (_19753_, _19715_, _19145_);
  and _65242_ (_19754_, _19753_, _19719_);
  and _65243_ (_19755_, _19754_, _19752_);
  and _65244_ (_19756_, _19702_, word_in[27]);
  or _65245_ (_36836_, _19756_, _19755_);
  and _65246_ (_19757_, _19038_, _18811_);
  and _65247_ (_19758_, _19706_, word_in[4]);
  not _65248_ (_19759_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor _65249_ (_19760_, _19706_, _19759_);
  nor _65250_ (_19761_, _19760_, _19758_);
  nor _65251_ (_19762_, _19761_, _19704_);
  and _65252_ (_19763_, _19704_, _19454_);
  or _65253_ (_19764_, _19763_, _19762_);
  or _65254_ (_19765_, _19764_, _19703_);
  or _65255_ (_19766_, _19715_, _19158_);
  and _65256_ (_19767_, _19766_, _19719_);
  and _65257_ (_19768_, _19767_, _19765_);
  or _65258_ (_36837_, _19768_, _19757_);
  and _65259_ (_19769_, _19706_, word_in[5]);
  not _65260_ (_19770_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor _65261_ (_19771_, _19706_, _19770_);
  nor _65262_ (_19772_, _19771_, _19769_);
  nor _65263_ (_19773_, _19772_, _19704_);
  and _65264_ (_19774_, _19704_, _19472_);
  or _65265_ (_19775_, _19774_, _19773_);
  and _65266_ (_19776_, _19775_, _19715_);
  and _65267_ (_19777_, _19703_, word_in[21]);
  or _65268_ (_19778_, _19777_, _19776_);
  and _65269_ (_19779_, _19778_, _19719_);
  and _65270_ (_19780_, _19702_, word_in[29]);
  or _65271_ (_36838_, _19780_, _19779_);
  and _65272_ (_19781_, _19702_, word_in[30]);
  not _65273_ (_19782_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor _65274_ (_19783_, _19706_, _19782_);
  and _65275_ (_19784_, _19706_, _19177_);
  or _65276_ (_19785_, _19784_, _19783_);
  or _65277_ (_19786_, _19785_, _19704_);
  or _65278_ (_19787_, _19711_, _19485_);
  and _65279_ (_19788_, _19787_, _19786_);
  or _65280_ (_19789_, _19788_, _19703_);
  or _65281_ (_19790_, _19715_, word_in[22]);
  and _65282_ (_19791_, _19790_, _19719_);
  and _65283_ (_19792_, _19791_, _19789_);
  or _65284_ (_36839_, _19792_, _19781_);
  and _65285_ (_19793_, _19702_, word_in[31]);
  and _65286_ (_19794_, _19706_, word_in[7]);
  nor _65287_ (_19795_, _19706_, _18451_);
  nor _65288_ (_19796_, _19795_, _19794_);
  nor _65289_ (_19797_, _19796_, _19704_);
  and _65290_ (_19798_, _19704_, _18791_);
  or _65291_ (_19799_, _19798_, _19797_);
  and _65292_ (_19800_, _19799_, _19715_);
  and _65293_ (_19801_, _19703_, word_in[23]);
  or _65294_ (_19802_, _19801_, _19800_);
  and _65295_ (_19803_, _19802_, _19719_);
  or _65296_ (_36840_, _19803_, _19793_);
  and _65297_ (_19804_, _18777_, _18616_);
  and _65298_ (_19805_, _19804_, _18981_);
  and _65299_ (_19806_, _18780_, _18503_);
  not _65300_ (_19807_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _65301_ (_19808_, _18785_, _18905_);
  nor _65302_ (_19809_, _19808_, _19807_);
  and _65303_ (_19810_, _19808_, _19096_);
  or _65304_ (_19811_, _19810_, _19809_);
  or _65305_ (_19812_, _19811_, _19806_);
  not _65306_ (_19813_, _19806_);
  or _65307_ (_19814_, _19813_, word_in[8]);
  nand _65308_ (_19815_, _19814_, _19812_);
  nor _65309_ (_19816_, _19815_, _19805_);
  and _65310_ (_19817_, _18976_, _18700_);
  and _65311_ (_19818_, _19817_, _18426_);
  and _65312_ (_19819_, _19805_, _19104_);
  or _65313_ (_19820_, _19819_, _19818_);
  or _65314_ (_19821_, _19820_, _19816_);
  not _65315_ (_19822_, _19818_);
  or _65316_ (_19823_, _19822_, _19414_);
  and _65317_ (_36841_, _19823_, _19821_);
  and _65318_ (_19824_, _19808_, word_in[1]);
  not _65319_ (_19825_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _65320_ (_19826_, _19808_, _19825_);
  nor _65321_ (_19827_, _19826_, _19824_);
  nor _65322_ (_19828_, _19827_, _19806_);
  and _65323_ (_19829_, _19806_, word_in[9]);
  nor _65324_ (_19830_, _19829_, _19828_);
  nor _65325_ (_19831_, _19830_, _19805_);
  and _65326_ (_19832_, _19805_, _19119_);
  or _65327_ (_19833_, _19832_, _19831_);
  and _65328_ (_19834_, _19833_, _19822_);
  and _65329_ (_19835_, _19818_, _19426_);
  or _65330_ (_36842_, _19835_, _19834_);
  and _65331_ (_19836_, _19808_, word_in[2]);
  not _65332_ (_19837_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _65333_ (_19838_, _19808_, _19837_);
  nor _65334_ (_19839_, _19838_, _19836_);
  nor _65335_ (_19840_, _19839_, _19806_);
  and _65336_ (_19841_, _19806_, word_in[10]);
  nor _65337_ (_19842_, _19841_, _19840_);
  nor _65338_ (_19843_, _19842_, _19805_);
  and _65339_ (_19844_, _19805_, _19132_);
  or _65340_ (_19845_, _19844_, _19843_);
  and _65341_ (_19846_, _19845_, _19822_);
  and _65342_ (_19847_, _19818_, _19439_);
  or _65343_ (_36843_, _19847_, _19846_);
  and _65344_ (_19848_, _19808_, word_in[3]);
  not _65345_ (_19849_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _65346_ (_19850_, _19808_, _19849_);
  nor _65347_ (_19851_, _19850_, _19848_);
  nor _65348_ (_19852_, _19851_, _19806_);
  and _65349_ (_19853_, _19806_, word_in[11]);
  nor _65350_ (_19854_, _19853_, _19852_);
  nor _65351_ (_19855_, _19854_, _19805_);
  and _65352_ (_19856_, _19805_, _19145_);
  or _65353_ (_19857_, _19856_, _19855_);
  and _65354_ (_19858_, _19857_, _19822_);
  and _65355_ (_19859_, _19818_, _19452_);
  or _65356_ (_36844_, _19859_, _19858_);
  not _65357_ (_19860_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _65358_ (_19861_, _19808_, _19860_);
  and _65359_ (_19862_, _19808_, _19151_);
  or _65360_ (_19863_, _19862_, _19861_);
  or _65361_ (_19864_, _19863_, _19806_);
  nand _65362_ (_19865_, _19806_, _19257_);
  nand _65363_ (_19866_, _19865_, _19864_);
  nor _65364_ (_19867_, _19866_, _19805_);
  and _65365_ (_19868_, _19805_, _19158_);
  or _65366_ (_19869_, _19868_, _19867_);
  or _65367_ (_19870_, _19869_, _19818_);
  or _65368_ (_19871_, _19822_, _19038_);
  and _65369_ (_36845_, _19871_, _19870_);
  and _65370_ (_19872_, _19808_, word_in[5]);
  not _65371_ (_19873_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _65372_ (_19874_, _19808_, _19873_);
  nor _65373_ (_19875_, _19874_, _19872_);
  nor _65374_ (_19876_, _19875_, _19806_);
  and _65375_ (_19877_, _19806_, word_in[13]);
  nor _65376_ (_19878_, _19877_, _19876_);
  nor _65377_ (_19879_, _19878_, _19805_);
  and _65378_ (_19880_, _19805_, _19171_);
  or _65379_ (_19881_, _19880_, _19879_);
  and _65380_ (_19882_, _19881_, _19822_);
  and _65381_ (_19883_, _19818_, _19479_);
  or _65382_ (_36846_, _19883_, _19882_);
  and _65383_ (_19884_, _19808_, word_in[6]);
  not _65384_ (_19885_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _65385_ (_19886_, _19808_, _19885_);
  nor _65386_ (_19887_, _19886_, _19884_);
  nor _65387_ (_19888_, _19887_, _19806_);
  and _65388_ (_19889_, _19806_, word_in[14]);
  nor _65389_ (_19890_, _19889_, _19888_);
  nor _65390_ (_19891_, _19890_, _19805_);
  and _65391_ (_19892_, _19805_, _19184_);
  or _65392_ (_19893_, _19892_, _19891_);
  and _65393_ (_19894_, _19893_, _19822_);
  and _65394_ (_19895_, _19818_, _19492_);
  or _65395_ (_36847_, _19895_, _19894_);
  and _65396_ (_19896_, _19808_, word_in[7]);
  nor _65397_ (_19897_, _19808_, _18581_);
  nor _65398_ (_19898_, _19897_, _19896_);
  nor _65399_ (_19899_, _19898_, _19806_);
  and _65400_ (_19900_, _19806_, word_in[15]);
  nor _65401_ (_19901_, _19900_, _19899_);
  nor _65402_ (_19902_, _19901_, _19805_);
  and _65403_ (_19903_, _19805_, _18795_);
  or _65404_ (_19904_, _19903_, _19902_);
  and _65405_ (_19905_, _19904_, _19822_);
  and _65406_ (_19906_, _19818_, _18768_);
  or _65407_ (_36848_, _19906_, _19905_);
  and _65408_ (_19907_, _19817_, _18437_);
  not _65409_ (_19908_, _19907_);
  and _65410_ (_19909_, _19804_, _19090_);
  and _65411_ (_19910_, _18780_, _18513_);
  and _65412_ (_19911_, _19910_, _18414_);
  and _65413_ (_19912_, _19096_, _18888_);
  not _65414_ (_19913_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _65415_ (_19914_, _18785_, _18888_);
  nor _65416_ (_19915_, _19914_, _19913_);
  nor _65417_ (_19916_, _19915_, _19912_);
  nor _65418_ (_19917_, _19916_, _19911_);
  and _65419_ (_19918_, _19911_, _19407_);
  nor _65420_ (_19919_, _19918_, _19917_);
  nor _65421_ (_19920_, _19919_, _19909_);
  and _65422_ (_19921_, _19909_, _19104_);
  or _65423_ (_19922_, _19921_, _19920_);
  and _65424_ (_19923_, _19922_, _19908_);
  and _65425_ (_19924_, _19907_, _19414_);
  or _65426_ (_36849_, _19924_, _19923_);
  not _65427_ (_19925_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _65428_ (_19926_, _19914_, _19925_);
  and _65429_ (_19927_, _19112_, _18888_);
  nor _65430_ (_19928_, _19927_, _19926_);
  nor _65431_ (_19929_, _19928_, _19911_);
  and _65432_ (_19930_, _19911_, _19001_);
  nor _65433_ (_19931_, _19930_, _19929_);
  nor _65434_ (_19932_, _19931_, _19909_);
  and _65435_ (_19933_, _19909_, _19119_);
  or _65436_ (_19934_, _19933_, _19932_);
  and _65437_ (_19935_, _19934_, _19908_);
  and _65438_ (_19936_, _19907_, _19426_);
  or _65439_ (_36850_, _19936_, _19935_);
  not _65440_ (_19937_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _65441_ (_19938_, _19914_, _19937_);
  and _65442_ (_19939_, _19125_, _18888_);
  or _65443_ (_19940_, _19939_, _19938_);
  or _65444_ (_19941_, _19940_, _19911_);
  not _65445_ (_19942_, _19911_);
  or _65446_ (_19943_, _19942_, _19432_);
  and _65447_ (_19944_, _19943_, _19941_);
  or _65448_ (_19945_, _19944_, _19909_);
  not _65449_ (_19946_, _19909_);
  or _65450_ (_19947_, _19946_, _19132_);
  and _65451_ (_19948_, _19947_, _19945_);
  or _65452_ (_19949_, _19948_, _19907_);
  or _65453_ (_19950_, _19908_, _19439_);
  and _65454_ (_36851_, _19950_, _19949_);
  not _65455_ (_19951_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _65456_ (_19952_, _19914_, _19951_);
  and _65457_ (_19953_, _19137_, _18888_);
  nor _65458_ (_19954_, _19953_, _19952_);
  nor _65459_ (_19955_, _19954_, _19911_);
  and _65460_ (_19956_, _19911_, _19445_);
  nor _65461_ (_19957_, _19956_, _19955_);
  nor _65462_ (_19958_, _19957_, _19909_);
  and _65463_ (_19959_, _19909_, _19145_);
  or _65464_ (_19960_, _19959_, _19907_);
  or _65465_ (_19961_, _19960_, _19958_);
  or _65466_ (_19962_, _19908_, _19452_);
  and _65467_ (_36852_, _19962_, _19961_);
  not _65468_ (_19963_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _65469_ (_19964_, _19914_, _19963_);
  and _65470_ (_19965_, _19151_, _18888_);
  or _65471_ (_19966_, _19965_, _19964_);
  or _65472_ (_19967_, _19966_, _19911_);
  or _65473_ (_19968_, _19942_, _19454_);
  and _65474_ (_19969_, _19968_, _19967_);
  or _65475_ (_19970_, _19969_, _19909_);
  or _65476_ (_19971_, _19946_, _19158_);
  and _65477_ (_19972_, _19971_, _19970_);
  or _65478_ (_19973_, _19972_, _19907_);
  or _65479_ (_19974_, _19908_, _19038_);
  and _65480_ (_36853_, _19974_, _19973_);
  not _65481_ (_19975_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _65482_ (_19976_, _19914_, _19975_);
  and _65483_ (_19977_, _19163_, _18888_);
  or _65484_ (_19978_, _19977_, _19976_);
  or _65485_ (_19979_, _19978_, _19911_);
  or _65486_ (_19980_, _19942_, _19472_);
  nand _65487_ (_19981_, _19980_, _19979_);
  nor _65488_ (_19982_, _19981_, _19909_);
  and _65489_ (_19983_, _19909_, _19171_);
  or _65490_ (_19984_, _19983_, _19907_);
  or _65491_ (_19985_, _19984_, _19982_);
  or _65492_ (_19986_, _19908_, _19479_);
  and _65493_ (_36854_, _19986_, _19985_);
  and _65494_ (_19987_, _19914_, word_in[6]);
  not _65495_ (_19988_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _65496_ (_19989_, _19914_, _19988_);
  nor _65497_ (_19990_, _19989_, _19987_);
  nor _65498_ (_19991_, _19990_, _19911_);
  and _65499_ (_19992_, _19911_, _19485_);
  nor _65500_ (_19993_, _19992_, _19991_);
  nor _65501_ (_19994_, _19993_, _19909_);
  and _65502_ (_19995_, _19909_, _19184_);
  or _65503_ (_19996_, _19995_, _19994_);
  and _65504_ (_19997_, _19996_, _19908_);
  and _65505_ (_19998_, _19907_, _19492_);
  or _65506_ (_36855_, _19998_, _19997_);
  nor _65507_ (_19999_, _19914_, _18472_);
  and _65508_ (_20000_, _19914_, _19189_);
  or _65509_ (_20001_, _20000_, _19999_);
  or _65510_ (_20002_, _20001_, _19911_);
  or _65511_ (_20003_, _19942_, _18791_);
  and _65512_ (_20004_, _20003_, _20002_);
  or _65513_ (_20005_, _20004_, _19909_);
  or _65514_ (_20006_, _19946_, _18795_);
  and _65515_ (_20007_, _20006_, _19908_);
  and _65516_ (_20008_, _20007_, _20005_);
  and _65517_ (_20009_, _19907_, _18768_);
  or _65518_ (_36856_, _20009_, _20008_);
  and _65519_ (_20010_, _18976_, _18499_);
  not _65520_ (_20011_, _20010_);
  and _65521_ (_20012_, _19804_, _19205_);
  and _65522_ (_20013_, _19910_, _18426_);
  and _65523_ (_20014_, _18785_, _18900_);
  and _65524_ (_20015_, _20014_, _19096_);
  not _65525_ (_20016_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor _65526_ (_20017_, _20014_, _20016_);
  nor _65527_ (_20018_, _20017_, _20015_);
  nor _65528_ (_20019_, _20018_, _20013_);
  and _65529_ (_20020_, _20013_, _19407_);
  nor _65530_ (_20021_, _20020_, _20019_);
  nor _65531_ (_20022_, _20021_, _20012_);
  and _65532_ (_20023_, _20012_, _19104_);
  or _65533_ (_20024_, _20023_, _20022_);
  and _65534_ (_20025_, _20024_, _20011_);
  and _65535_ (_20026_, _20010_, word_in[24]);
  or _65536_ (_36738_, _20026_, _20025_);
  and _65537_ (_20027_, _20014_, word_in[1]);
  not _65538_ (_20028_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _65539_ (_20029_, _20014_, _20028_);
  nor _65540_ (_20030_, _20029_, _20027_);
  nor _65541_ (_20031_, _20030_, _20013_);
  and _65542_ (_20032_, _20013_, _19001_);
  nor _65543_ (_20033_, _20032_, _20031_);
  nor _65544_ (_20034_, _20033_, _20012_);
  and _65545_ (_20035_, _20012_, _19119_);
  or _65546_ (_20036_, _20035_, _20010_);
  or _65547_ (_20037_, _20036_, _20034_);
  or _65548_ (_20038_, _20011_, _19426_);
  and _65549_ (_36739_, _20038_, _20037_);
  and _65550_ (_20039_, _20014_, word_in[2]);
  not _65551_ (_20040_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _65552_ (_20041_, _20014_, _20040_);
  nor _65553_ (_20042_, _20041_, _20039_);
  nor _65554_ (_20043_, _20042_, _20013_);
  and _65555_ (_20044_, _20013_, _19432_);
  nor _65556_ (_20045_, _20044_, _20043_);
  nor _65557_ (_20046_, _20045_, _20012_);
  and _65558_ (_20047_, _20012_, _19132_);
  or _65559_ (_20048_, _20047_, _20010_);
  or _65560_ (_20049_, _20048_, _20046_);
  or _65561_ (_20050_, _20011_, _19439_);
  and _65562_ (_36740_, _20050_, _20049_);
  and _65563_ (_20051_, _20014_, word_in[3]);
  not _65564_ (_20052_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _65565_ (_20053_, _20014_, _20052_);
  nor _65566_ (_20054_, _20053_, _20051_);
  nor _65567_ (_20055_, _20054_, _20013_);
  and _65568_ (_20056_, _20013_, _19445_);
  nor _65569_ (_20057_, _20056_, _20055_);
  nor _65570_ (_20058_, _20057_, _20012_);
  and _65571_ (_20059_, _20012_, _19145_);
  or _65572_ (_20060_, _20059_, _20058_);
  and _65573_ (_20061_, _20060_, _20011_);
  and _65574_ (_20062_, _20010_, word_in[27]);
  or _65575_ (_36741_, _20062_, _20061_);
  and _65576_ (_20063_, _20014_, word_in[4]);
  not _65577_ (_20064_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor _65578_ (_20065_, _20014_, _20064_);
  nor _65579_ (_20066_, _20065_, _20063_);
  nor _65580_ (_20067_, _20066_, _20013_);
  and _65581_ (_20068_, _20013_, _19454_);
  nor _65582_ (_20069_, _20068_, _20067_);
  nor _65583_ (_20070_, _20069_, _20012_);
  and _65584_ (_20071_, _20012_, _19158_);
  or _65585_ (_20072_, _20071_, _20070_);
  and _65586_ (_20073_, _20072_, _20011_);
  and _65587_ (_20074_, _20010_, word_in[28]);
  or _65588_ (_36742_, _20074_, _20073_);
  and _65589_ (_20075_, _20014_, word_in[5]);
  not _65590_ (_20076_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _65591_ (_20077_, _20014_, _20076_);
  nor _65592_ (_20078_, _20077_, _20075_);
  nor _65593_ (_20079_, _20078_, _20013_);
  and _65594_ (_20080_, _20013_, _19472_);
  nor _65595_ (_20081_, _20080_, _20079_);
  nor _65596_ (_20082_, _20081_, _20012_);
  and _65597_ (_20083_, _20012_, _19171_);
  or _65598_ (_20084_, _20083_, _20082_);
  and _65599_ (_20085_, _20084_, _20011_);
  and _65600_ (_20086_, _20010_, word_in[29]);
  or _65601_ (_36743_, _20086_, _20085_);
  not _65602_ (_20087_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _65603_ (_20088_, _20014_, _20087_);
  and _65604_ (_20089_, _20014_, word_in[6]);
  nor _65605_ (_20090_, _20089_, _20088_);
  nor _65606_ (_20091_, _20090_, _20013_);
  and _65607_ (_20092_, _20013_, _19485_);
  nor _65608_ (_20093_, _20092_, _20091_);
  nor _65609_ (_20094_, _20093_, _20012_);
  and _65610_ (_20095_, _20012_, _19184_);
  or _65611_ (_20096_, _20095_, _20094_);
  and _65612_ (_20097_, _20096_, _20011_);
  and _65613_ (_20098_, _20010_, word_in[30]);
  or _65614_ (_36744_, _20098_, _20097_);
  and _65615_ (_20099_, _20014_, word_in[7]);
  nor _65616_ (_20100_, _20014_, _18586_);
  nor _65617_ (_20101_, _20100_, _20099_);
  nor _65618_ (_20102_, _20101_, _20013_);
  and _65619_ (_20103_, _20013_, _18791_);
  nor _65620_ (_20104_, _20103_, _20102_);
  nor _65621_ (_20105_, _20104_, _20012_);
  and _65622_ (_20106_, _20012_, _18795_);
  or _65623_ (_20107_, _20106_, _20010_);
  or _65624_ (_20108_, _20107_, _20105_);
  or _65625_ (_20109_, _20011_, _18768_);
  and _65626_ (_36745_, _20109_, _20108_);
  and _65627_ (_20110_, _18767_, _18905_);
  not _65628_ (_20111_, _20110_);
  and _65629_ (_20112_, _19804_, _18774_);
  and _65630_ (_20113_, _19910_, _18437_);
  and _65631_ (_20114_, _18785_, _18926_);
  and _65632_ (_20115_, _20114_, word_in[0]);
  not _65633_ (_20116_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor _65634_ (_20117_, _20114_, _20116_);
  nor _65635_ (_20118_, _20117_, _20115_);
  nor _65636_ (_20119_, _20118_, _20113_);
  and _65637_ (_20120_, _20113_, _19407_);
  nor _65638_ (_20121_, _20120_, _20119_);
  nor _65639_ (_20122_, _20121_, _20112_);
  and _65640_ (_20123_, _20112_, _19104_);
  or _65641_ (_20124_, _20123_, _20122_);
  and _65642_ (_20125_, _20124_, _20111_);
  and _65643_ (_20126_, _20110_, word_in[24]);
  or _65644_ (_36746_, _20126_, _20125_);
  not _65645_ (_20127_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _65646_ (_20128_, _20114_, _20127_);
  and _65647_ (_20129_, _20114_, word_in[1]);
  or _65648_ (_20130_, _20129_, _20128_);
  or _65649_ (_20131_, _20130_, _20113_);
  not _65650_ (_20132_, _20113_);
  or _65651_ (_20133_, _20132_, _19001_);
  and _65652_ (_20134_, _20133_, _20131_);
  or _65653_ (_20135_, _20134_, _20112_);
  not _65654_ (_20136_, _20112_);
  or _65655_ (_20137_, _20136_, _19119_);
  and _65656_ (_20138_, _20137_, _20111_);
  and _65657_ (_20139_, _20138_, _20135_);
  and _65658_ (_20140_, _20110_, word_in[25]);
  or _65659_ (_36747_, _20140_, _20139_);
  and _65660_ (_20141_, _20114_, word_in[2]);
  not _65661_ (_20142_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _65662_ (_20143_, _20114_, _20142_);
  nor _65663_ (_20144_, _20143_, _20141_);
  nor _65664_ (_20145_, _20144_, _20113_);
  and _65665_ (_20146_, _20113_, _19432_);
  nor _65666_ (_20147_, _20146_, _20145_);
  nor _65667_ (_20148_, _20147_, _20112_);
  and _65668_ (_20149_, _20112_, _19132_);
  or _65669_ (_20150_, _20149_, _20148_);
  and _65670_ (_20151_, _20150_, _20111_);
  and _65671_ (_20152_, _20110_, word_in[26]);
  or _65672_ (_36748_, _20152_, _20151_);
  and _65673_ (_20153_, _20114_, word_in[3]);
  not _65674_ (_20154_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _65675_ (_20155_, _20114_, _20154_);
  nor _65676_ (_20156_, _20155_, _20153_);
  nor _65677_ (_20157_, _20156_, _20113_);
  and _65678_ (_20158_, _20113_, _19445_);
  nor _65679_ (_20159_, _20158_, _20157_);
  nor _65680_ (_20160_, _20159_, _20112_);
  and _65681_ (_20161_, _20112_, _19145_);
  or _65682_ (_20162_, _20161_, _20160_);
  and _65683_ (_20163_, _20162_, _20111_);
  and _65684_ (_20164_, _20110_, word_in[27]);
  or _65685_ (_36749_, _20164_, _20163_);
  not _65686_ (_20165_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _65687_ (_20166_, _20114_, _20165_);
  and _65688_ (_20167_, _20114_, word_in[4]);
  or _65689_ (_20168_, _20167_, _20166_);
  or _65690_ (_20169_, _20168_, _20113_);
  or _65691_ (_20170_, _20132_, _19454_);
  and _65692_ (_20171_, _20170_, _20169_);
  or _65693_ (_20172_, _20171_, _20112_);
  or _65694_ (_20173_, _20136_, _19158_);
  and _65695_ (_20174_, _20173_, _20111_);
  and _65696_ (_20175_, _20174_, _20172_);
  and _65697_ (_20176_, _20110_, word_in[28]);
  or _65698_ (_36750_, _20176_, _20175_);
  and _65699_ (_20177_, _20114_, word_in[5]);
  not _65700_ (_20178_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _65701_ (_20179_, _20114_, _20178_);
  nor _65702_ (_20180_, _20179_, _20177_);
  nor _65703_ (_20181_, _20180_, _20113_);
  and _65704_ (_20182_, _20113_, _19472_);
  nor _65705_ (_20183_, _20182_, _20181_);
  nor _65706_ (_20184_, _20183_, _20112_);
  and _65707_ (_20185_, _20112_, _19171_);
  or _65708_ (_20186_, _20185_, _20184_);
  and _65709_ (_20187_, _20186_, _20111_);
  and _65710_ (_20188_, _20110_, word_in[29]);
  or _65711_ (_36751_, _20188_, _20187_);
  and _65712_ (_20189_, _20114_, word_in[6]);
  not _65713_ (_20190_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _65714_ (_20191_, _20114_, _20190_);
  nor _65715_ (_20192_, _20191_, _20189_);
  nor _65716_ (_20193_, _20192_, _20113_);
  and _65717_ (_20194_, _20113_, _19485_);
  nor _65718_ (_20195_, _20194_, _20193_);
  nor _65719_ (_20196_, _20195_, _20112_);
  and _65720_ (_20197_, _20112_, _19184_);
  or _65721_ (_20198_, _20197_, _20196_);
  and _65722_ (_20199_, _20198_, _20111_);
  and _65723_ (_20200_, _20110_, word_in[30]);
  or _65724_ (_36752_, _20200_, _20199_);
  nor _65725_ (_20201_, _20114_, _18489_);
  and _65726_ (_20202_, _20114_, word_in[7]);
  or _65727_ (_20203_, _20202_, _20201_);
  or _65728_ (_20204_, _20203_, _20113_);
  or _65729_ (_20205_, _20132_, _18791_);
  and _65730_ (_20206_, _20205_, _20204_);
  or _65731_ (_20207_, _20206_, _20112_);
  or _65732_ (_20208_, _20136_, _18795_);
  and _65733_ (_20209_, _20208_, _20111_);
  and _65734_ (_20210_, _20209_, _20207_);
  and _65735_ (_20211_, _20110_, word_in[31]);
  or _65736_ (_36753_, _20211_, _20210_);
  and _65737_ (_20212_, _18975_, _18695_);
  and _65738_ (_20213_, _20212_, _18426_);
  and _65739_ (_20214_, _18981_, _18778_);
  and _65740_ (_20215_, _18780_, _18926_);
  and _65741_ (_20216_, _18785_, _18769_);
  and _65742_ (_20217_, _20216_, _19096_);
  not _65743_ (_20218_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _65744_ (_20219_, _20216_, _20218_);
  or _65745_ (_20220_, _20219_, _20217_);
  or _65746_ (_20221_, _20220_, _20215_);
  not _65747_ (_20222_, _20215_);
  or _65748_ (_20223_, _20222_, word_in[8]);
  and _65749_ (_20224_, _20223_, _20221_);
  or _65750_ (_20225_, _20224_, _20214_);
  not _65751_ (_20226_, _20214_);
  or _65752_ (_20227_, _20226_, _19104_);
  and _65753_ (_20228_, _20227_, _20225_);
  or _65754_ (_20229_, _20228_, _20213_);
  not _65755_ (_20230_, _20213_);
  or _65756_ (_20231_, _20230_, word_in[24]);
  and _65757_ (_36754_, _20231_, _20229_);
  not _65758_ (_20232_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _65759_ (_20233_, _20216_, _20232_);
  and _65760_ (_20234_, _20216_, _19112_);
  nor _65761_ (_20235_, _20234_, _20233_);
  nor _65762_ (_20236_, _20235_, _20215_);
  and _65763_ (_20237_, _20215_, word_in[9]);
  nor _65764_ (_20238_, _20237_, _20236_);
  nor _65765_ (_20239_, _20238_, _20214_);
  and _65766_ (_20240_, _20214_, _19119_);
  or _65767_ (_20241_, _20240_, _20239_);
  and _65768_ (_20242_, _20241_, _20230_);
  and _65769_ (_20243_, _20213_, word_in[25]);
  or _65770_ (_36755_, _20243_, _20242_);
  and _65771_ (_20244_, _20216_, _19125_);
  not _65772_ (_20245_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _65773_ (_20246_, _20216_, _20245_);
  nor _65774_ (_20247_, _20246_, _20244_);
  nor _65775_ (_20248_, _20247_, _20215_);
  and _65776_ (_20249_, _20215_, word_in[10]);
  nor _65777_ (_20250_, _20249_, _20248_);
  nor _65778_ (_20251_, _20250_, _20214_);
  and _65779_ (_20252_, _20214_, _19132_);
  or _65780_ (_20253_, _20252_, _20251_);
  and _65781_ (_20254_, _20253_, _20230_);
  and _65782_ (_20255_, _20213_, word_in[26]);
  or _65783_ (_36756_, _20255_, _20254_);
  and _65784_ (_20256_, _20216_, word_in[3]);
  not _65785_ (_20257_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _65786_ (_20258_, _20216_, _20257_);
  nor _65787_ (_20259_, _20258_, _20256_);
  nor _65788_ (_20260_, _20259_, _20215_);
  and _65789_ (_20261_, _20215_, word_in[11]);
  nor _65790_ (_20262_, _20261_, _20260_);
  nor _65791_ (_20263_, _20262_, _20214_);
  and _65792_ (_20264_, _20214_, _19145_);
  or _65793_ (_20265_, _20264_, _20263_);
  and _65794_ (_20266_, _20265_, _20230_);
  and _65795_ (_20267_, _20213_, word_in[27]);
  or _65796_ (_36757_, _20267_, _20266_);
  and _65797_ (_20268_, _20216_, word_in[4]);
  not _65798_ (_20269_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _65799_ (_20270_, _20216_, _20269_);
  nor _65800_ (_20271_, _20270_, _20268_);
  nor _65801_ (_20272_, _20271_, _20215_);
  and _65802_ (_20273_, _20215_, word_in[12]);
  nor _65803_ (_20274_, _20273_, _20272_);
  nor _65804_ (_20275_, _20274_, _20214_);
  and _65805_ (_20276_, _20214_, _19158_);
  or _65806_ (_20277_, _20276_, _20275_);
  and _65807_ (_20278_, _20277_, _20230_);
  and _65808_ (_20279_, _20213_, word_in[28]);
  or _65809_ (_36758_, _20279_, _20278_);
  and _65810_ (_20280_, _20216_, word_in[5]);
  not _65811_ (_20281_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _65812_ (_20282_, _20216_, _20281_);
  nor _65813_ (_20283_, _20282_, _20280_);
  nor _65814_ (_20284_, _20283_, _20215_);
  and _65815_ (_20285_, _20215_, word_in[13]);
  nor _65816_ (_20286_, _20285_, _20284_);
  nor _65817_ (_20287_, _20286_, _20214_);
  and _65818_ (_20288_, _20214_, _19171_);
  or _65819_ (_20289_, _20288_, _20287_);
  and _65820_ (_20290_, _20289_, _20230_);
  and _65821_ (_20291_, _20213_, word_in[29]);
  or _65822_ (_36759_, _20291_, _20290_);
  not _65823_ (_20292_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _65824_ (_20293_, _20216_, _20292_);
  and _65825_ (_20294_, _20216_, _19177_);
  or _65826_ (_20295_, _20294_, _20293_);
  or _65827_ (_20296_, _20295_, _20215_);
  or _65828_ (_20297_, _20222_, word_in[14]);
  and _65829_ (_20298_, _20297_, _20296_);
  or _65830_ (_20299_, _20298_, _20214_);
  or _65831_ (_20300_, _20226_, _19184_);
  and _65832_ (_20301_, _20300_, _20299_);
  or _65833_ (_20302_, _20301_, _20213_);
  or _65834_ (_20303_, _20230_, word_in[30]);
  and _65835_ (_36760_, _20303_, _20302_);
  and _65836_ (_20304_, _20216_, word_in[7]);
  nor _65837_ (_20305_, _20216_, _18593_);
  nor _65838_ (_20306_, _20305_, _20304_);
  nor _65839_ (_20307_, _20306_, _20215_);
  and _65840_ (_20308_, _20215_, word_in[15]);
  nor _65841_ (_20309_, _20308_, _20307_);
  nor _65842_ (_20310_, _20309_, _20214_);
  and _65843_ (_20311_, _20214_, _18795_);
  or _65844_ (_20312_, _20311_, _20310_);
  and _65845_ (_20313_, _20312_, _20230_);
  and _65846_ (_20314_, _20213_, word_in[31]);
  or _65847_ (_36761_, _20314_, _20313_);
  and _65848_ (_20315_, _20212_, _18437_);
  and _65849_ (_20316_, _19090_, _18778_);
  and _65850_ (_20317_, _18782_, _18414_);
  not _65851_ (_20318_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _65852_ (_20319_, _18785_, _18966_);
  nor _65853_ (_20320_, _20319_, _20318_);
  and _65854_ (_20321_, _19096_, _18966_);
  or _65855_ (_20322_, _20321_, _20320_);
  or _65856_ (_20323_, _20322_, _20317_);
  not _65857_ (_20324_, _20317_);
  or _65858_ (_20325_, _20324_, _19407_);
  and _65859_ (_20326_, _20325_, _20323_);
  or _65860_ (_20327_, _20326_, _20316_);
  not _65861_ (_20328_, _20316_);
  or _65862_ (_20329_, _20328_, _19104_);
  and _65863_ (_20330_, _20329_, _20327_);
  or _65864_ (_20331_, _20330_, _20315_);
  not _65865_ (_20332_, _20315_);
  or _65866_ (_20333_, _20332_, _19414_);
  and _65867_ (_36762_, _20333_, _20331_);
  not _65868_ (_20334_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _65869_ (_20335_, _20319_, _20334_);
  and _65870_ (_20336_, _19112_, _18966_);
  nor _65871_ (_20337_, _20336_, _20335_);
  nor _65872_ (_20338_, _20337_, _20317_);
  and _65873_ (_20339_, _20317_, _19001_);
  or _65874_ (_20340_, _20339_, _20338_);
  or _65875_ (_20341_, _20340_, _20316_);
  or _65876_ (_20342_, _20328_, _19119_);
  and _65877_ (_20343_, _20342_, _20332_);
  and _65878_ (_20344_, _20343_, _20341_);
  and _65879_ (_20345_, _20315_, _19426_);
  or _65880_ (_36763_, _20345_, _20344_);
  not _65881_ (_20346_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _65882_ (_20347_, _20319_, _20346_);
  and _65883_ (_20348_, _19125_, _18966_);
  or _65884_ (_20349_, _20348_, _20347_);
  or _65885_ (_20350_, _20349_, _20317_);
  or _65886_ (_20351_, _20324_, _19432_);
  and _65887_ (_20352_, _20351_, _20350_);
  or _65888_ (_20353_, _20352_, _20316_);
  or _65889_ (_20354_, _20328_, _19132_);
  and _65890_ (_20355_, _20354_, _20353_);
  or _65891_ (_20356_, _20355_, _20315_);
  or _65892_ (_20357_, _20332_, _19439_);
  and _65893_ (_36764_, _20357_, _20356_);
  or _65894_ (_20358_, _20324_, _19445_);
  not _65895_ (_20359_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _65896_ (_20360_, _20319_, _20359_);
  and _65897_ (_20361_, _20319_, word_in[3]);
  or _65898_ (_20362_, _20361_, _20360_);
  or _65899_ (_20363_, _20362_, _20317_);
  and _65900_ (_20364_, _20363_, _20358_);
  or _65901_ (_20365_, _20364_, _20316_);
  or _65902_ (_20366_, _20328_, _19145_);
  and _65903_ (_20367_, _20366_, _20365_);
  or _65904_ (_20368_, _20367_, _20315_);
  or _65905_ (_20369_, _20332_, _19452_);
  and _65906_ (_36765_, _20369_, _20368_);
  or _65907_ (_20370_, _20324_, _19454_);
  and _65908_ (_20371_, _20319_, word_in[4]);
  not _65909_ (_20372_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _65910_ (_20373_, _20319_, _20372_);
  or _65911_ (_20374_, _20373_, _20371_);
  or _65912_ (_20375_, _20374_, _20317_);
  and _65913_ (_20376_, _20375_, _20370_);
  or _65914_ (_20377_, _20376_, _20316_);
  or _65915_ (_20378_, _20328_, _19158_);
  and _65916_ (_20379_, _20378_, _20332_);
  and _65917_ (_20380_, _20379_, _20377_);
  and _65918_ (_20381_, _20315_, _19038_);
  or _65919_ (_36766_, _20381_, _20380_);
  not _65920_ (_20382_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _65921_ (_20383_, _20319_, _20382_);
  and _65922_ (_20384_, _20319_, _19163_);
  or _65923_ (_20385_, _20384_, _20383_);
  or _65924_ (_20386_, _20385_, _20317_);
  or _65925_ (_20387_, _20324_, _19472_);
  and _65926_ (_20388_, _20387_, _20386_);
  or _65927_ (_20389_, _20388_, _20316_);
  or _65928_ (_20390_, _20328_, _19171_);
  and _65929_ (_20391_, _20390_, _20332_);
  and _65930_ (_20392_, _20391_, _20389_);
  and _65931_ (_20393_, _20315_, _19479_);
  or _65932_ (_36767_, _20393_, _20392_);
  and _65933_ (_20394_, _20317_, _19485_);
  not _65934_ (_20395_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  or _65935_ (_20396_, _20319_, _20395_);
  nand _65936_ (_20397_, _20319_, _19177_);
  and _65937_ (_20398_, _20397_, _20396_);
  nor _65938_ (_20399_, _20398_, _20317_);
  nor _65939_ (_20400_, _20399_, _20394_);
  nor _65940_ (_20401_, _20400_, _20316_);
  and _65941_ (_20402_, _20316_, _19184_);
  or _65942_ (_20403_, _20402_, _20401_);
  and _65943_ (_20404_, _20403_, _20332_);
  and _65944_ (_20405_, _20315_, _19492_);
  or _65945_ (_36768_, _20405_, _20404_);
  nor _65946_ (_20406_, _20319_, _18478_);
  and _65947_ (_20407_, _20319_, _19189_);
  or _65948_ (_20408_, _20407_, _20406_);
  or _65949_ (_20409_, _20408_, _20317_);
  or _65950_ (_20410_, _20324_, _18791_);
  and _65951_ (_20411_, _20410_, _20409_);
  or _65952_ (_20412_, _20411_, _20316_);
  or _65953_ (_20413_, _20328_, _18795_);
  and _65954_ (_20414_, _20413_, _20332_);
  and _65955_ (_20415_, _20414_, _20412_);
  and _65956_ (_20416_, _20315_, _18768_);
  or _65957_ (_36769_, _20416_, _20415_);
  and _65958_ (_20417_, _20212_, _18404_);
  and _65959_ (_20418_, _19205_, _18778_);
  and _65960_ (_20419_, _18782_, _18426_);
  not _65961_ (_20420_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _65962_ (_20421_, _18785_, _18804_);
  nor _65963_ (_20422_, _20421_, _20420_);
  and _65964_ (_20423_, _20421_, _19096_);
  or _65965_ (_20424_, _20423_, _20422_);
  or _65966_ (_20425_, _20424_, _20419_);
  not _65967_ (_20426_, _20419_);
  or _65968_ (_20427_, _20426_, _19407_);
  and _65969_ (_20428_, _20427_, _20425_);
  or _65970_ (_20429_, _20428_, _20418_);
  not _65971_ (_20430_, _20418_);
  or _65972_ (_20431_, _20430_, _19104_);
  and _65973_ (_20432_, _20431_, _20429_);
  or _65974_ (_20433_, _20432_, _20417_);
  not _65975_ (_20434_, _20417_);
  or _65976_ (_20435_, _20434_, word_in[24]);
  and _65977_ (_36770_, _20435_, _20433_);
  or _65978_ (_20436_, _20426_, _19001_);
  and _65979_ (_20437_, _20421_, word_in[1]);
  not _65980_ (_20438_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor _65981_ (_20439_, _20421_, _20438_);
  or _65982_ (_20440_, _20439_, _20437_);
  or _65983_ (_20441_, _20440_, _20419_);
  and _65984_ (_20442_, _20441_, _20436_);
  or _65985_ (_20443_, _20442_, _20418_);
  or _65986_ (_20444_, _20430_, _19119_);
  and _65987_ (_20445_, _20444_, _20443_);
  or _65988_ (_20446_, _20445_, _20417_);
  or _65989_ (_20447_, _20434_, word_in[25]);
  and _65990_ (_36771_, _20447_, _20446_);
  or _65991_ (_20448_, _20426_, _19432_);
  and _65992_ (_20449_, _20421_, word_in[2]);
  not _65993_ (_20450_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor _65994_ (_20451_, _20421_, _20450_);
  or _65995_ (_20452_, _20451_, _20449_);
  or _65996_ (_20453_, _20452_, _20419_);
  and _65997_ (_20454_, _20453_, _20448_);
  or _65998_ (_20455_, _20454_, _20418_);
  or _65999_ (_20456_, _20430_, _19132_);
  and _66000_ (_20457_, _20456_, _20434_);
  and _66001_ (_20458_, _20457_, _20455_);
  and _66002_ (_20459_, _20417_, _19439_);
  or _66003_ (_36772_, _20459_, _20458_);
  and _66004_ (_20460_, _20418_, _19145_);
  not _66005_ (_20461_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor _66006_ (_20462_, _20421_, _20461_);
  and _66007_ (_20463_, _20421_, word_in[3]);
  nor _66008_ (_20464_, _20463_, _20462_);
  nor _66009_ (_20465_, _20464_, _20419_);
  and _66010_ (_20466_, _20419_, _19445_);
  nor _66011_ (_20467_, _20466_, _20465_);
  nor _66012_ (_20468_, _20467_, _20418_);
  or _66013_ (_20469_, _20468_, _20460_);
  and _66014_ (_20470_, _20469_, _20434_);
  and _66015_ (_20471_, _20417_, word_in[27]);
  or _66016_ (_36773_, _20471_, _20470_);
  or _66017_ (_20472_, _20430_, _19158_);
  not _66018_ (_20473_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor _66019_ (_20474_, _20421_, _20473_);
  and _66020_ (_20475_, _20421_, _19151_);
  or _66021_ (_20476_, _20475_, _20474_);
  or _66022_ (_20477_, _20476_, _20419_);
  or _66023_ (_20478_, _20426_, _19454_);
  and _66024_ (_20479_, _20478_, _20477_);
  or _66025_ (_20480_, _20479_, _20418_);
  and _66026_ (_20481_, _20480_, _20472_);
  or _66027_ (_20482_, _20481_, _20417_);
  or _66028_ (_20483_, _20434_, word_in[28]);
  and _66029_ (_36774_, _20483_, _20482_);
  or _66030_ (_20484_, _20426_, _19472_);
  and _66031_ (_20485_, _20421_, word_in[5]);
  not _66032_ (_20486_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor _66033_ (_20487_, _20421_, _20486_);
  or _66034_ (_20488_, _20487_, _20485_);
  or _66035_ (_20489_, _20488_, _20419_);
  and _66036_ (_20490_, _20489_, _20484_);
  or _66037_ (_20491_, _20490_, _20418_);
  or _66038_ (_20492_, _20430_, _19171_);
  and _66039_ (_20493_, _20492_, _20434_);
  and _66040_ (_20494_, _20493_, _20491_);
  and _66041_ (_20495_, _20417_, _19479_);
  or _66042_ (_36775_, _20495_, _20494_);
  or _66043_ (_20496_, _20426_, _19485_);
  and _66044_ (_20497_, _20421_, word_in[6]);
  not _66045_ (_20498_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor _66046_ (_20499_, _20421_, _20498_);
  or _66047_ (_20500_, _20499_, _20497_);
  or _66048_ (_20501_, _20500_, _20419_);
  and _66049_ (_20502_, _20501_, _20496_);
  or _66050_ (_20503_, _20502_, _20418_);
  or _66051_ (_20504_, _20430_, _19184_);
  and _66052_ (_20505_, _20504_, _20503_);
  or _66053_ (_20506_, _20505_, _20417_);
  or _66054_ (_20507_, _20434_, word_in[30]);
  and _66055_ (_36776_, _20507_, _20506_);
  and _66056_ (_20508_, _20421_, word_in[7]);
  nor _66057_ (_20509_, _20421_, _18598_);
  nor _66058_ (_20510_, _20509_, _20508_);
  nor _66059_ (_20511_, _20510_, _20419_);
  and _66060_ (_20512_, _20419_, _18791_);
  nor _66061_ (_20513_, _20512_, _20511_);
  nor _66062_ (_20514_, _20513_, _20418_);
  and _66063_ (_20515_, _20418_, _18795_);
  or _66064_ (_20516_, _20515_, _20514_);
  and _66065_ (_20517_, _20516_, _20434_);
  and _66066_ (_20518_, _20417_, word_in[31]);
  or _66067_ (_36777_, _20518_, _20517_);
  and _66068_ (_20519_, _19414_, _18770_);
  and _66069_ (_20520_, _18786_, word_in[0]);
  not _66070_ (_20521_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor _66071_ (_20522_, _18786_, _20521_);
  nor _66072_ (_20523_, _20522_, _20520_);
  nor _66073_ (_20524_, _20523_, _18783_);
  and _66074_ (_20525_, _19407_, _18783_);
  nor _66075_ (_20526_, _20525_, _20524_);
  nor _66076_ (_20527_, _20526_, _18779_);
  and _66077_ (_20528_, _19104_, _18779_);
  or _66078_ (_20529_, _20528_, _20527_);
  and _66079_ (_20530_, _20529_, _18772_);
  or _66080_ (_36778_, _20530_, _20519_);
  not _66081_ (_20531_, _18783_);
  or _66082_ (_20532_, _19001_, _20531_);
  and _66083_ (_20533_, _18786_, word_in[1]);
  not _66084_ (_20534_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor _66085_ (_20535_, _18786_, _20534_);
  or _66086_ (_20536_, _20535_, _20533_);
  or _66087_ (_20537_, _20536_, _18783_);
  and _66088_ (_20538_, _20537_, _20532_);
  or _66089_ (_20539_, _20538_, _18779_);
  not _66090_ (_20540_, _18779_);
  or _66091_ (_20541_, _19119_, _20540_);
  and _66092_ (_20542_, _20541_, _18772_);
  and _66093_ (_20543_, _20542_, _20539_);
  and _66094_ (_20544_, _19426_, _18770_);
  or _66095_ (_36779_, _20544_, _20543_);
  and _66096_ (_20545_, _19439_, _18770_);
  and _66097_ (_20546_, _18786_, word_in[2]);
  not _66098_ (_20547_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _66099_ (_20548_, _18786_, _20547_);
  nor _66100_ (_20549_, _20548_, _20546_);
  nor _66101_ (_20550_, _20549_, _18783_);
  and _66102_ (_20551_, _19432_, _18783_);
  nor _66103_ (_20552_, _20551_, _20550_);
  nor _66104_ (_20553_, _20552_, _18779_);
  and _66105_ (_20554_, _19132_, _18779_);
  or _66106_ (_20555_, _20554_, _20553_);
  and _66107_ (_20556_, _20555_, _18772_);
  or _66108_ (_36780_, _20556_, _20545_);
  or _66109_ (_20557_, _19445_, _20531_);
  and _66110_ (_20558_, _18786_, word_in[3]);
  not _66111_ (_20559_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor _66112_ (_20560_, _18786_, _20559_);
  or _66113_ (_20561_, _20560_, _20558_);
  or _66114_ (_20562_, _20561_, _18783_);
  and _66115_ (_20563_, _20562_, _20557_);
  or _66116_ (_20564_, _20563_, _18779_);
  or _66117_ (_20565_, _19145_, _20540_);
  and _66118_ (_20566_, _20565_, _20564_);
  or _66119_ (_20567_, _20566_, _18770_);
  or _66120_ (_20568_, _18772_, word_in[27]);
  and _66121_ (_36781_, _20568_, _20567_);
  and _66122_ (_20569_, _19038_, _18770_);
  and _66123_ (_20570_, _18786_, word_in[4]);
  not _66124_ (_20571_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor _66125_ (_20572_, _18786_, _20571_);
  nor _66126_ (_20573_, _20572_, _20570_);
  nor _66127_ (_20574_, _20573_, _18783_);
  and _66128_ (_20575_, _19454_, _18783_);
  nor _66129_ (_20576_, _20575_, _20574_);
  nor _66130_ (_20577_, _20576_, _18779_);
  and _66131_ (_20578_, _19158_, _18779_);
  or _66132_ (_20579_, _20578_, _20577_);
  and _66133_ (_20580_, _20579_, _18772_);
  or _66134_ (_36782_, _20580_, _20569_);
  and _66135_ (_20581_, _18770_, word_in[29]);
  or _66136_ (_20582_, _19472_, _20531_);
  and _66137_ (_20583_, _18786_, word_in[5]);
  not _66138_ (_20584_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor _66139_ (_20585_, _18786_, _20584_);
  or _66140_ (_20586_, _20585_, _20583_);
  or _66141_ (_20587_, _20586_, _18783_);
  and _66142_ (_20588_, _20587_, _20582_);
  or _66143_ (_20589_, _20588_, _18779_);
  or _66144_ (_20590_, _19171_, _20540_);
  and _66145_ (_20591_, _20590_, _18772_);
  and _66146_ (_20592_, _20591_, _20589_);
  or _66147_ (_36783_, _20592_, _20581_);
  not _66148_ (_20593_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor _66149_ (_20594_, _18786_, _20593_);
  and _66150_ (_20595_, _19177_, _18786_);
  or _66151_ (_20596_, _20595_, _20594_);
  or _66152_ (_20597_, _20596_, _18783_);
  or _66153_ (_20598_, _19485_, _20531_);
  and _66154_ (_20599_, _20598_, _20597_);
  or _66155_ (_20600_, _20599_, _18779_);
  or _66156_ (_20601_, _19184_, _20540_);
  and _66157_ (_20602_, _20601_, _18772_);
  and _66158_ (_20603_, _20602_, _20600_);
  and _66159_ (_20604_, _18770_, word_in[30]);
  or _66160_ (_36784_, _20604_, _20603_);
  and _66161_ (_20605_, _18441_, word_in[0]);
  not _66162_ (_20606_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand _66163_ (_20607_, _18400_, _20606_);
  or _66164_ (_20608_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _66165_ (_20609_, _20608_, _20607_);
  and _66166_ (_20610_, _20609_, _18447_);
  nor _66167_ (_20611_, _20610_, _18385_);
  not _66168_ (_20612_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nand _66169_ (_20613_, _18400_, _20612_);
  or _66170_ (_20614_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _66171_ (_20615_, _20614_, _20613_);
  and _66172_ (_20616_, _20615_, _18456_);
  nand _66173_ (_20617_, _18400_, _19705_);
  or _66174_ (_20618_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _66175_ (_20619_, _20618_, _20617_);
  and _66176_ (_20620_, _20619_, _18450_);
  not _66177_ (_20621_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand _66178_ (_20622_, _18400_, _20621_);
  or _66179_ (_20623_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _66180_ (_20624_, _20623_, _20622_);
  and _66181_ (_20625_, _20624_, _18466_);
  or _66182_ (_20626_, _20625_, _20620_);
  nor _66183_ (_20627_, _20626_, _20616_);
  and _66184_ (_20628_, _20627_, _20611_);
  nand _66185_ (_20629_, _18400_, _19913_);
  or _66186_ (_20630_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _66187_ (_20631_, _20630_, _20629_);
  and _66188_ (_20632_, _20631_, _18447_);
  nor _66189_ (_20633_, _20632_, _18471_);
  nand _66190_ (_20634_, _18400_, _20318_);
  or _66191_ (_20635_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _66192_ (_20636_, _20635_, _20634_);
  and _66193_ (_20637_, _20636_, _18456_);
  nand _66194_ (_20638_, _18400_, _20521_);
  or _66195_ (_20639_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _66196_ (_20640_, _20639_, _20638_);
  and _66197_ (_20641_, _20640_, _18450_);
  nand _66198_ (_20642_, _18400_, _20116_);
  or _66199_ (_20643_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _66200_ (_20644_, _20643_, _20642_);
  and _66201_ (_20645_, _20644_, _18466_);
  or _66202_ (_20646_, _20645_, _20641_);
  nor _66203_ (_20647_, _20646_, _20637_);
  and _66204_ (_20648_, _20647_, _20633_);
  or _66205_ (_20649_, _20648_, _20628_);
  nor _66206_ (_20650_, _20649_, _18441_);
  or _66207_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _20650_, _20605_);
  and _66208_ (_20651_, _18441_, word_in[1]);
  not _66209_ (_20652_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nand _66210_ (_20653_, _18400_, _20652_);
  or _66211_ (_20654_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _66212_ (_20655_, _20654_, _20653_);
  and _66213_ (_20656_, _20655_, _18447_);
  nor _66214_ (_20657_, _20656_, _18385_);
  not _66215_ (_20658_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nand _66216_ (_20659_, _18400_, _20658_);
  or _66217_ (_20660_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _66218_ (_20661_, _20660_, _20659_);
  and _66219_ (_20662_, _20661_, _18456_);
  nand _66220_ (_20663_, _18400_, _19721_);
  or _66221_ (_20664_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _66222_ (_20665_, _20664_, _20663_);
  and _66223_ (_20666_, _20665_, _18450_);
  not _66224_ (_20667_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nand _66225_ (_20668_, _18400_, _20667_);
  or _66226_ (_20669_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _66227_ (_20670_, _20669_, _20668_);
  and _66228_ (_20671_, _20670_, _18466_);
  or _66229_ (_20672_, _20671_, _20666_);
  nor _66230_ (_20673_, _20672_, _20662_);
  and _66231_ (_20674_, _20673_, _20657_);
  nand _66232_ (_20675_, _18400_, _19925_);
  or _66233_ (_20676_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _66234_ (_20677_, _20676_, _20675_);
  and _66235_ (_20678_, _20677_, _18447_);
  nor _66236_ (_20679_, _20678_, _18471_);
  nand _66237_ (_20680_, _18400_, _20334_);
  or _66238_ (_20681_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _66239_ (_20682_, _20681_, _20680_);
  and _66240_ (_20683_, _20682_, _18456_);
  nand _66241_ (_20684_, _18400_, _20534_);
  or _66242_ (_20685_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _66243_ (_20686_, _20685_, _20684_);
  and _66244_ (_20687_, _20686_, _18450_);
  nand _66245_ (_20688_, _18400_, _20127_);
  or _66246_ (_20689_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _66247_ (_20690_, _20689_, _20688_);
  and _66248_ (_20691_, _20690_, _18466_);
  or _66249_ (_20692_, _20691_, _20687_);
  nor _66250_ (_20693_, _20692_, _20683_);
  and _66251_ (_20694_, _20693_, _20679_);
  or _66252_ (_20695_, _20694_, _20674_);
  nor _66253_ (_20696_, _20695_, _18441_);
  or _66254_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _20696_, _20651_);
  and _66255_ (_20697_, _18441_, word_in[2]);
  not _66256_ (_20698_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand _66257_ (_20699_, _18400_, _20698_);
  or _66258_ (_20700_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _66259_ (_20701_, _20700_, _20699_);
  and _66260_ (_20702_, _20701_, _18447_);
  nor _66261_ (_20703_, _20702_, _18385_);
  not _66262_ (_20704_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand _66263_ (_20705_, _18400_, _20704_);
  or _66264_ (_20706_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _66265_ (_20707_, _20706_, _20705_);
  and _66266_ (_20708_, _20707_, _18456_);
  nand _66267_ (_20709_, _18400_, _19735_);
  or _66268_ (_20710_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _66269_ (_20711_, _20710_, _20709_);
  and _66270_ (_20712_, _20711_, _18450_);
  not _66271_ (_20713_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand _66272_ (_20714_, _18400_, _20713_);
  or _66273_ (_20715_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _66274_ (_20716_, _20715_, _20714_);
  and _66275_ (_20717_, _20716_, _18466_);
  or _66276_ (_20718_, _20717_, _20712_);
  nor _66277_ (_20719_, _20718_, _20708_);
  and _66278_ (_20720_, _20719_, _20703_);
  nand _66279_ (_20721_, _18400_, _19937_);
  or _66280_ (_20722_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _66281_ (_20723_, _20722_, _20721_);
  and _66282_ (_20724_, _20723_, _18447_);
  nor _66283_ (_20725_, _20724_, _18471_);
  nand _66284_ (_20726_, _18400_, _20547_);
  or _66285_ (_20727_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _66286_ (_20728_, _20727_, _20726_);
  and _66287_ (_20729_, _20728_, _18450_);
  nand _66288_ (_20730_, _18400_, _20346_);
  or _66289_ (_20731_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _66290_ (_20732_, _20731_, _20730_);
  and _66291_ (_20733_, _20732_, _18456_);
  or _66292_ (_20734_, _20733_, _20729_);
  nand _66293_ (_20735_, _18400_, _20142_);
  or _66294_ (_20736_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _66295_ (_20737_, _20736_, _20735_);
  and _66296_ (_20738_, _20737_, _18466_);
  nor _66297_ (_20739_, _20738_, _20734_);
  and _66298_ (_20740_, _20739_, _20725_);
  or _66299_ (_20741_, _20740_, _20720_);
  nor _66300_ (_20742_, _20741_, _18441_);
  or _66301_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _20742_, _20697_);
  and _66302_ (_20743_, _18441_, word_in[3]);
  not _66303_ (_20744_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nand _66304_ (_20745_, _18400_, _20744_);
  or _66305_ (_20746_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _66306_ (_20747_, _20746_, _20745_);
  and _66307_ (_20748_, _20747_, _18447_);
  nor _66308_ (_20749_, _20748_, _18385_);
  not _66309_ (_20750_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nand _66310_ (_20751_, _18400_, _20750_);
  or _66311_ (_20752_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _66312_ (_20753_, _20752_, _20751_);
  and _66313_ (_20754_, _20753_, _18456_);
  nand _66314_ (_20755_, _18400_, _19745_);
  or _66315_ (_20756_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _66316_ (_20757_, _20756_, _20755_);
  and _66317_ (_20758_, _20757_, _18450_);
  not _66318_ (_20759_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nand _66319_ (_20760_, _18400_, _20759_);
  or _66320_ (_20761_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _66321_ (_20762_, _20761_, _20760_);
  and _66322_ (_20763_, _20762_, _18466_);
  or _66323_ (_20764_, _20763_, _20758_);
  nor _66324_ (_20765_, _20764_, _20754_);
  and _66325_ (_20766_, _20765_, _20749_);
  nand _66326_ (_20767_, _18400_, _19951_);
  or _66327_ (_20768_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and _66328_ (_20769_, _20768_, _20767_);
  and _66329_ (_20770_, _20769_, _18447_);
  nor _66330_ (_20771_, _20770_, _18471_);
  nand _66331_ (_20772_, _18400_, _20359_);
  or _66332_ (_20773_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and _66333_ (_20774_, _20773_, _20772_);
  and _66334_ (_20775_, _20774_, _18456_);
  nand _66335_ (_20776_, _18400_, _20559_);
  or _66336_ (_20777_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _66337_ (_20778_, _20777_, _20776_);
  and _66338_ (_20779_, _20778_, _18450_);
  nand _66339_ (_20780_, _18400_, _20154_);
  or _66340_ (_20781_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _66341_ (_20782_, _20781_, _20780_);
  and _66342_ (_20783_, _20782_, _18466_);
  or _66343_ (_20784_, _20783_, _20779_);
  nor _66344_ (_20785_, _20784_, _20775_);
  and _66345_ (_20786_, _20785_, _20771_);
  or _66346_ (_20787_, _20786_, _20766_);
  nor _66347_ (_20788_, _20787_, _18441_);
  or _66348_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _20788_, _20743_);
  and _66349_ (_20789_, _18441_, word_in[4]);
  not _66350_ (_20790_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nand _66351_ (_20791_, _18400_, _20790_);
  or _66352_ (_20792_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _66353_ (_20793_, _20792_, _20791_);
  and _66354_ (_20794_, _20793_, _18447_);
  nor _66355_ (_20795_, _20794_, _18385_);
  not _66356_ (_20796_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nand _66357_ (_20797_, _18400_, _20796_);
  or _66358_ (_20798_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _66359_ (_20799_, _20798_, _20797_);
  and _66360_ (_20800_, _20799_, _18456_);
  nand _66361_ (_20801_, _18400_, _19759_);
  or _66362_ (_20802_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _66363_ (_20803_, _20802_, _20801_);
  and _66364_ (_20804_, _20803_, _18450_);
  not _66365_ (_20805_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nand _66366_ (_20806_, _18400_, _20805_);
  or _66367_ (_20807_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _66368_ (_20808_, _20807_, _20806_);
  and _66369_ (_20809_, _20808_, _18466_);
  or _66370_ (_20810_, _20809_, _20804_);
  nor _66371_ (_20811_, _20810_, _20800_);
  and _66372_ (_20812_, _20811_, _20795_);
  nand _66373_ (_20813_, _18400_, _19963_);
  or _66374_ (_20814_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and _66375_ (_20815_, _20814_, _20813_);
  and _66376_ (_20816_, _20815_, _18447_);
  nor _66377_ (_20817_, _20816_, _18471_);
  nand _66378_ (_20818_, _18400_, _20372_);
  or _66379_ (_20819_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and _66380_ (_20820_, _20819_, _20818_);
  and _66381_ (_20821_, _20820_, _18456_);
  nand _66382_ (_20822_, _18400_, _20571_);
  or _66383_ (_20823_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _66384_ (_20824_, _20823_, _20822_);
  and _66385_ (_20825_, _20824_, _18450_);
  nand _66386_ (_20826_, _18400_, _20165_);
  or _66387_ (_20827_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _66388_ (_20828_, _20827_, _20826_);
  and _66389_ (_20829_, _20828_, _18466_);
  or _66390_ (_20830_, _20829_, _20825_);
  nor _66391_ (_20831_, _20830_, _20821_);
  and _66392_ (_20832_, _20831_, _20817_);
  or _66393_ (_20833_, _20832_, _20812_);
  nor _66394_ (_20834_, _20833_, _18441_);
  or _66395_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _20834_, _20789_);
  and _66396_ (_20835_, _18441_, word_in[5]);
  not _66397_ (_20836_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nand _66398_ (_20837_, _18400_, _20836_);
  or _66399_ (_20838_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _66400_ (_20839_, _20838_, _20837_);
  and _66401_ (_20840_, _20839_, _18447_);
  nor _66402_ (_20841_, _20840_, _18385_);
  not _66403_ (_20842_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nand _66404_ (_20843_, _18400_, _20842_);
  or _66405_ (_20844_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _66406_ (_20845_, _20844_, _20843_);
  and _66407_ (_20846_, _20845_, _18456_);
  nand _66408_ (_20847_, _18400_, _19770_);
  or _66409_ (_20848_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _66410_ (_20849_, _20848_, _20847_);
  and _66411_ (_20850_, _20849_, _18450_);
  not _66412_ (_20851_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nand _66413_ (_20852_, _18400_, _20851_);
  or _66414_ (_20853_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _66415_ (_20854_, _20853_, _20852_);
  and _66416_ (_20855_, _20854_, _18466_);
  or _66417_ (_20856_, _20855_, _20850_);
  nor _66418_ (_20857_, _20856_, _20846_);
  and _66419_ (_20858_, _20857_, _20841_);
  nand _66420_ (_20859_, _18400_, _19975_);
  or _66421_ (_20860_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _66422_ (_20861_, _20860_, _20859_);
  and _66423_ (_20862_, _20861_, _18447_);
  nor _66424_ (_20863_, _20862_, _18471_);
  nand _66425_ (_20864_, _18400_, _20382_);
  or _66426_ (_20865_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _66427_ (_20866_, _20865_, _20864_);
  and _66428_ (_20867_, _20866_, _18456_);
  nand _66429_ (_20868_, _18400_, _20584_);
  or _66430_ (_20869_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _66431_ (_20870_, _20869_, _20868_);
  and _66432_ (_20871_, _20870_, _18450_);
  nand _66433_ (_20872_, _18400_, _20178_);
  or _66434_ (_20873_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _66435_ (_20874_, _20873_, _20872_);
  and _66436_ (_20875_, _20874_, _18466_);
  or _66437_ (_20876_, _20875_, _20871_);
  nor _66438_ (_20877_, _20876_, _20867_);
  and _66439_ (_20878_, _20877_, _20863_);
  or _66440_ (_20879_, _20878_, _20858_);
  nor _66441_ (_20880_, _20879_, _18441_);
  or _66442_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _20880_, _20835_);
  and _66443_ (_20881_, _18441_, word_in[6]);
  not _66444_ (_20882_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nand _66445_ (_20883_, _18400_, _20882_);
  or _66446_ (_20884_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _66447_ (_20885_, _20884_, _20883_);
  and _66448_ (_20886_, _20885_, _18447_);
  nor _66449_ (_20887_, _20886_, _18385_);
  not _66450_ (_20888_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nand _66451_ (_20889_, _18400_, _20888_);
  or _66452_ (_20890_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _66453_ (_20891_, _20890_, _20889_);
  and _66454_ (_20892_, _20891_, _18456_);
  nand _66455_ (_20893_, _18400_, _19782_);
  or _66456_ (_20894_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _66457_ (_20895_, _20894_, _20893_);
  and _66458_ (_20896_, _20895_, _18450_);
  not _66459_ (_20897_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nand _66460_ (_20898_, _18400_, _20897_);
  or _66461_ (_20899_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _66462_ (_20900_, _20899_, _20898_);
  and _66463_ (_20901_, _20900_, _18466_);
  or _66464_ (_20902_, _20901_, _20896_);
  nor _66465_ (_20903_, _20902_, _20892_);
  and _66466_ (_20904_, _20903_, _20887_);
  nand _66467_ (_20905_, _18400_, _19988_);
  or _66468_ (_20906_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _66469_ (_20907_, _20906_, _20905_);
  and _66470_ (_20908_, _20907_, _18447_);
  nor _66471_ (_20909_, _20908_, _18471_);
  nand _66472_ (_20910_, _18400_, _20593_);
  or _66473_ (_20911_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _66474_ (_20912_, _20911_, _20910_);
  and _66475_ (_20913_, _20912_, _18450_);
  nand _66476_ (_20914_, _18400_, _20395_);
  or _66477_ (_20915_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _66478_ (_20916_, _20915_, _20914_);
  and _66479_ (_20917_, _20916_, _18456_);
  or _66480_ (_20918_, _20917_, _20913_);
  nand _66481_ (_20919_, _18400_, _20190_);
  or _66482_ (_20920_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _66483_ (_20921_, _20920_, _20919_);
  and _66484_ (_20922_, _20921_, _18466_);
  nor _66485_ (_20923_, _20922_, _20918_);
  and _66486_ (_20924_, _20923_, _20909_);
  or _66487_ (_20925_, _20924_, _20904_);
  nor _66488_ (_20926_, _20925_, _18441_);
  or _66489_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _20926_, _20881_);
  and _66490_ (_20927_, _18553_, word_in[8]);
  nand _66491_ (_20928_, _18400_, _18987_);
  or _66492_ (_20929_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _66493_ (_20930_, _20929_, _20928_);
  and _66494_ (_20931_, _20930_, _18555_);
  and _66495_ (_20932_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor _66496_ (_20933_, _18400_, _20621_);
  or _66497_ (_20934_, _20933_, _20932_);
  and _66498_ (_20935_, _20934_, _18561_);
  nor _66499_ (_20936_, _20935_, _20931_);
  nor _66500_ (_20937_, _20936_, _18500_);
  and _66501_ (_20938_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _66502_ (_20939_, _18400_, _20612_);
  or _66503_ (_20940_, _20939_, _20938_);
  and _66504_ (_20941_, _20940_, _18555_);
  nand _66505_ (_20942_, _18400_, _19604_);
  or _66506_ (_20943_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _66507_ (_20944_, _20943_, _20942_);
  and _66508_ (_20945_, _20944_, _18561_);
  or _66509_ (_20946_, _20945_, _20941_);
  and _66510_ (_20947_, _20946_, _18500_);
  or _66511_ (_20948_, _20947_, _20937_);
  and _66512_ (_20949_, _20948_, _18504_);
  nand _66513_ (_20950_, _18400_, _19807_);
  or _66514_ (_20951_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _66515_ (_20952_, _20951_, _20950_);
  and _66516_ (_20953_, _20952_, _18555_);
  nand _66517_ (_20954_, _18400_, _20016_);
  or _66518_ (_20955_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _66519_ (_20956_, _20955_, _20954_);
  and _66520_ (_20957_, _20956_, _18561_);
  nor _66521_ (_20958_, _20957_, _20953_);
  nor _66522_ (_20959_, _20958_, _18500_);
  nand _66523_ (_20960_, _18400_, _20218_);
  or _66524_ (_20961_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _66525_ (_20962_, _20961_, _20960_);
  and _66526_ (_20963_, _20962_, _18555_);
  nand _66527_ (_20964_, _18400_, _20420_);
  or _66528_ (_20965_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _66529_ (_20966_, _20965_, _20964_);
  and _66530_ (_20967_, _20966_, _18561_);
  or _66531_ (_20968_, _20967_, _20963_);
  and _66532_ (_20969_, _20968_, _18500_);
  nor _66533_ (_20970_, _20969_, _20959_);
  nor _66534_ (_20971_, _20970_, _18504_);
  nor _66535_ (_20972_, _20971_, _20949_);
  nor _66536_ (_20973_, _20972_, _18553_);
  or _66537_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _20973_, _20927_);
  and _66538_ (_20974_, _18553_, word_in[9]);
  nand _66539_ (_20975_, _18400_, _19003_);
  or _66540_ (_20976_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _66541_ (_20977_, _20976_, _20975_);
  and _66542_ (_20978_, _20977_, _18555_);
  and _66543_ (_20979_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _66544_ (_20980_, _18400_, _20667_);
  or _66545_ (_20981_, _20980_, _20979_);
  and _66546_ (_20982_, _20981_, _18561_);
  nor _66547_ (_20983_, _20982_, _20978_);
  nor _66548_ (_20984_, _20983_, _18500_);
  and _66549_ (_20985_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _66550_ (_20986_, _18400_, _20658_);
  or _66551_ (_20987_, _20986_, _20985_);
  and _66552_ (_20988_, _20987_, _18555_);
  nand _66553_ (_20989_, _18400_, _19618_);
  or _66554_ (_20990_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _66555_ (_20991_, _20990_, _20989_);
  and _66556_ (_20992_, _20991_, _18561_);
  or _66557_ (_20993_, _20992_, _20988_);
  and _66558_ (_20994_, _20993_, _18500_);
  or _66559_ (_20995_, _20994_, _20984_);
  and _66560_ (_20996_, _20995_, _18504_);
  nand _66561_ (_20997_, _18400_, _19825_);
  or _66562_ (_20998_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _66563_ (_20999_, _20998_, _20997_);
  and _66564_ (_21000_, _20999_, _18555_);
  nand _66565_ (_21001_, _18400_, _20028_);
  or _66566_ (_21002_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _66567_ (_21003_, _21002_, _21001_);
  and _66568_ (_21004_, _21003_, _18561_);
  nor _66569_ (_21005_, _21004_, _21000_);
  nor _66570_ (_21006_, _21005_, _18500_);
  nand _66571_ (_21007_, _18400_, _20232_);
  or _66572_ (_21008_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _66573_ (_21009_, _21008_, _21007_);
  and _66574_ (_21010_, _21009_, _18555_);
  nand _66575_ (_21011_, _18400_, _20438_);
  or _66576_ (_21012_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _66577_ (_21013_, _21012_, _21011_);
  and _66578_ (_21014_, _21013_, _18561_);
  or _66579_ (_21015_, _21014_, _21010_);
  and _66580_ (_21016_, _21015_, _18500_);
  nor _66581_ (_21017_, _21016_, _21006_);
  nor _66582_ (_21018_, _21017_, _18504_);
  nor _66583_ (_21019_, _21018_, _20996_);
  nor _66584_ (_21020_, _21019_, _18553_);
  or _66585_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _21020_, _20974_);
  and _66586_ (_21021_, _18553_, word_in[10]);
  nand _66587_ (_21022_, _18400_, _19016_);
  or _66588_ (_21023_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _66589_ (_21024_, _21023_, _21022_);
  and _66590_ (_21025_, _21024_, _18555_);
  and _66591_ (_21026_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _66592_ (_21027_, _18400_, _20713_);
  or _66593_ (_21028_, _21027_, _21026_);
  and _66594_ (_21029_, _21028_, _18561_);
  nor _66595_ (_21030_, _21029_, _21025_);
  nor _66596_ (_21031_, _21030_, _18500_);
  and _66597_ (_21032_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _66598_ (_21033_, _18400_, _20704_);
  or _66599_ (_21034_, _21033_, _21032_);
  and _66600_ (_21035_, _21034_, _18555_);
  nand _66601_ (_21036_, _18400_, _19632_);
  or _66602_ (_21037_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _66603_ (_21038_, _21037_, _21036_);
  and _66604_ (_21039_, _21038_, _18561_);
  or _66605_ (_21040_, _21039_, _21035_);
  and _66606_ (_21041_, _21040_, _18500_);
  or _66607_ (_21042_, _21041_, _21031_);
  and _66608_ (_21043_, _21042_, _18504_);
  nand _66609_ (_21044_, _18400_, _19837_);
  or _66610_ (_21045_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _66611_ (_21046_, _21045_, _21044_);
  and _66612_ (_21047_, _21046_, _18555_);
  nand _66613_ (_21048_, _18400_, _20040_);
  or _66614_ (_21049_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _66615_ (_21050_, _21049_, _21048_);
  and _66616_ (_21051_, _21050_, _18561_);
  nor _66617_ (_21052_, _21051_, _21047_);
  nor _66618_ (_21053_, _21052_, _18500_);
  nand _66619_ (_21054_, _18400_, _20245_);
  or _66620_ (_21055_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and _66621_ (_21056_, _21055_, _21054_);
  and _66622_ (_21057_, _21056_, _18555_);
  nand _66623_ (_21058_, _18400_, _20450_);
  or _66624_ (_21059_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _66625_ (_21060_, _21059_, _21058_);
  and _66626_ (_21061_, _21060_, _18561_);
  or _66627_ (_21062_, _21061_, _21057_);
  and _66628_ (_21063_, _21062_, _18500_);
  nor _66629_ (_21064_, _21063_, _21053_);
  nor _66630_ (_21065_, _21064_, _18504_);
  nor _66631_ (_21066_, _21065_, _21043_);
  nor _66632_ (_21067_, _21066_, _18553_);
  or _66633_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _21067_, _21021_);
  and _66634_ (_21068_, _18553_, word_in[11]);
  nand _66635_ (_21069_, _18400_, _19027_);
  or _66636_ (_21070_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and _66637_ (_21071_, _21070_, _21069_);
  and _66638_ (_21072_, _21071_, _18555_);
  and _66639_ (_21073_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor _66640_ (_21074_, _18400_, _20759_);
  or _66641_ (_21075_, _21074_, _21073_);
  and _66642_ (_21076_, _21075_, _18561_);
  nor _66643_ (_21077_, _21076_, _21072_);
  nor _66644_ (_21078_, _21077_, _18500_);
  and _66645_ (_21079_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _66646_ (_21080_, _18400_, _20750_);
  or _66647_ (_21081_, _21080_, _21079_);
  and _66648_ (_21082_, _21081_, _18555_);
  nand _66649_ (_21083_, _18400_, _19645_);
  or _66650_ (_21084_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _66651_ (_21085_, _21084_, _21083_);
  and _66652_ (_21086_, _21085_, _18561_);
  or _66653_ (_21087_, _21086_, _21082_);
  and _66654_ (_21088_, _21087_, _18500_);
  or _66655_ (_21089_, _21088_, _21078_);
  and _66656_ (_21090_, _21089_, _18504_);
  nand _66657_ (_21091_, _18400_, _19849_);
  or _66658_ (_21092_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _66659_ (_21093_, _21092_, _21091_);
  and _66660_ (_21094_, _21093_, _18555_);
  nand _66661_ (_21095_, _18400_, _20052_);
  or _66662_ (_21096_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _66663_ (_21097_, _21096_, _21095_);
  and _66664_ (_21098_, _21097_, _18561_);
  nor _66665_ (_21099_, _21098_, _21094_);
  nor _66666_ (_21100_, _21099_, _18500_);
  nand _66667_ (_21101_, _18400_, _20257_);
  or _66668_ (_21102_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _66669_ (_21103_, _21102_, _21101_);
  and _66670_ (_21104_, _21103_, _18555_);
  nand _66671_ (_21105_, _18400_, _20461_);
  or _66672_ (_21106_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _66673_ (_21107_, _21106_, _21105_);
  and _66674_ (_21108_, _21107_, _18561_);
  or _66675_ (_21109_, _21108_, _21104_);
  and _66676_ (_21110_, _21109_, _18500_);
  nor _66677_ (_21111_, _21110_, _21100_);
  nor _66678_ (_21112_, _21111_, _18504_);
  nor _66679_ (_21113_, _21112_, _21090_);
  nor _66680_ (_21114_, _21113_, _18553_);
  or _66681_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _21114_, _21068_);
  and _66682_ (_21115_, _18553_, word_in[12]);
  nand _66683_ (_21116_, _18400_, _19042_);
  or _66684_ (_21117_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _66685_ (_21118_, _21117_, _21116_);
  and _66686_ (_21119_, _21118_, _18555_);
  and _66687_ (_21120_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _66688_ (_21121_, _18400_, _20805_);
  or _66689_ (_21122_, _21121_, _21120_);
  and _66690_ (_21123_, _21122_, _18561_);
  nor _66691_ (_21124_, _21123_, _21119_);
  nor _66692_ (_21125_, _21124_, _18500_);
  and _66693_ (_21126_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _66694_ (_21127_, _18400_, _20796_);
  or _66695_ (_21128_, _21127_, _21126_);
  and _66696_ (_21129_, _21128_, _18555_);
  nand _66697_ (_21130_, _18400_, _19657_);
  or _66698_ (_21131_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _66699_ (_21132_, _21131_, _21130_);
  and _66700_ (_21133_, _21132_, _18561_);
  or _66701_ (_21134_, _21133_, _21129_);
  and _66702_ (_21135_, _21134_, _18500_);
  or _66703_ (_21136_, _21135_, _21125_);
  and _66704_ (_21137_, _21136_, _18504_);
  nand _66705_ (_21138_, _18400_, _19860_);
  or _66706_ (_21139_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _66707_ (_21140_, _21139_, _21138_);
  and _66708_ (_21141_, _21140_, _18555_);
  nand _66709_ (_21142_, _18400_, _20064_);
  or _66710_ (_21143_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _66711_ (_21144_, _21143_, _21142_);
  and _66712_ (_21145_, _21144_, _18561_);
  nor _66713_ (_21146_, _21145_, _21141_);
  nor _66714_ (_21147_, _21146_, _18500_);
  nand _66715_ (_21148_, _18400_, _20269_);
  or _66716_ (_21149_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and _66717_ (_21150_, _21149_, _21148_);
  and _66718_ (_21151_, _21150_, _18555_);
  nand _66719_ (_21152_, _18400_, _20473_);
  or _66720_ (_21153_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _66721_ (_21154_, _21153_, _21152_);
  and _66722_ (_21155_, _21154_, _18561_);
  or _66723_ (_21156_, _21155_, _21151_);
  and _66724_ (_21157_, _21156_, _18500_);
  nor _66725_ (_21158_, _21157_, _21147_);
  nor _66726_ (_21159_, _21158_, _18504_);
  nor _66727_ (_21160_, _21159_, _21137_);
  nor _66728_ (_21161_, _21160_, _18553_);
  or _66729_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _21161_, _21115_);
  and _66730_ (_21162_, _18553_, word_in[13]);
  nand _66731_ (_21163_, _18400_, _19054_);
  or _66732_ (_21164_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _66733_ (_21165_, _21164_, _21163_);
  and _66734_ (_21166_, _21165_, _18555_);
  and _66735_ (_21167_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _66736_ (_21168_, _18400_, _20851_);
  or _66737_ (_21169_, _21168_, _21167_);
  and _66738_ (_21170_, _21169_, _18561_);
  nor _66739_ (_21171_, _21170_, _21166_);
  nor _66740_ (_21172_, _21171_, _18500_);
  and _66741_ (_21173_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _66742_ (_21174_, _18400_, _20842_);
  or _66743_ (_21175_, _21174_, _21173_);
  and _66744_ (_21176_, _21175_, _18555_);
  nand _66745_ (_21177_, _18400_, _19667_);
  or _66746_ (_21178_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _66747_ (_21179_, _21178_, _21177_);
  and _66748_ (_21180_, _21179_, _18561_);
  or _66749_ (_21181_, _21180_, _21176_);
  and _66750_ (_21182_, _21181_, _18500_);
  or _66751_ (_21183_, _21182_, _21172_);
  and _66752_ (_21184_, _21183_, _18504_);
  nand _66753_ (_21185_, _18400_, _19873_);
  or _66754_ (_21186_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _66755_ (_21187_, _21186_, _21185_);
  and _66756_ (_21188_, _21187_, _18555_);
  nand _66757_ (_21189_, _18400_, _20076_);
  or _66758_ (_21190_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _66759_ (_21191_, _21190_, _21189_);
  and _66760_ (_21192_, _21191_, _18561_);
  nor _66761_ (_21193_, _21192_, _21188_);
  nor _66762_ (_21194_, _21193_, _18500_);
  nand _66763_ (_21195_, _18400_, _20281_);
  or _66764_ (_21196_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _66765_ (_21197_, _21196_, _21195_);
  and _66766_ (_21198_, _21197_, _18555_);
  nand _66767_ (_21199_, _18400_, _20486_);
  or _66768_ (_21200_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _66769_ (_21201_, _21200_, _21199_);
  and _66770_ (_21202_, _21201_, _18561_);
  or _66771_ (_21203_, _21202_, _21198_);
  and _66772_ (_21204_, _21203_, _18500_);
  nor _66773_ (_21205_, _21204_, _21194_);
  nor _66774_ (_21206_, _21205_, _18504_);
  nor _66775_ (_21207_, _21206_, _21184_);
  nor _66776_ (_21208_, _21207_, _18553_);
  or _66777_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _21208_, _21162_);
  and _66778_ (_21209_, _18553_, word_in[14]);
  nand _66779_ (_21210_, _18400_, _19065_);
  or _66780_ (_21211_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _66781_ (_21212_, _21211_, _21210_);
  and _66782_ (_21213_, _21212_, _18555_);
  and _66783_ (_21214_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _66784_ (_21215_, _18400_, _20897_);
  or _66785_ (_21216_, _21215_, _21214_);
  and _66786_ (_21217_, _21216_, _18561_);
  nor _66787_ (_21218_, _21217_, _21213_);
  nor _66788_ (_21219_, _21218_, _18500_);
  and _66789_ (_21220_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _66790_ (_21221_, _18400_, _20888_);
  or _66791_ (_21222_, _21221_, _21220_);
  and _66792_ (_21223_, _21222_, _18555_);
  nand _66793_ (_21224_, _18400_, _19679_);
  or _66794_ (_21225_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _66795_ (_21226_, _21225_, _21224_);
  and _66796_ (_21227_, _21226_, _18561_);
  or _66797_ (_21228_, _21227_, _21223_);
  and _66798_ (_21229_, _21228_, _18500_);
  or _66799_ (_21230_, _21229_, _21219_);
  and _66800_ (_21231_, _21230_, _18504_);
  nand _66801_ (_21232_, _18400_, _19885_);
  or _66802_ (_21233_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _66803_ (_21234_, _21233_, _21232_);
  and _66804_ (_21235_, _21234_, _18555_);
  nand _66805_ (_21236_, _18400_, _20087_);
  or _66806_ (_21237_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _66807_ (_21238_, _21237_, _21236_);
  and _66808_ (_21239_, _21238_, _18561_);
  nor _66809_ (_21240_, _21239_, _21235_);
  nor _66810_ (_21241_, _21240_, _18500_);
  nand _66811_ (_21242_, _18400_, _20292_);
  or _66812_ (_21243_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _66813_ (_21244_, _21243_, _21242_);
  and _66814_ (_21245_, _21244_, _18555_);
  nand _66815_ (_21246_, _18400_, _20498_);
  or _66816_ (_21247_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _66817_ (_21248_, _21247_, _21246_);
  and _66818_ (_21249_, _21248_, _18561_);
  or _66819_ (_21250_, _21249_, _21245_);
  and _66820_ (_21251_, _21250_, _18500_);
  nor _66821_ (_21252_, _21251_, _21241_);
  nor _66822_ (_21253_, _21252_, _18504_);
  nor _66823_ (_21254_, _21253_, _21231_);
  nor _66824_ (_21255_, _21254_, _18553_);
  or _66825_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _21255_, _21209_);
  and _66826_ (_21256_, _18672_, word_in[16]);
  and _66827_ (_21257_, _20636_, _18466_);
  and _66828_ (_21258_, _20640_, _18456_);
  or _66829_ (_21259_, _21258_, _21257_);
  and _66830_ (_21260_, _20631_, _18450_);
  and _66831_ (_21261_, _20644_, _18447_);
  or _66832_ (_21262_, _21261_, _21260_);
  or _66833_ (_21263_, _21262_, _21259_);
  or _66834_ (_21264_, _21263_, _18613_);
  and _66835_ (_21265_, _20615_, _18466_);
  and _66836_ (_21266_, _20619_, _18456_);
  or _66837_ (_21267_, _21266_, _21265_);
  and _66838_ (_21268_, _20609_, _18450_);
  and _66839_ (_21269_, _20624_, _18447_);
  or _66840_ (_21270_, _21269_, _21268_);
  nor _66841_ (_21271_, _21270_, _21267_);
  nand _66842_ (_21272_, _21271_, _18613_);
  and _66843_ (_21273_, _21272_, _21264_);
  and _66844_ (_21274_, _21273_, _18671_);
  or _66845_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _21274_, _21256_);
  and _66846_ (_21275_, _18672_, word_in[17]);
  and _66847_ (_21276_, _20686_, _18456_);
  and _66848_ (_21277_, _20682_, _18466_);
  or _66849_ (_21278_, _21277_, _21276_);
  and _66850_ (_21279_, _20690_, _18447_);
  and _66851_ (_21280_, _20677_, _18450_);
  or _66852_ (_21281_, _21280_, _21279_);
  or _66853_ (_21282_, _21281_, _21278_);
  or _66854_ (_21283_, _21282_, _18613_);
  and _66855_ (_21284_, _20665_, _18456_);
  and _66856_ (_21285_, _20661_, _18466_);
  or _66857_ (_21286_, _21285_, _21284_);
  and _66858_ (_21287_, _20670_, _18447_);
  and _66859_ (_21288_, _20655_, _18450_);
  or _66860_ (_21289_, _21288_, _21287_);
  nor _66861_ (_21290_, _21289_, _21286_);
  nand _66862_ (_21291_, _21290_, _18613_);
  and _66863_ (_21292_, _21291_, _21283_);
  and _66864_ (_21293_, _21292_, _18671_);
  or _66865_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _21293_, _21275_);
  and _66866_ (_21294_, _18672_, word_in[18]);
  and _66867_ (_21295_, _20732_, _18466_);
  and _66868_ (_21296_, _20728_, _18456_);
  or _66869_ (_21297_, _21296_, _21295_);
  and _66870_ (_21298_, _20723_, _18450_);
  and _66871_ (_21299_, _20737_, _18447_);
  or _66872_ (_21300_, _21299_, _21298_);
  or _66873_ (_21301_, _21300_, _21297_);
  or _66874_ (_21302_, _21301_, _18613_);
  and _66875_ (_21303_, _20707_, _18466_);
  and _66876_ (_21304_, _20711_, _18456_);
  or _66877_ (_21305_, _21304_, _21303_);
  and _66878_ (_21306_, _20701_, _18450_);
  and _66879_ (_21307_, _20716_, _18447_);
  or _66880_ (_21308_, _21307_, _21306_);
  nor _66881_ (_21309_, _21308_, _21305_);
  nand _66882_ (_21310_, _21309_, _18613_);
  and _66883_ (_21311_, _21310_, _21302_);
  and _66884_ (_21312_, _21311_, _18671_);
  or _66885_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _21312_, _21294_);
  and _66886_ (_21313_, _18672_, word_in[19]);
  and _66887_ (_21314_, _20774_, _18466_);
  and _66888_ (_21315_, _20778_, _18456_);
  or _66889_ (_21316_, _21315_, _21314_);
  and _66890_ (_21317_, _20769_, _18450_);
  and _66891_ (_21318_, _20782_, _18447_);
  or _66892_ (_21319_, _21318_, _21317_);
  or _66893_ (_21320_, _21319_, _21316_);
  or _66894_ (_21321_, _21320_, _18613_);
  and _66895_ (_21322_, _20757_, _18456_);
  and _66896_ (_21323_, _20753_, _18466_);
  or _66897_ (_21324_, _21323_, _21322_);
  and _66898_ (_21325_, _20762_, _18447_);
  and _66899_ (_21326_, _20747_, _18450_);
  or _66900_ (_21327_, _21326_, _21325_);
  nor _66901_ (_21328_, _21327_, _21324_);
  nand _66902_ (_21329_, _21328_, _18613_);
  and _66903_ (_21330_, _21329_, _21321_);
  and _66904_ (_21331_, _21330_, _18671_);
  or _66905_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _21331_, _21313_);
  and _66906_ (_21332_, _18672_, word_in[20]);
  and _66907_ (_21333_, _20824_, _18456_);
  and _66908_ (_21334_, _20820_, _18466_);
  or _66909_ (_21335_, _21334_, _21333_);
  and _66910_ (_21336_, _20828_, _18447_);
  and _66911_ (_21337_, _20815_, _18450_);
  or _66912_ (_21338_, _21337_, _21336_);
  or _66913_ (_21339_, _21338_, _21335_);
  or _66914_ (_21340_, _21339_, _18613_);
  and _66915_ (_21341_, _20799_, _18466_);
  and _66916_ (_21342_, _20803_, _18456_);
  or _66917_ (_21343_, _21342_, _21341_);
  and _66918_ (_21344_, _20793_, _18450_);
  and _66919_ (_21345_, _20808_, _18447_);
  or _66920_ (_21346_, _21345_, _21344_);
  nor _66921_ (_21347_, _21346_, _21343_);
  nand _66922_ (_21348_, _21347_, _18613_);
  and _66923_ (_21349_, _21348_, _21340_);
  and _66924_ (_21350_, _21349_, _18671_);
  or _66925_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _21350_, _21332_);
  and _66926_ (_21351_, _18672_, word_in[21]);
  and _66927_ (_21352_, _20866_, _18466_);
  and _66928_ (_21353_, _20870_, _18456_);
  or _66929_ (_21354_, _21353_, _21352_);
  and _66930_ (_21355_, _20861_, _18450_);
  and _66931_ (_21356_, _20874_, _18447_);
  or _66932_ (_21357_, _21356_, _21355_);
  or _66933_ (_21358_, _21357_, _21354_);
  or _66934_ (_21359_, _21358_, _18613_);
  and _66935_ (_21360_, _20845_, _18466_);
  and _66936_ (_21361_, _20849_, _18456_);
  or _66937_ (_21362_, _21361_, _21360_);
  and _66938_ (_21363_, _20839_, _18450_);
  and _66939_ (_21364_, _20854_, _18447_);
  or _66940_ (_21365_, _21364_, _21363_);
  nor _66941_ (_21366_, _21365_, _21362_);
  nand _66942_ (_21367_, _21366_, _18613_);
  and _66943_ (_21368_, _21367_, _21359_);
  and _66944_ (_21369_, _21368_, _18671_);
  or _66945_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _21369_, _21351_);
  and _66946_ (_21370_, _18672_, word_in[22]);
  and _66947_ (_21371_, _20916_, _18466_);
  and _66948_ (_21372_, _20912_, _18456_);
  or _66949_ (_21373_, _21372_, _21371_);
  and _66950_ (_21374_, _20907_, _18450_);
  and _66951_ (_21375_, _20921_, _18447_);
  or _66952_ (_21376_, _21375_, _21374_);
  or _66953_ (_21377_, _21376_, _21373_);
  or _66954_ (_21378_, _21377_, _18613_);
  and _66955_ (_21379_, _20895_, _18456_);
  and _66956_ (_21380_, _20891_, _18466_);
  or _66957_ (_21381_, _21380_, _21379_);
  and _66958_ (_21382_, _20900_, _18447_);
  and _66959_ (_21383_, _20885_, _18450_);
  or _66960_ (_21384_, _21383_, _21382_);
  nor _66961_ (_21385_, _21384_, _21381_);
  nand _66962_ (_21386_, _21385_, _18613_);
  and _66963_ (_21387_, _21386_, _21378_);
  and _66964_ (_21388_, _21387_, _18671_);
  or _66965_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _21388_, _21370_);
  and _66966_ (_21389_, _18741_, word_in[24]);
  and _66967_ (_21390_, _20966_, _18555_);
  and _66968_ (_21391_, _20962_, _18561_);
  or _66969_ (_21392_, _21391_, _21390_);
  and _66970_ (_21393_, _21392_, _18699_);
  and _66971_ (_21394_, _20956_, _18555_);
  and _66972_ (_21395_, _20952_, _18561_);
  nor _66973_ (_21396_, _21395_, _21394_);
  nor _66974_ (_21397_, _21396_, _18699_);
  or _66975_ (_21398_, _21397_, _21393_);
  and _66976_ (_21399_, _21398_, _18695_);
  and _66977_ (_21400_, _20944_, _18555_);
  and _66978_ (_21401_, _20940_, _18561_);
  or _66979_ (_21402_, _21401_, _21400_);
  and _66980_ (_21403_, _21402_, _18699_);
  and _66981_ (_21404_, _20930_, _18561_);
  and _66982_ (_21405_, _20934_, _18555_);
  nor _66983_ (_21406_, _21405_, _21404_);
  nor _66984_ (_21407_, _21406_, _18699_);
  or _66985_ (_21408_, _21407_, _21403_);
  and _66986_ (_21409_, _21408_, _18752_);
  nor _66987_ (_21410_, _21409_, _21399_);
  nor _66988_ (_21411_, _21410_, _18741_);
  or _66989_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _21411_, _21389_);
  and _66990_ (_21412_, _18741_, word_in[25]);
  and _66991_ (_21413_, _21013_, _18555_);
  and _66992_ (_21414_, _21009_, _18561_);
  or _66993_ (_21415_, _21414_, _21413_);
  and _66994_ (_21416_, _21415_, _18699_);
  and _66995_ (_21417_, _20999_, _18561_);
  and _66996_ (_21418_, _21003_, _18555_);
  nor _66997_ (_21419_, _21418_, _21417_);
  nor _66998_ (_21420_, _21419_, _18699_);
  or _66999_ (_21421_, _21420_, _21416_);
  and _67000_ (_21422_, _21421_, _18695_);
  and _67001_ (_21423_, _20991_, _18555_);
  and _67002_ (_21424_, _20987_, _18561_);
  or _67003_ (_21425_, _21424_, _21423_);
  and _67004_ (_21426_, _21425_, _18699_);
  and _67005_ (_21427_, _20977_, _18561_);
  and _67006_ (_21428_, _20981_, _18555_);
  nor _67007_ (_21429_, _21428_, _21427_);
  nor _67008_ (_21430_, _21429_, _18699_);
  or _67009_ (_21431_, _21430_, _21426_);
  and _67010_ (_21432_, _21431_, _18752_);
  nor _67011_ (_21433_, _21432_, _21422_);
  nor _67012_ (_21434_, _21433_, _18741_);
  or _67013_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _21434_, _21412_);
  and _67014_ (_21435_, _18741_, word_in[26]);
  and _67015_ (_21436_, _21060_, _18555_);
  and _67016_ (_21437_, _21056_, _18561_);
  or _67017_ (_21438_, _21437_, _21436_);
  and _67018_ (_21439_, _21438_, _18699_);
  and _67019_ (_21440_, _21046_, _18561_);
  and _67020_ (_21441_, _21050_, _18555_);
  nor _67021_ (_21442_, _21441_, _21440_);
  nor _67022_ (_21443_, _21442_, _18699_);
  or _67023_ (_21444_, _21443_, _21439_);
  and _67024_ (_21445_, _21444_, _18695_);
  and _67025_ (_21446_, _21038_, _18555_);
  and _67026_ (_21447_, _21034_, _18561_);
  or _67027_ (_21448_, _21447_, _21446_);
  and _67028_ (_21449_, _21448_, _18699_);
  and _67029_ (_21450_, _21024_, _18561_);
  and _67030_ (_21451_, _21028_, _18555_);
  nor _67031_ (_21452_, _21451_, _21450_);
  nor _67032_ (_21453_, _21452_, _18699_);
  or _67033_ (_21454_, _21453_, _21449_);
  and _67034_ (_21455_, _21454_, _18752_);
  nor _67035_ (_21456_, _21455_, _21445_);
  nor _67036_ (_21457_, _21456_, _18741_);
  or _67037_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _21457_, _21435_);
  and _67038_ (_21458_, _18741_, word_in[27]);
  and _67039_ (_21459_, _21107_, _18555_);
  and _67040_ (_21460_, _21103_, _18561_);
  or _67041_ (_21461_, _21460_, _21459_);
  and _67042_ (_21462_, _21461_, _18699_);
  and _67043_ (_21463_, _21093_, _18561_);
  and _67044_ (_21464_, _21097_, _18555_);
  nor _67045_ (_21465_, _21464_, _21463_);
  nor _67046_ (_21466_, _21465_, _18699_);
  or _67047_ (_21467_, _21466_, _21462_);
  and _67048_ (_21468_, _21467_, _18695_);
  and _67049_ (_21469_, _21075_, _18555_);
  and _67050_ (_21470_, _21071_, _18561_);
  nor _67051_ (_21471_, _21470_, _21469_);
  nor _67052_ (_21472_, _21471_, _18699_);
  and _67053_ (_21473_, _21085_, _18555_);
  and _67054_ (_21474_, _21081_, _18561_);
  or _67055_ (_21475_, _21474_, _21473_);
  and _67056_ (_21476_, _21475_, _18699_);
  or _67057_ (_21477_, _21476_, _21472_);
  and _67058_ (_21478_, _21477_, _18752_);
  nor _67059_ (_21479_, _21478_, _21468_);
  nor _67060_ (_21480_, _21479_, _18741_);
  or _67061_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _21480_, _21458_);
  and _67062_ (_21481_, _18741_, word_in[28]);
  and _67063_ (_21482_, _21154_, _18555_);
  and _67064_ (_21483_, _21150_, _18561_);
  or _67065_ (_21484_, _21483_, _21482_);
  and _67066_ (_21485_, _21484_, _18699_);
  and _67067_ (_21486_, _21140_, _18561_);
  and _67068_ (_21487_, _21144_, _18555_);
  nor _67069_ (_21488_, _21487_, _21486_);
  nor _67070_ (_21489_, _21488_, _18699_);
  or _67071_ (_21490_, _21489_, _21485_);
  and _67072_ (_21491_, _21490_, _18695_);
  and _67073_ (_21492_, _21132_, _18555_);
  and _67074_ (_21493_, _21128_, _18561_);
  or _67075_ (_21494_, _21493_, _21492_);
  and _67076_ (_21495_, _21494_, _18699_);
  and _67077_ (_21496_, _21118_, _18561_);
  and _67078_ (_21497_, _21122_, _18555_);
  nor _67079_ (_21498_, _21497_, _21496_);
  nor _67080_ (_21499_, _21498_, _18699_);
  or _67081_ (_21500_, _21499_, _21495_);
  and _67082_ (_21501_, _21500_, _18752_);
  nor _67083_ (_21502_, _21501_, _21491_);
  nor _67084_ (_21503_, _21502_, _18741_);
  or _67085_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _21503_, _21481_);
  and _67086_ (_21504_, _18741_, word_in[29]);
  and _67087_ (_21505_, _21201_, _18555_);
  and _67088_ (_21506_, _21197_, _18561_);
  or _67089_ (_21507_, _21506_, _21505_);
  and _67090_ (_21508_, _21507_, _18699_);
  and _67091_ (_21509_, _21187_, _18561_);
  and _67092_ (_21510_, _21191_, _18555_);
  nor _67093_ (_21511_, _21510_, _21509_);
  nor _67094_ (_21512_, _21511_, _18699_);
  or _67095_ (_21513_, _21512_, _21508_);
  and _67096_ (_21514_, _21513_, _18695_);
  and _67097_ (_21515_, _21179_, _18555_);
  and _67098_ (_21516_, _21175_, _18561_);
  or _67099_ (_21517_, _21516_, _21515_);
  and _67100_ (_21518_, _21517_, _18699_);
  and _67101_ (_21519_, _21165_, _18561_);
  and _67102_ (_21520_, _21169_, _18555_);
  nor _67103_ (_21521_, _21520_, _21519_);
  nor _67104_ (_21522_, _21521_, _18699_);
  or _67105_ (_21523_, _21522_, _21518_);
  and _67106_ (_21524_, _21523_, _18752_);
  nor _67107_ (_21525_, _21524_, _21514_);
  nor _67108_ (_21526_, _21525_, _18741_);
  or _67109_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _21526_, _21504_);
  and _67110_ (_21527_, _18741_, word_in[30]);
  and _67111_ (_21528_, _21248_, _18555_);
  and _67112_ (_21529_, _21244_, _18561_);
  or _67113_ (_21530_, _21529_, _21528_);
  and _67114_ (_21531_, _21530_, _18699_);
  and _67115_ (_21532_, _21238_, _18555_);
  and _67116_ (_21533_, _21234_, _18561_);
  nor _67117_ (_21534_, _21533_, _21532_);
  nor _67118_ (_21535_, _21534_, _18699_);
  or _67119_ (_21536_, _21535_, _21531_);
  and _67120_ (_21537_, _21536_, _18695_);
  and _67121_ (_21538_, _21226_, _18555_);
  and _67122_ (_21539_, _21222_, _18561_);
  or _67123_ (_21540_, _21539_, _21538_);
  and _67124_ (_21541_, _21540_, _18699_);
  and _67125_ (_21542_, _21212_, _18561_);
  and _67126_ (_21543_, _21216_, _18555_);
  nor _67127_ (_21544_, _21543_, _21542_);
  nor _67128_ (_21545_, _21544_, _18699_);
  or _67129_ (_21546_, _21545_, _21541_);
  and _67130_ (_21547_, _21546_, _18752_);
  nor _67131_ (_21548_, _21547_, _21537_);
  nor _67132_ (_21549_, _21548_, _18741_);
  or _67133_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _21549_, _21527_);
  and _67134_ (_21550_, _15585_, iram_op1[6]);
  and _67135_ (_21551_, _15589_, iram_op1_reg[6]);
  or _67136_ (_21552_, _21551_, _21550_);
  and _67137_ (_00004_[6], _21552_, _38997_);
  and _67138_ (_21553_, _15585_, iram_op1[5]);
  and _67139_ (_21554_, _15589_, iram_op1_reg[5]);
  or _67140_ (_21555_, _21554_, _21553_);
  and _67141_ (_00004_[5], _21555_, _38997_);
  and _67142_ (_21556_, _15585_, iram_op1[4]);
  and _67143_ (_21557_, _15589_, iram_op1_reg[4]);
  or _67144_ (_21558_, _21557_, _21556_);
  and _67145_ (_00004_[4], _21558_, _38997_);
  and _67146_ (_21559_, _15585_, iram_op1[3]);
  and _67147_ (_21560_, _15589_, iram_op1_reg[3]);
  or _67148_ (_21561_, _21560_, _21559_);
  and _67149_ (_00004_[3], _21561_, _38997_);
  and _67150_ (_21562_, _15585_, iram_op1[2]);
  and _67151_ (_21563_, _15589_, iram_op1_reg[2]);
  or _67152_ (_21564_, _21563_, _21562_);
  and _67153_ (_00004_[2], _21564_, _38997_);
  and _67154_ (_21565_, _15585_, iram_op1[1]);
  not _67155_ (_21566_, iram_op1_reg[1]);
  nor _67156_ (_21567_, _15585_, _21566_);
  or _67157_ (_21568_, _21567_, _21565_);
  and _67158_ (_00004_[1], _21568_, _38997_);
  and _67159_ (_21569_, _15585_, iram_op1[0]);
  not _67160_ (_21570_, iram_op1_reg[0]);
  nor _67161_ (_21571_, _15585_, _21570_);
  or _67162_ (_21572_, _21571_, _21569_);
  and _67163_ (_00004_[0], _21572_, _38997_);
  and _67164_ (_21573_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not _67165_ (_21574_, pc_change_r);
  and _67166_ (_21575_, _21574_, acc_reg[6]);
  or _67167_ (_21576_, _21575_, _21573_);
  and _67168_ (_00000_[6], _21576_, _38997_);
  and _67169_ (_21577_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _67170_ (_21578_, _21574_, acc_reg[5]);
  or _67171_ (_21579_, _21578_, _21577_);
  and _67172_ (_00000_[5], _21579_, _38997_);
  and _67173_ (_21580_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _67174_ (_21581_, _21574_, acc_reg[4]);
  or _67175_ (_21582_, _21581_, _21580_);
  and _67176_ (_00000_[4], _21582_, _38997_);
  and _67177_ (_21583_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _67178_ (_21584_, _21574_, acc_reg[3]);
  or _67179_ (_21585_, _21584_, _21583_);
  and _67180_ (_00000_[3], _21585_, _38997_);
  and _67181_ (_21586_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _67182_ (_21587_, _21574_, acc_reg[2]);
  or _67183_ (_21588_, _21587_, _21586_);
  and _67184_ (_00000_[2], _21588_, _38997_);
  and _67185_ (_21589_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _67186_ (_21590_, _21574_, acc_reg[1]);
  or _67187_ (_21591_, _21590_, _21589_);
  and _67188_ (_00000_[1], _21591_, _38997_);
  and _67189_ (_21592_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _67190_ (_21593_, _21574_, acc_reg[0]);
  or _67191_ (_21594_, _21593_, _21592_);
  and _67192_ (_00000_[0], _21594_, _38997_);
  and _67193_ (_21595_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _67194_ (_21596_, _21595_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _67195_ (_21597_, _21596_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _67196_ (_21598_, _21596_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _67197_ (_21599_, _21598_, _21597_);
  not _67198_ (_21600_, _21599_);
  nor _67199_ (_21601_, _21595_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _67200_ (_21602_, _21596_, _21601_);
  and _67201_ (_21603_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], _16190_);
  and _67202_ (_21604_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _67203_ (_21605_, _16194_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _67204_ (_21606_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _67205_ (_21607_, _21606_, _21604_);
  nor _67206_ (_21608_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _67207_ (_21609_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _67208_ (_21610_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _67209_ (_21611_, _21610_, _21609_);
  and _67210_ (_21612_, _21611_, _21607_);
  nor _67211_ (_21613_, _21612_, _21602_);
  not _67212_ (_21614_, _21602_);
  and _67213_ (_21615_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _67214_ (_21616_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _67215_ (_21617_, _21616_, _21615_);
  and _67216_ (_21618_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _67217_ (_21619_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _67218_ (_21620_, _21619_, _21618_);
  and _67219_ (_21621_, _21620_, _21617_);
  nor _67220_ (_21622_, _21621_, _21614_);
  or _67221_ (_21623_, _21622_, _21613_);
  and _67222_ (_21624_, _21623_, _21600_);
  and _67223_ (_21625_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _67224_ (_21626_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _67225_ (_21627_, _21626_, _21625_);
  and _67226_ (_21628_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _67227_ (_21629_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _67228_ (_21630_, _21629_, _21628_);
  and _67229_ (_21631_, _21630_, _21627_);
  nor _67230_ (_21632_, _21631_, _21602_);
  and _67231_ (_21633_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _67232_ (_21634_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _67233_ (_21635_, _21634_, _21633_);
  and _67234_ (_21636_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _67235_ (_21637_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _67236_ (_21638_, _21637_, _21636_);
  and _67237_ (_21639_, _21638_, _21635_);
  nor _67238_ (_21640_, _21639_, _21614_);
  nor _67239_ (_21641_, _21640_, _21632_);
  nor _67240_ (_21642_, _21641_, _21600_);
  nor _67241_ (_21643_, _21642_, _21624_);
  not _67242_ (_21644_, _21643_);
  not _67243_ (_21645_, _21603_);
  nor _67244_ (_21646_, _21599_, _18609_);
  and _67245_ (_21647_, _21599_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _67246_ (_21648_, _21647_, _21646_);
  nor _67247_ (_21649_, _21648_, _21645_);
  or _67248_ (_21650_, _21649_, _21602_);
  not _67249_ (_21651_, _21595_);
  nor _67250_ (_21652_, _21599_, _18657_);
  and _67251_ (_21653_, _21599_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _67252_ (_21654_, _21653_, _21652_);
  nor _67253_ (_21655_, _21654_, _21651_);
  not _67254_ (_21656_, _21608_);
  nor _67255_ (_21657_, _21599_, _18635_);
  and _67256_ (_21658_, _21599_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _67257_ (_21659_, _21658_, _21657_);
  nor _67258_ (_21660_, _21659_, _21656_);
  not _67259_ (_21661_, _21605_);
  nor _67260_ (_21662_, _21599_, _18644_);
  and _67261_ (_21663_, _21599_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _67262_ (_21664_, _21663_, _21662_);
  nor _67263_ (_21665_, _21664_, _21661_);
  or _67264_ (_21666_, _21665_, _21660_);
  or _67265_ (_21667_, _21666_, _21655_);
  or _67266_ (_21668_, _21667_, _21650_);
  and _67267_ (_21669_, _21599_, _18622_);
  nor _67268_ (_21670_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _67269_ (_21671_, _21670_, _21645_);
  nor _67270_ (_21672_, _21671_, _21669_);
  or _67271_ (_21673_, _21672_, _21614_);
  and _67272_ (_21674_, _21599_, _18663_);
  nor _67273_ (_21675_, \oc8051_symbolic_cxrom1.regvalid [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _67274_ (_21676_, _21675_, _21651_);
  nor _67275_ (_21677_, _21676_, _21674_);
  and _67276_ (_21678_, _21599_, _18630_);
  nor _67277_ (_21679_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _67278_ (_21680_, _21679_, _21656_);
  nor _67279_ (_21681_, _21680_, _21678_);
  and _67280_ (_21682_, _21599_, _18651_);
  nor _67281_ (_21683_, \oc8051_symbolic_cxrom1.regvalid [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _67282_ (_21684_, _21683_, _21661_);
  nor _67283_ (_21685_, _21684_, _21682_);
  or _67284_ (_21686_, _21685_, _21681_);
  or _67285_ (_21687_, _21686_, _21677_);
  or _67286_ (_21688_, _21687_, _21673_);
  and _67287_ (_21689_, _21688_, _21668_);
  and _67288_ (_21690_, _21689_, _21644_);
  or _67289_ (_21691_, _21690_, _15589_);
  or _67290_ (_21692_, _15585_, op1_out_r[6]);
  and _67291_ (_21693_, _21692_, _38997_);
  and _67292_ (_00005_[6], _21693_, _21691_);
  and _67293_ (_21694_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _67294_ (_21695_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _67295_ (_21696_, _21695_, _21694_);
  and _67296_ (_21697_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _67297_ (_21698_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _67298_ (_21699_, _21698_, _21697_);
  and _67299_ (_21700_, _21699_, _21696_);
  and _67300_ (_21701_, _21700_, _21614_);
  and _67301_ (_21702_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _67302_ (_21703_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _67303_ (_21704_, _21703_, _21702_);
  and _67304_ (_21705_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _67305_ (_21706_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _67306_ (_21707_, _21706_, _21705_);
  and _67307_ (_21708_, _21707_, _21704_);
  and _67308_ (_21709_, _21708_, _21602_);
  or _67309_ (_21710_, _21709_, _21599_);
  nor _67310_ (_21711_, _21710_, _21701_);
  and _67311_ (_21712_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _67312_ (_21713_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _67313_ (_21714_, _21713_, _21712_);
  and _67314_ (_21715_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _67315_ (_21716_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _67316_ (_21717_, _21716_, _21715_);
  and _67317_ (_21718_, _21717_, _21714_);
  nor _67318_ (_21719_, _21718_, _21602_);
  and _67319_ (_21720_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _67320_ (_21721_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _67321_ (_21722_, _21721_, _21720_);
  and _67322_ (_21723_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _67323_ (_21724_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _67324_ (_21725_, _21724_, _21723_);
  and _67325_ (_21726_, _21725_, _21722_);
  nor _67326_ (_21727_, _21726_, _21614_);
  or _67327_ (_21728_, _21727_, _21719_);
  and _67328_ (_21729_, _21728_, _21599_);
  nor _67329_ (_21730_, _21729_, _21711_);
  not _67330_ (_21731_, _21730_);
  and _67331_ (_21732_, _21731_, _21689_);
  or _67332_ (_21733_, _21732_, _15589_);
  or _67333_ (_21734_, _15585_, op1_out_r[5]);
  and _67334_ (_21735_, _21734_, _38997_);
  and _67335_ (_00005_[5], _21735_, _21733_);
  and _67336_ (_21736_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _67337_ (_21737_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _67338_ (_21738_, _21737_, _21736_);
  and _67339_ (_21739_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _67340_ (_21740_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _67341_ (_21741_, _21740_, _21739_);
  and _67342_ (_21742_, _21741_, _21738_);
  and _67343_ (_21743_, _21742_, _21614_);
  and _67344_ (_21744_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _67345_ (_21745_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _67346_ (_21746_, _21745_, _21744_);
  and _67347_ (_21747_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _67348_ (_21748_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _67349_ (_21749_, _21748_, _21747_);
  and _67350_ (_21750_, _21749_, _21746_);
  and _67351_ (_21751_, _21750_, _21602_);
  or _67352_ (_21752_, _21751_, _21599_);
  nor _67353_ (_21753_, _21752_, _21743_);
  and _67354_ (_21754_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _67355_ (_21755_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _67356_ (_21756_, _21755_, _21754_);
  and _67357_ (_21757_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _67358_ (_21758_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _67359_ (_21759_, _21758_, _21757_);
  and _67360_ (_21760_, _21759_, _21756_);
  and _67361_ (_21761_, _21760_, _21614_);
  and _67362_ (_21762_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _67363_ (_21763_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _67364_ (_21764_, _21763_, _21762_);
  and _67365_ (_21765_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _67366_ (_21766_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _67367_ (_21767_, _21766_, _21765_);
  and _67368_ (_21768_, _21767_, _21764_);
  and _67369_ (_21769_, _21768_, _21602_);
  or _67370_ (_21770_, _21769_, _21600_);
  nor _67371_ (_21771_, _21770_, _21761_);
  nor _67372_ (_21772_, _21771_, _21753_);
  not _67373_ (_21773_, _21772_);
  and _67374_ (_21774_, _21773_, _21689_);
  or _67375_ (_21775_, _21774_, _15589_);
  or _67376_ (_21776_, _15585_, op1_out_r[4]);
  and _67377_ (_21777_, _21776_, _38997_);
  and _67378_ (_00005_[4], _21777_, _21775_);
  and _67379_ (_21778_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _67380_ (_21779_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _67381_ (_21780_, _21779_, _21778_);
  and _67382_ (_21781_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and _67383_ (_21782_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _67384_ (_21783_, _21782_, _21781_);
  and _67385_ (_21784_, _21783_, _21780_);
  nor _67386_ (_21785_, _21784_, _21602_);
  and _67387_ (_21786_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _67388_ (_21787_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _67389_ (_21788_, _21787_, _21786_);
  and _67390_ (_21789_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _67391_ (_21790_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _67392_ (_21791_, _21790_, _21789_);
  and _67393_ (_21792_, _21791_, _21788_);
  nor _67394_ (_21793_, _21792_, _21614_);
  or _67395_ (_21794_, _21793_, _21785_);
  and _67396_ (_21795_, _21794_, _21600_);
  and _67397_ (_21796_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _67398_ (_21797_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _67399_ (_21798_, _21797_, _21796_);
  and _67400_ (_21799_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _67401_ (_21800_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _67402_ (_21801_, _21800_, _21799_);
  and _67403_ (_21802_, _21801_, _21798_);
  nor _67404_ (_21803_, _21802_, _21602_);
  and _67405_ (_21804_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _67406_ (_21805_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor _67407_ (_21806_, _21805_, _21804_);
  and _67408_ (_21807_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _67409_ (_21808_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _67410_ (_21809_, _21808_, _21807_);
  and _67411_ (_21810_, _21809_, _21806_);
  nor _67412_ (_21811_, _21810_, _21614_);
  or _67413_ (_21812_, _21811_, _21803_);
  and _67414_ (_21813_, _21812_, _21599_);
  nor _67415_ (_21814_, _21813_, _21795_);
  not _67416_ (_21815_, _21814_);
  and _67417_ (_21816_, _21815_, _21689_);
  or _67418_ (_21817_, _21816_, _15589_);
  or _67419_ (_21818_, _15585_, op1_out_r[3]);
  and _67420_ (_21819_, _21818_, _38997_);
  and _67421_ (_00005_[3], _21819_, _21817_);
  and _67422_ (_21820_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _67423_ (_21821_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _67424_ (_21822_, _21821_, _21820_);
  and _67425_ (_21823_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _67426_ (_21824_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _67427_ (_21825_, _21824_, _21823_);
  and _67428_ (_21826_, _21825_, _21822_);
  and _67429_ (_21827_, _21826_, _21602_);
  and _67430_ (_21828_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _67431_ (_21829_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _67432_ (_21830_, _21829_, _21828_);
  and _67433_ (_21831_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _67434_ (_21832_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _67435_ (_21833_, _21832_, _21831_);
  and _67436_ (_21834_, _21833_, _21830_);
  and _67437_ (_21835_, _21834_, _21614_);
  nor _67438_ (_21836_, _21835_, _21827_);
  nor _67439_ (_21837_, _21836_, _21600_);
  and _67440_ (_21838_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _67441_ (_21839_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _67442_ (_21840_, _21839_, _21838_);
  and _67443_ (_21841_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _67444_ (_21842_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _67445_ (_21843_, _21842_, _21841_);
  and _67446_ (_21844_, _21843_, _21840_);
  and _67447_ (_21845_, _21844_, _21614_);
  and _67448_ (_21846_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _67449_ (_21847_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _67450_ (_21848_, _21847_, _21846_);
  and _67451_ (_21849_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _67452_ (_21850_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _67453_ (_21851_, _21850_, _21849_);
  and _67454_ (_21852_, _21851_, _21848_);
  and _67455_ (_21853_, _21852_, _21602_);
  nor _67456_ (_21854_, _21853_, _21845_);
  nor _67457_ (_21855_, _21854_, _21599_);
  nor _67458_ (_21856_, _21855_, _21837_);
  and _67459_ (_21857_, _21856_, _21689_);
  or _67460_ (_21858_, _21857_, _15589_);
  or _67461_ (_21859_, _15585_, op1_out_r[2]);
  and _67462_ (_21860_, _21859_, _38997_);
  and _67463_ (_00005_[2], _21860_, _21858_);
  and _67464_ (_21861_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _67465_ (_21862_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _67466_ (_21863_, _21862_, _21861_);
  and _67467_ (_21864_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _67468_ (_21865_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _67469_ (_21866_, _21865_, _21864_);
  and _67470_ (_21867_, _21866_, _21863_);
  and _67471_ (_21868_, _21867_, _21614_);
  and _67472_ (_21869_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _67473_ (_21870_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _67474_ (_21871_, _21870_, _21869_);
  and _67475_ (_21872_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _67476_ (_21873_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _67477_ (_21874_, _21873_, _21872_);
  and _67478_ (_21875_, _21874_, _21871_);
  and _67479_ (_21876_, _21875_, _21602_);
  nor _67480_ (_21877_, _21876_, _21868_);
  nor _67481_ (_21878_, _21877_, _21600_);
  and _67482_ (_21879_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _67483_ (_21880_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _67484_ (_21881_, _21880_, _21879_);
  and _67485_ (_21882_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _67486_ (_21883_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _67487_ (_21884_, _21883_, _21882_);
  and _67488_ (_21885_, _21884_, _21881_);
  and _67489_ (_21886_, _21885_, _21614_);
  and _67490_ (_21887_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _67491_ (_21888_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _67492_ (_21889_, _21888_, _21887_);
  and _67493_ (_21890_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _67494_ (_21891_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _67495_ (_21892_, _21891_, _21890_);
  and _67496_ (_21893_, _21892_, _21889_);
  and _67497_ (_21894_, _21893_, _21602_);
  nor _67498_ (_21895_, _21894_, _21886_);
  nor _67499_ (_21896_, _21895_, _21599_);
  nor _67500_ (_21897_, _21896_, _21878_);
  and _67501_ (_21898_, _21897_, _21689_);
  or _67502_ (_21899_, _21898_, _15589_);
  or _67503_ (_21900_, _15585_, op1_out_r[1]);
  and _67504_ (_21901_, _21900_, _38997_);
  and _67505_ (_00005_[1], _21901_, _21899_);
  and _67506_ (_21902_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _67507_ (_21903_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor _67508_ (_21904_, _21903_, _21902_);
  and _67509_ (_21905_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _67510_ (_21906_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _67511_ (_21907_, _21906_, _21905_);
  and _67512_ (_21908_, _21907_, _21904_);
  and _67513_ (_21909_, _21908_, _21614_);
  and _67514_ (_21910_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _67515_ (_21911_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _67516_ (_21912_, _21911_, _21910_);
  and _67517_ (_21913_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _67518_ (_21914_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _67519_ (_21915_, _21914_, _21913_);
  and _67520_ (_21916_, _21915_, _21912_);
  and _67521_ (_21917_, _21916_, _21602_);
  or _67522_ (_21918_, _21917_, _21599_);
  nor _67523_ (_21919_, _21918_, _21909_);
  and _67524_ (_21920_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _67525_ (_21921_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor _67526_ (_21922_, _21921_, _21920_);
  and _67527_ (_21923_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _67528_ (_21924_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _67529_ (_21925_, _21924_, _21923_);
  and _67530_ (_21926_, _21925_, _21922_);
  and _67531_ (_21927_, _21926_, _21614_);
  and _67532_ (_21928_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _67533_ (_21929_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _67534_ (_21930_, _21929_, _21928_);
  and _67535_ (_21931_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _67536_ (_21932_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _67537_ (_21933_, _21932_, _21931_);
  and _67538_ (_21934_, _21933_, _21930_);
  and _67539_ (_21935_, _21934_, _21602_);
  or _67540_ (_21936_, _21935_, _21600_);
  nor _67541_ (_21937_, _21936_, _21927_);
  nor _67542_ (_21938_, _21937_, _21919_);
  not _67543_ (_21939_, _21938_);
  and _67544_ (_21940_, _21939_, _21689_);
  or _67545_ (_21941_, _21940_, _15589_);
  or _67546_ (_21942_, _15585_, op1_out_r[0]);
  and _67547_ (_21943_, _21942_, _38997_);
  and _67548_ (_00005_[0], _21943_, _21941_);
  and _67549_ (_21944_, _15589_, iram_op1[6]);
  and _67550_ (_21945_, _21774_, _21732_);
  and _67551_ (_21946_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _67552_ (_21947_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor _67553_ (_21948_, _21947_, _21946_);
  and _67554_ (_21949_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _67555_ (_21950_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor _67556_ (_21951_, _21950_, _21949_);
  and _67557_ (_21952_, _21951_, _21948_);
  and _67558_ (_21953_, _21952_, _21614_);
  and _67559_ (_21954_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _67560_ (_21955_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _67561_ (_21956_, _21955_, _21954_);
  and _67562_ (_21957_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _67563_ (_21958_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _67564_ (_21959_, _21958_, _21957_);
  and _67565_ (_21960_, _21959_, _21956_);
  and _67566_ (_21961_, _21960_, _21602_);
  nor _67567_ (_21962_, _21961_, _21953_);
  nor _67568_ (_21963_, _21962_, _21600_);
  and _67569_ (_21964_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _67570_ (_21965_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor _67571_ (_21966_, _21965_, _21964_);
  and _67572_ (_21967_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _67573_ (_21968_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _67574_ (_21969_, _21968_, _21967_);
  and _67575_ (_21970_, _21969_, _21966_);
  and _67576_ (_21971_, _21970_, _21614_);
  and _67577_ (_21972_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _67578_ (_21973_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor _67579_ (_21974_, _21973_, _21972_);
  and _67580_ (_21975_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _67581_ (_21976_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _67582_ (_21977_, _21976_, _21975_);
  and _67583_ (_21978_, _21977_, _21974_);
  and _67584_ (_21979_, _21978_, _21602_);
  nor _67585_ (_21980_, _21979_, _21971_);
  nor _67586_ (_21981_, _21980_, _21599_);
  nor _67587_ (_21982_, _21981_, _21963_);
  and _67588_ (_21983_, _21982_, _21689_);
  and _67589_ (_21984_, _21983_, _21690_);
  and _67590_ (_21985_, _21984_, _21945_);
  nor _67591_ (_21986_, _21857_, _21816_);
  and _67592_ (_21987_, _21938_, _21898_);
  and _67593_ (_21988_, _21987_, _21986_);
  and _67594_ (_21989_, _21988_, _21985_);
  and _67595_ (_21990_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  not _67596_ (_21991_, _21898_);
  and _67597_ (_21992_, _21940_, _21991_);
  and _67598_ (_21993_, _21986_, _21992_);
  and _67599_ (_21994_, _21993_, _21985_);
  and _67600_ (_21995_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or _67601_ (_21996_, _21995_, _21990_);
  nor _67602_ (_21997_, _21940_, _21898_);
  and _67603_ (_21998_, _21986_, _21997_);
  and _67604_ (_21999_, _21998_, _21985_);
  and _67605_ (_22000_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and _67606_ (_22001_, _21857_, _21816_);
  and _67607_ (_22002_, _21940_, _21898_);
  and _67608_ (_22003_, _22002_, _22001_);
  and _67609_ (_22004_, _21772_, _21732_);
  and _67610_ (_22005_, _22004_, _21984_);
  and _67611_ (_22006_, _22005_, _22003_);
  and _67612_ (_22007_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  or _67613_ (_22008_, _22007_, _22000_);
  or _67614_ (_22009_, _22008_, _21996_);
  not _67615_ (_22010_, _21816_);
  and _67616_ (_22011_, _21857_, _22010_);
  and _67617_ (_22012_, _22011_, _21992_);
  and _67618_ (_22013_, _22012_, _21985_);
  and _67619_ (_22014_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  and _67620_ (_22015_, _21987_, _22011_);
  and _67621_ (_22016_, _22015_, _21985_);
  and _67622_ (_22017_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or _67623_ (_22018_, _22017_, _22014_);
  and _67624_ (_22019_, _22011_, _21997_);
  and _67625_ (_22020_, _22019_, _21985_);
  and _67626_ (_22021_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and _67627_ (_22022_, _21986_, _22002_);
  and _67628_ (_22023_, _22022_, _21985_);
  and _67629_ (_22024_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  or _67630_ (_22025_, _22024_, _22021_);
  or _67631_ (_22026_, _22025_, _22018_);
  or _67632_ (_22027_, _22026_, _22009_);
  and _67633_ (_22028_, _21987_, _22001_);
  and _67634_ (_22029_, _22028_, _21985_);
  and _67635_ (_22030_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and _67636_ (_22031_, _21992_, _22001_);
  and _67637_ (_22032_, _22031_, _21985_);
  and _67638_ (_22033_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  or _67639_ (_22034_, _22033_, _22030_);
  and _67640_ (_22035_, _22001_, _21997_);
  and _67641_ (_22036_, _22035_, _21985_);
  and _67642_ (_22037_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  nor _67643_ (_22038_, _21857_, _22010_);
  and _67644_ (_22039_, _22002_, _22038_);
  and _67645_ (_22040_, _22039_, _21985_);
  and _67646_ (_22041_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or _67647_ (_22042_, _22041_, _22037_);
  or _67648_ (_22043_, _22042_, _22034_);
  and _67649_ (_22044_, _21987_, _22038_);
  and _67650_ (_22045_, _22044_, _21985_);
  and _67651_ (_22046_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and _67652_ (_22047_, _21992_, _22038_);
  and _67653_ (_22048_, _22047_, _21985_);
  and _67654_ (_22049_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  or _67655_ (_22050_, _22049_, _22046_);
  and _67656_ (_22051_, _22038_, _21997_);
  and _67657_ (_22052_, _22051_, _21985_);
  and _67658_ (_22053_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  and _67659_ (_22054_, _22011_, _22002_);
  and _67660_ (_22055_, _22054_, _21985_);
  and _67661_ (_22056_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  or _67662_ (_22057_, _22056_, _22053_);
  or _67663_ (_22058_, _22057_, _22050_);
  or _67664_ (_22059_, _22058_, _22043_);
  or _67665_ (_22060_, _22059_, _22027_);
  and _67666_ (_22061_, _22005_, _21993_);
  and _67667_ (_22062_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and _67668_ (_22063_, _22005_, _21988_);
  and _67669_ (_22064_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  or _67670_ (_22065_, _22064_, _22062_);
  and _67671_ (_22066_, _21774_, _21730_);
  and _67672_ (_22067_, _22066_, _21984_);
  and _67673_ (_22068_, _22067_, _22003_);
  and _67674_ (_22069_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  and _67675_ (_22070_, _22005_, _21998_);
  and _67676_ (_22071_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or _67677_ (_22072_, _22071_, _22069_);
  or _67678_ (_22073_, _22072_, _22065_);
  and _67679_ (_22074_, _22005_, _22015_);
  and _67680_ (_22075_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and _67681_ (_22076_, _22005_, _22012_);
  and _67682_ (_22077_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  or _67683_ (_22078_, _22077_, _22075_);
  and _67684_ (_22079_, _22005_, _22022_);
  and _67685_ (_22080_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  and _67686_ (_22081_, _22005_, _22019_);
  and _67687_ (_22082_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or _67688_ (_22083_, _22082_, _22080_);
  or _67689_ (_22084_, _22083_, _22078_);
  or _67690_ (_22085_, _22084_, _22073_);
  and _67691_ (_22086_, _22005_, _22031_);
  and _67692_ (_22087_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  and _67693_ (_22088_, _22005_, _22028_);
  and _67694_ (_22089_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or _67695_ (_22090_, _22089_, _22087_);
  and _67696_ (_22091_, _22005_, _22039_);
  and _67697_ (_22092_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and _67698_ (_22093_, _22005_, _22035_);
  and _67699_ (_22094_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  or _67700_ (_22095_, _22094_, _22092_);
  or _67701_ (_22096_, _22095_, _22090_);
  and _67702_ (_22097_, _22005_, _22044_);
  and _67703_ (_22098_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  and _67704_ (_22099_, _22005_, _22047_);
  and _67705_ (_22100_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or _67706_ (_22101_, _22100_, _22098_);
  and _67707_ (_22102_, _22005_, _22051_);
  and _67708_ (_22103_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and _67709_ (_22104_, _22005_, _22054_);
  and _67710_ (_22105_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or _67711_ (_22106_, _22105_, _22103_);
  or _67712_ (_22107_, _22106_, _22101_);
  or _67713_ (_22108_, _22107_, _22096_);
  or _67714_ (_22109_, _22108_, _22085_);
  or _67715_ (_22110_, _22109_, _22060_);
  and _67716_ (_22111_, _22067_, _22028_);
  and _67717_ (_22112_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and _67718_ (_22113_, _22067_, _22031_);
  and _67719_ (_22114_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  or _67720_ (_22115_, _22114_, _22112_);
  and _67721_ (_22116_, _22067_, _22039_);
  and _67722_ (_22117_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  and _67723_ (_22118_, _22067_, _22035_);
  and _67724_ (_22119_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or _67725_ (_22120_, _22119_, _22117_);
  or _67726_ (_22121_, _22120_, _22115_);
  and _67727_ (_22122_, _22067_, _22044_);
  and _67728_ (_22123_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and _67729_ (_22124_, _22067_, _22047_);
  and _67730_ (_22125_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  or _67731_ (_22126_, _22125_, _22123_);
  and _67732_ (_22127_, _22067_, _22051_);
  and _67733_ (_22128_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  and _67734_ (_22129_, _22067_, _22054_);
  and _67735_ (_22130_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  or _67736_ (_22131_, _22130_, _22128_);
  or _67737_ (_22132_, _22131_, _22126_);
  or _67738_ (_22133_, _22132_, _22121_);
  and _67739_ (_22134_, _22067_, _21993_);
  and _67740_ (_22135_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  and _67741_ (_22136_, _22067_, _21988_);
  and _67742_ (_22137_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or _67743_ (_22138_, _22137_, _22135_);
  nor _67744_ (_22139_, _21774_, _21732_);
  and _67745_ (_22140_, _22139_, _21984_);
  and _67746_ (_22141_, _22003_, _22140_);
  and _67747_ (_22142_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and _67748_ (_22143_, _22067_, _21998_);
  and _67749_ (_22144_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  or _67750_ (_22145_, _22144_, _22142_);
  or _67751_ (_22146_, _22145_, _22138_);
  and _67752_ (_22147_, _22067_, _22015_);
  and _67753_ (_22148_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  and _67754_ (_22149_, _22067_, _22012_);
  and _67755_ (_22150_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or _67756_ (_22151_, _22150_, _22148_);
  and _67757_ (_22152_, _22067_, _22019_);
  and _67758_ (_22153_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and _67759_ (_22154_, _22067_, _22022_);
  and _67760_ (_22155_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  or _67761_ (_22156_, _22155_, _22153_);
  or _67762_ (_22157_, _22156_, _22151_);
  or _67763_ (_22158_, _22157_, _22146_);
  or _67764_ (_22159_, _22158_, _22133_);
  and _67765_ (_22160_, _22031_, _22140_);
  and _67766_ (_22161_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  and _67767_ (_22162_, _22028_, _22140_);
  and _67768_ (_22163_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or _67769_ (_22164_, _22163_, _22161_);
  and _67770_ (_22165_, _22039_, _22140_);
  and _67771_ (_22166_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and _67772_ (_22167_, _22140_, _22035_);
  and _67773_ (_22168_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  or _67774_ (_22169_, _22168_, _22166_);
  or _67775_ (_22170_, _22169_, _22164_);
  and _67776_ (_22171_, _22047_, _22140_);
  and _67777_ (_22172_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  and _67778_ (_22173_, _22044_, _22140_);
  and _67779_ (_22174_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or _67780_ (_22175_, _22174_, _22172_);
  and _67781_ (_22176_, _22140_, _22051_);
  and _67782_ (_22177_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and _67783_ (_22178_, _22054_, _22140_);
  and _67784_ (_22179_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or _67785_ (_22180_, _22179_, _22177_);
  or _67786_ (_22181_, _22180_, _22175_);
  or _67787_ (_22182_, _22181_, _22170_);
  and _67788_ (_22183_, _22015_, _22140_);
  and _67789_ (_22184_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and _67790_ (_22185_, _22012_, _22140_);
  and _67791_ (_22186_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  or _67792_ (_22187_, _22186_, _22184_);
  and _67793_ (_22188_, _22022_, _22140_);
  and _67794_ (_22189_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  and _67795_ (_22190_, _22019_, _22140_);
  and _67796_ (_22191_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or _67797_ (_22192_, _22191_, _22189_);
  or _67798_ (_22193_, _22192_, _22187_);
  and _67799_ (_22194_, _21988_, _22140_);
  and _67800_ (_22195_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and _67801_ (_22196_, _21993_, _22140_);
  and _67802_ (_22197_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  or _67803_ (_22198_, _22197_, _22195_);
  not _67804_ (_22199_, _21983_);
  nor _67805_ (_22200_, _22199_, _21690_);
  and _67806_ (_22201_, _22200_, _21945_);
  and _67807_ (_22202_, _22201_, _22003_);
  and _67808_ (_22203_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  and _67809_ (_22204_, _21998_, _22140_);
  and _67810_ (_22205_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or _67811_ (_22206_, _22205_, _22203_);
  or _67812_ (_22207_, _22206_, _22198_);
  or _67813_ (_22208_, _22207_, _22193_);
  or _67814_ (_22209_, _22208_, _22182_);
  or _67815_ (_22210_, _22209_, _22159_);
  or _67816_ (_22211_, _22210_, _22110_);
  and _67817_ (_22212_, _22201_, _22012_);
  and _67818_ (_22213_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  and _67819_ (_22214_, _22201_, _22015_);
  and _67820_ (_22215_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or _67821_ (_22216_, _22215_, _22213_);
  and _67822_ (_22217_, _22201_, _22019_);
  and _67823_ (_22218_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and _67824_ (_22219_, _22201_, _22022_);
  and _67825_ (_22220_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  or _67826_ (_22221_, _22220_, _22218_);
  or _67827_ (_22222_, _22221_, _22216_);
  and _67828_ (_22223_, _22201_, _21993_);
  and _67829_ (_22224_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  and _67830_ (_22225_, _22201_, _21988_);
  and _67831_ (_22226_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or _67832_ (_22227_, _22226_, _22224_);
  and _67833_ (_22228_, _22004_, _22200_);
  and _67834_ (_22229_, _22003_, _22228_);
  and _67835_ (_22230_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and _67836_ (_22231_, _22201_, _21998_);
  and _67837_ (_22232_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  or _67838_ (_22233_, _22232_, _22230_);
  or _67839_ (_22234_, _22233_, _22227_);
  or _67840_ (_22235_, _22234_, _22222_);
  and _67841_ (_22236_, _22201_, _22044_);
  and _67842_ (_22237_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and _67843_ (_22238_, _22201_, _22047_);
  and _67844_ (_22239_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  or _67845_ (_22240_, _22239_, _22237_);
  and _67846_ (_22241_, _22201_, _22051_);
  and _67847_ (_22242_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  and _67848_ (_22243_, _22201_, _22054_);
  and _67849_ (_22244_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  or _67850_ (_22245_, _22244_, _22242_);
  or _67851_ (_22246_, _22245_, _22240_);
  and _67852_ (_22247_, _22201_, _22028_);
  and _67853_ (_22248_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and _67854_ (_22249_, _22201_, _22031_);
  and _67855_ (_22250_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  or _67856_ (_22251_, _22250_, _22248_);
  and _67857_ (_22252_, _22201_, _22039_);
  and _67858_ (_22253_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  and _67859_ (_22254_, _22201_, _22035_);
  and _67860_ (_22255_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or _67861_ (_22256_, _22255_, _22253_);
  or _67862_ (_22257_, _22256_, _22251_);
  or _67863_ (_22258_, _22257_, _22246_);
  or _67864_ (_22259_, _22258_, _22235_);
  and _67865_ (_22260_, _22047_, _22228_);
  and _67866_ (_22261_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  and _67867_ (_22262_, _22044_, _22228_);
  and _67868_ (_22263_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or _67869_ (_22264_, _22263_, _22261_);
  and _67870_ (_22265_, _22054_, _22228_);
  and _67871_ (_22266_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  and _67872_ (_22267_, _22228_, _22051_);
  and _67873_ (_22268_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  or _67874_ (_22269_, _22268_, _22266_);
  or _67875_ (_22270_, _22269_, _22264_);
  and _67876_ (_22271_, _22228_, _22031_);
  and _67877_ (_22272_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  and _67878_ (_22273_, _22028_, _22228_);
  and _67879_ (_22274_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or _67880_ (_22275_, _22274_, _22272_);
  and _67881_ (_22276_, _22228_, _22039_);
  and _67882_ (_22277_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and _67883_ (_22278_, _22228_, _22035_);
  and _67884_ (_22279_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  or _67885_ (_22280_, _22279_, _22277_);
  or _67886_ (_22281_, _22280_, _22275_);
  or _67887_ (_22282_, _22281_, _22270_);
  and _67888_ (_22283_, _22012_, _22228_);
  and _67889_ (_22284_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and _67890_ (_22285_, _22015_, _22228_);
  and _67891_ (_22286_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  or _67892_ (_22287_, _22286_, _22284_);
  and _67893_ (_22288_, _22022_, _22228_);
  and _67894_ (_22289_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  and _67895_ (_22290_, _22019_, _22228_);
  and _67896_ (_22291_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or _67897_ (_22292_, _22291_, _22289_);
  or _67898_ (_22293_, _22292_, _22287_);
  and _67899_ (_22294_, _21988_, _22228_);
  and _67900_ (_22295_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and _67901_ (_22296_, _21993_, _22228_);
  and _67902_ (_22297_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  or _67903_ (_22298_, _22297_, _22295_);
  and _67904_ (_22299_, _22066_, _22200_);
  and _67905_ (_22300_, _22299_, _22003_);
  and _67906_ (_22301_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  and _67907_ (_22302_, _21998_, _22228_);
  and _67908_ (_22303_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or _67909_ (_22304_, _22303_, _22301_);
  or _67910_ (_22305_, _22304_, _22298_);
  or _67911_ (_22306_, _22305_, _22293_);
  or _67912_ (_22307_, _22306_, _22282_);
  or _67913_ (_22308_, _22307_, _22259_);
  and _67914_ (_22309_, _22299_, _21988_);
  and _67915_ (_22310_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  and _67916_ (_22311_, _22299_, _21993_);
  and _67917_ (_22312_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or _67918_ (_22313_, _22312_, _22310_);
  and _67919_ (_22314_, _22299_, _21998_);
  and _67920_ (_22315_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and _67921_ (_22316_, _22200_, _22139_);
  and _67922_ (_22317_, _22003_, _22316_);
  and _67923_ (_22318_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  or _67924_ (_22319_, _22318_, _22315_);
  or _67925_ (_22320_, _22319_, _22313_);
  and _67926_ (_22321_, _22299_, _22015_);
  and _67927_ (_22322_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  and _67928_ (_22323_, _22299_, _22012_);
  and _67929_ (_22324_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or _67930_ (_22325_, _22324_, _22322_);
  and _67931_ (_22326_, _22299_, _22019_);
  and _67932_ (_22327_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and _67933_ (_22328_, _22299_, _22022_);
  and _67934_ (_22329_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  or _67935_ (_22330_, _22329_, _22327_);
  or _67936_ (_22331_, _22330_, _22325_);
  or _67937_ (_22332_, _22331_, _22320_);
  and _67938_ (_22333_, _22299_, _22031_);
  and _67939_ (_22334_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and _67940_ (_22335_, _22299_, _22028_);
  and _67941_ (_22336_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  or _67942_ (_22337_, _22336_, _22334_);
  and _67943_ (_22338_, _22299_, _22035_);
  and _67944_ (_22339_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  and _67945_ (_22340_, _22299_, _22039_);
  and _67946_ (_22341_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or _67947_ (_22342_, _22341_, _22339_);
  or _67948_ (_22343_, _22342_, _22337_);
  and _67949_ (_22344_, _22299_, _22047_);
  and _67950_ (_22345_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and _67951_ (_22346_, _22299_, _22044_);
  and _67952_ (_22347_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  or _67953_ (_22348_, _22347_, _22345_);
  and _67954_ (_22349_, _22299_, _22051_);
  and _67955_ (_22350_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  and _67956_ (_22351_, _22299_, _22054_);
  and _67957_ (_22352_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  or _67958_ (_22353_, _22352_, _22350_);
  or _67959_ (_22354_, _22353_, _22348_);
  or _67960_ (_22355_, _22354_, _22343_);
  or _67961_ (_22356_, _22355_, _22332_);
  and _67962_ (_22357_, _21993_, _22316_);
  and _67963_ (_22358_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and _67964_ (_22359_, _21988_, _22316_);
  and _67965_ (_22360_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  or _67966_ (_22361_, _22360_, _22358_);
  and _67967_ (_22362_, _21998_, _22316_);
  and _67968_ (_22363_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  and _67969_ (_22364_, _22199_, _21690_);
  and _67970_ (_22365_, _22364_, _21945_);
  and _67971_ (_22366_, _22003_, _22365_);
  and _67972_ (_22367_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or _67973_ (_22368_, _22367_, _22363_);
  or _67974_ (_22369_, _22368_, _22361_);
  and _67975_ (_22370_, _22015_, _22316_);
  and _67976_ (_22371_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and _67977_ (_22372_, _22012_, _22316_);
  and _67978_ (_22373_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  or _67979_ (_22374_, _22373_, _22371_);
  and _67980_ (_22375_, _22019_, _22316_);
  and _67981_ (_22376_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  and _67982_ (_22377_, _22022_, _22316_);
  and _67983_ (_22378_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or _67984_ (_22379_, _22378_, _22376_);
  or _67985_ (_22380_, _22379_, _22374_);
  or _67986_ (_22381_, _22380_, _22369_);
  and _67987_ (_22382_, _22031_, _22316_);
  and _67988_ (_22383_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  and _67989_ (_22384_, _22028_, _22316_);
  and _67990_ (_22385_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or _67991_ (_22386_, _22385_, _22383_);
  and _67992_ (_22387_, _22316_, _22035_);
  and _67993_ (_22388_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and _67994_ (_22389_, _22039_, _22316_);
  and _67995_ (_22390_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  or _67996_ (_22391_, _22390_, _22388_);
  or _67997_ (_22392_, _22391_, _22386_);
  and _67998_ (_22393_, _22044_, _22316_);
  and _67999_ (_22394_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  and _68000_ (_22395_, _22047_, _22316_);
  and _68001_ (_22396_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or _68002_ (_22397_, _22396_, _22394_);
  and _68003_ (_22398_, _22054_, _22316_);
  and _68004_ (_22399_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  and _68005_ (_22400_, _22316_, _22051_);
  and _68006_ (_22401_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  or _68007_ (_22402_, _22401_, _22399_);
  or _68008_ (_22403_, _22402_, _22397_);
  or _68009_ (_22404_, _22403_, _22392_);
  or _68010_ (_22405_, _22404_, _22381_);
  or _68011_ (_22406_, _22405_, _22356_);
  or _68012_ (_22407_, _22406_, _22308_);
  or _68013_ (_22408_, _22407_, _22211_);
  and _68014_ (_22409_, _22365_, _22012_);
  and _68015_ (_22410_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  and _68016_ (_22411_, _22365_, _22015_);
  and _68017_ (_22412_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or _68018_ (_22413_, _22412_, _22410_);
  and _68019_ (_22414_, _22365_, _22019_);
  and _68020_ (_22415_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and _68021_ (_22416_, _22365_, _22022_);
  and _68022_ (_22417_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  or _68023_ (_22418_, _22417_, _22415_);
  or _68024_ (_22419_, _22418_, _22413_);
  and _68025_ (_22420_, _22365_, _21993_);
  and _68026_ (_22421_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  and _68027_ (_22422_, _21988_, _22365_);
  and _68028_ (_22423_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or _68029_ (_22424_, _22423_, _22421_);
  and _68030_ (_22425_, _22364_, _22004_);
  and _68031_ (_22426_, _22003_, _22425_);
  and _68032_ (_22427_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and _68033_ (_22428_, _22365_, _21998_);
  and _68034_ (_22429_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  or _68035_ (_22430_, _22429_, _22427_);
  or _68036_ (_22431_, _22430_, _22424_);
  or _68037_ (_22432_, _22431_, _22419_);
  and _68038_ (_22433_, _22365_, _22044_);
  and _68039_ (_22434_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and _68040_ (_22435_, _22365_, _22047_);
  and _68041_ (_22436_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  or _68042_ (_22437_, _22436_, _22434_);
  and _68043_ (_22438_, _22365_, _22054_);
  and _68044_ (_22439_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and _68045_ (_22440_, _22365_, _22051_);
  and _68046_ (_22441_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or _68047_ (_22442_, _22441_, _22439_);
  or _68048_ (_22443_, _22442_, _22437_);
  and _68049_ (_22444_, _22365_, _22028_);
  and _68050_ (_22445_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and _68051_ (_22446_, _22365_, _22031_);
  and _68052_ (_22447_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  or _68053_ (_22448_, _22447_, _22445_);
  and _68054_ (_22449_, _22365_, _22039_);
  and _68055_ (_22450_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  and _68056_ (_22451_, _22365_, _22035_);
  and _68057_ (_22452_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or _68058_ (_22453_, _22452_, _22450_);
  or _68059_ (_22454_, _22453_, _22448_);
  or _68060_ (_22455_, _22454_, _22443_);
  or _68061_ (_22456_, _22455_, _22432_);
  and _68062_ (_22457_, _22425_, _22028_);
  and _68063_ (_22458_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  and _68064_ (_22459_, _22425_, _22031_);
  and _68065_ (_22460_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or _68066_ (_22461_, _22460_, _22458_);
  and _68067_ (_22462_, _22425_, _22035_);
  and _68068_ (_22463_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and _68069_ (_22464_, _22425_, _22039_);
  and _68070_ (_22465_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  or _68071_ (_22466_, _22465_, _22463_);
  or _68072_ (_22467_, _22466_, _22461_);
  and _68073_ (_22468_, _22425_, _22044_);
  and _68074_ (_22469_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  and _68075_ (_22470_, _22425_, _22047_);
  and _68076_ (_22471_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or _68077_ (_22472_, _22471_, _22469_);
  and _68078_ (_22473_, _22425_, _22051_);
  and _68079_ (_22474_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and _68080_ (_22475_, _22425_, _22054_);
  and _68081_ (_22476_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or _68082_ (_22477_, _22476_, _22474_);
  or _68083_ (_22478_, _22477_, _22472_);
  or _68084_ (_22479_, _22478_, _22467_);
  and _68085_ (_22480_, _22425_, _22012_);
  and _68086_ (_22481_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and _68087_ (_22482_, _22425_, _22015_);
  and _68088_ (_22483_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  or _68089_ (_22484_, _22483_, _22481_);
  and _68090_ (_22485_, _22019_, _22425_);
  and _68091_ (_22486_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  and _68092_ (_22487_, _22425_, _22022_);
  and _68093_ (_22488_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or _68094_ (_22489_, _22488_, _22486_);
  or _68095_ (_22490_, _22489_, _22484_);
  and _68096_ (_22491_, _21988_, _22425_);
  and _68097_ (_22492_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and _68098_ (_22493_, _22425_, _21993_);
  and _68099_ (_22494_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  or _68100_ (_22495_, _22494_, _22492_);
  and _68101_ (_22496_, _21998_, _22425_);
  and _68102_ (_22497_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  and _68103_ (_22498_, _22364_, _22066_);
  and _68104_ (_22499_, _22003_, _22498_);
  and _68105_ (_22500_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or _68106_ (_22501_, _22500_, _22497_);
  or _68107_ (_22502_, _22501_, _22495_);
  or _68108_ (_22503_, _22502_, _22490_);
  or _68109_ (_22504_, _22503_, _22479_);
  or _68110_ (_22505_, _22504_, _22456_);
  and _68111_ (_22506_, _22012_, _22498_);
  and _68112_ (_22507_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  and _68113_ (_22508_, _22015_, _22498_);
  and _68114_ (_22509_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or _68115_ (_22510_, _22509_, _22507_);
  and _68116_ (_22511_, _22019_, _22498_);
  and _68117_ (_22512_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and _68118_ (_22513_, _22022_, _22498_);
  and _68119_ (_22514_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  or _68120_ (_22515_, _22514_, _22512_);
  or _68121_ (_22516_, _22515_, _22510_);
  and _68122_ (_22517_, _21988_, _22498_);
  and _68123_ (_22518_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  and _68124_ (_22519_, _21993_, _22498_);
  and _68125_ (_22520_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or _68126_ (_22521_, _22520_, _22518_);
  and _68127_ (_22522_, _21998_, _22498_);
  and _68128_ (_22523_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and _68129_ (_22524_, _22364_, _22139_);
  and _68130_ (_22525_, _22003_, _22524_);
  and _68131_ (_22526_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  or _68132_ (_22527_, _22526_, _22523_);
  or _68133_ (_22528_, _22527_, _22521_);
  or _68134_ (_22529_, _22528_, _22516_);
  and _68135_ (_22530_, _22044_, _22498_);
  and _68136_ (_22531_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and _68137_ (_22532_, _22047_, _22498_);
  and _68138_ (_22533_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  or _68139_ (_22534_, _22533_, _22531_);
  and _68140_ (_22535_, _22498_, _22054_);
  and _68141_ (_22536_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and _68142_ (_22537_, _22498_, _22051_);
  and _68143_ (_22538_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or _68144_ (_22539_, _22538_, _22536_);
  or _68145_ (_22540_, _22539_, _22534_);
  and _68146_ (_22541_, _22498_, _22039_);
  and _68147_ (_22542_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  and _68148_ (_22543_, _22498_, _22035_);
  and _68149_ (_22544_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or _68150_ (_22545_, _22544_, _22542_);
  and _68151_ (_22546_, _22498_, _22031_);
  and _68152_ (_22547_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and _68153_ (_22548_, _22028_, _22498_);
  and _68154_ (_22549_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  or _68155_ (_22550_, _22549_, _22547_);
  or _68156_ (_22551_, _22550_, _22545_);
  or _68157_ (_22552_, _22551_, _22540_);
  or _68158_ (_22553_, _22552_, _22529_);
  and _68159_ (_22554_, _22524_, _21993_);
  and _68160_ (_22555_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and _68161_ (_22556_, _22524_, _21988_);
  and _68162_ (_22557_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  or _68163_ (_22558_, _22557_, _22555_);
  nor _68164_ (_22559_, _21983_, _21690_);
  and _68165_ (_22560_, _22559_, _21945_);
  and _68166_ (_22561_, _22003_, _22560_);
  and _68167_ (_22562_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  and _68168_ (_22563_, _22524_, _21998_);
  and _68169_ (_22564_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or _68170_ (_22565_, _22564_, _22562_);
  or _68171_ (_22566_, _22565_, _22558_);
  and _68172_ (_22567_, _22524_, _22015_);
  and _68173_ (_22568_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and _68174_ (_22569_, _22524_, _22012_);
  and _68175_ (_22570_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  or _68176_ (_22571_, _22570_, _22568_);
  and _68177_ (_22572_, _22524_, _22022_);
  and _68178_ (_22573_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  and _68179_ (_22574_, _22524_, _22019_);
  and _68180_ (_22575_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or _68181_ (_22576_, _22575_, _22573_);
  or _68182_ (_22577_, _22576_, _22571_);
  or _68183_ (_22578_, _22577_, _22566_);
  and _68184_ (_22579_, _22524_, _22044_);
  and _68185_ (_22580_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  and _68186_ (_22581_, _22524_, _22047_);
  and _68187_ (_22582_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or _68188_ (_22583_, _22582_, _22580_);
  and _68189_ (_22584_, _22524_, _22054_);
  and _68190_ (_22585_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  and _68191_ (_22586_, _22524_, _22051_);
  and _68192_ (_22587_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  or _68193_ (_22588_, _22587_, _22585_);
  or _68194_ (_22589_, _22588_, _22583_);
  and _68195_ (_22590_, _22524_, _22031_);
  and _68196_ (_22591_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  and _68197_ (_22592_, _22524_, _22028_);
  and _68198_ (_22593_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or _68199_ (_22594_, _22593_, _22591_);
  and _68200_ (_22595_, _22524_, _22035_);
  and _68201_ (_22596_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and _68202_ (_22597_, _22524_, _22039_);
  and _68203_ (_22598_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  or _68204_ (_22599_, _22598_, _22596_);
  or _68205_ (_22600_, _22599_, _22594_);
  or _68206_ (_22601_, _22600_, _22589_);
  or _68207_ (_22602_, _22601_, _22578_);
  or _68208_ (_22603_, _22602_, _22553_);
  or _68209_ (_22604_, _22603_, _22505_);
  and _68210_ (_22605_, _22047_, _22560_);
  and _68211_ (_22606_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and _68212_ (_22607_, _22044_, _22560_);
  and _68213_ (_22608_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  or _68214_ (_22609_, _22608_, _22606_);
  and _68215_ (_22610_, _22560_, _22054_);
  and _68216_ (_22611_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and _68217_ (_22612_, _22560_, _22051_);
  and _68218_ (_22613_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or _68219_ (_22614_, _22613_, _22611_);
  or _68220_ (_22615_, _22614_, _22609_);
  and _68221_ (_22616_, _22028_, _22560_);
  and _68222_ (_22617_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and _68223_ (_22618_, _22560_, _22031_);
  and _68224_ (_22619_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  or _68225_ (_22620_, _22619_, _22617_);
  and _68226_ (_22621_, _22560_, _22039_);
  and _68227_ (_22622_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  and _68228_ (_22623_, _22560_, _22035_);
  and _68229_ (_22624_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or _68230_ (_22625_, _22624_, _22622_);
  or _68231_ (_22626_, _22625_, _22620_);
  or _68232_ (_22627_, _22626_, _22615_);
  and _68233_ (_22628_, _22012_, _22560_);
  and _68234_ (_22629_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  and _68235_ (_22630_, _22015_, _22560_);
  and _68236_ (_22631_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or _68237_ (_22632_, _22631_, _22629_);
  and _68238_ (_22633_, _22019_, _22560_);
  and _68239_ (_22634_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and _68240_ (_22635_, _22560_, _22022_);
  and _68241_ (_22636_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  or _68242_ (_22637_, _22636_, _22634_);
  or _68243_ (_22638_, _22637_, _22632_);
  and _68244_ (_22639_, _21988_, _22560_);
  and _68245_ (_22640_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  and _68246_ (_22641_, _22560_, _21993_);
  and _68247_ (_22642_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or _68248_ (_22643_, _22642_, _22640_);
  and _68249_ (_22644_, _21998_, _22560_);
  and _68250_ (_22645_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and _68251_ (_22646_, _22559_, _22004_);
  and _68252_ (_22647_, _22003_, _22646_);
  and _68253_ (_22648_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  or _68254_ (_22649_, _22648_, _22645_);
  or _68255_ (_22650_, _22649_, _22643_);
  or _68256_ (_22651_, _22650_, _22638_);
  or _68257_ (_22652_, _22651_, _22627_);
  and _68258_ (_22653_, _22646_, _22028_);
  and _68259_ (_22654_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  and _68260_ (_22655_, _22646_, _22031_);
  and _68261_ (_22656_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or _68262_ (_22657_, _22656_, _22654_);
  and _68263_ (_22658_, _22646_, _22035_);
  and _68264_ (_22659_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and _68265_ (_22660_, _22646_, _22039_);
  and _68266_ (_22661_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  or _68267_ (_22662_, _22661_, _22659_);
  or _68268_ (_22663_, _22662_, _22657_);
  and _68269_ (_22664_, _22047_, _22646_);
  and _68270_ (_22665_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  and _68271_ (_22666_, _22044_, _22646_);
  and _68272_ (_22667_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or _68273_ (_22668_, _22667_, _22665_);
  and _68274_ (_22669_, _22646_, _22051_);
  and _68275_ (_22670_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and _68276_ (_22671_, _22646_, _22054_);
  and _68277_ (_22672_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or _68278_ (_22673_, _22672_, _22670_);
  or _68279_ (_22674_, _22673_, _22668_);
  or _68280_ (_22675_, _22674_, _22663_);
  and _68281_ (_22676_, _22015_, _22646_);
  and _68282_ (_22677_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and _68283_ (_22678_, _22012_, _22646_);
  and _68284_ (_22679_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  or _68285_ (_22680_, _22679_, _22677_);
  and _68286_ (_22681_, _22019_, _22646_);
  and _68287_ (_22682_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  and _68288_ (_22683_, _22646_, _22022_);
  and _68289_ (_22684_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or _68290_ (_22685_, _22684_, _22682_);
  or _68291_ (_22686_, _22685_, _22680_);
  and _68292_ (_22687_, _21988_, _22646_);
  and _68293_ (_22688_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and _68294_ (_22689_, _22646_, _21993_);
  and _68295_ (_22690_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  or _68296_ (_22691_, _22690_, _22688_);
  and _68297_ (_22692_, _22559_, _22066_);
  and _68298_ (_22693_, _22003_, _22692_);
  and _68299_ (_22694_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  and _68300_ (_22695_, _21998_, _22646_);
  and _68301_ (_22696_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or _68302_ (_22697_, _22696_, _22694_);
  or _68303_ (_22698_, _22697_, _22691_);
  or _68304_ (_22699_, _22698_, _22686_);
  or _68305_ (_22700_, _22699_, _22675_);
  or _68306_ (_22701_, _22700_, _22652_);
  and _68307_ (_22702_, _22559_, _22139_);
  and _68308_ (_22703_, _22012_, _22702_);
  and _68309_ (_22704_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and _68310_ (_22705_, _22015_, _22702_);
  and _68311_ (_22706_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or _68312_ (_22707_, _22706_, _22704_);
  and _68313_ (_22708_, _22019_, _22702_);
  and _68314_ (_22709_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _68315_ (_22710_, _22709_, _22707_);
  and _68316_ (_22711_, _21988_, _22702_);
  and _68317_ (_22712_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and _68318_ (_22713_, _21998_, _22702_);
  and _68319_ (_22714_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or _68320_ (_22715_, _22714_, _22712_);
  and _68321_ (_22716_, _22702_, _21993_);
  and _68322_ (_22717_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and _68323_ (_22718_, _22702_, _22022_);
  and _68324_ (_22719_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or _68325_ (_22720_, _22719_, _22717_);
  or _68326_ (_22721_, _22720_, _22715_);
  or _68327_ (_22722_, _22721_, _22710_);
  and _68328_ (_22723_, _22044_, _22702_);
  and _68329_ (_22724_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and _68330_ (_22725_, _22047_, _22702_);
  and _68331_ (_22726_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or _68332_ (_22727_, _22726_, _22724_);
  and _68333_ (_22728_, _22702_, _22051_);
  and _68334_ (_22729_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and _68335_ (_22730_, _22702_, _22054_);
  and _68336_ (_22731_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or _68337_ (_22732_, _22731_, _22729_);
  or _68338_ (_22733_, _22732_, _22727_);
  and _68339_ (_22734_, _22702_, _22031_);
  and _68340_ (_22735_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and _68341_ (_22736_, _22028_, _22702_);
  and _68342_ (_22737_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or _68343_ (_22738_, _22737_, _22735_);
  and _68344_ (_22739_, _22702_, _22039_);
  and _68345_ (_22740_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and _68346_ (_22741_, _22702_, _22035_);
  and _68347_ (_22742_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or _68348_ (_22743_, _22742_, _22740_);
  or _68349_ (_22744_, _22743_, _22738_);
  or _68350_ (_22745_, _22744_, _22733_);
  or _68351_ (_22746_, _22745_, _22722_);
  and _68352_ (_22747_, _22692_, _22028_);
  and _68353_ (_22748_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and _68354_ (_22749_, _22692_, _22031_);
  and _68355_ (_22750_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  or _68356_ (_22751_, _22750_, _22748_);
  and _68357_ (_22752_, _22692_, _22035_);
  and _68358_ (_22753_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  and _68359_ (_22754_, _22692_, _22039_);
  and _68360_ (_22755_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or _68361_ (_22756_, _22755_, _22753_);
  or _68362_ (_22757_, _22756_, _22751_);
  and _68363_ (_22758_, _22692_, _22044_);
  and _68364_ (_22759_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and _68365_ (_22760_, _22692_, _22047_);
  and _68366_ (_22761_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  or _68367_ (_22762_, _22761_, _22759_);
  and _68368_ (_22763_, _22692_, _22051_);
  and _68369_ (_22764_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  and _68370_ (_22765_, _22692_, _22054_);
  and _68371_ (_22766_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  or _68372_ (_22767_, _22766_, _22764_);
  or _68373_ (_22768_, _22767_, _22762_);
  or _68374_ (_22769_, _22768_, _22757_);
  and _68375_ (_22770_, _22692_, _22015_);
  and _68376_ (_22771_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  and _68377_ (_22772_, _22692_, _22012_);
  and _68378_ (_22773_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or _68379_ (_22774_, _22773_, _22771_);
  and _68380_ (_22775_, _22692_, _22022_);
  and _68381_ (_22776_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and _68382_ (_22777_, _22692_, _22019_);
  and _68383_ (_22778_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  or _68384_ (_22779_, _22778_, _22776_);
  or _68385_ (_22780_, _22779_, _22774_);
  and _68386_ (_22781_, _22003_, _22702_);
  and _68387_ (_22782_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and _68388_ (_22783_, _22692_, _21998_);
  and _68389_ (_22784_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  or _68390_ (_22785_, _22784_, _22782_);
  and _68391_ (_22786_, _21988_, _22692_);
  and _68392_ (_22787_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  and _68393_ (_22788_, _22692_, _21993_);
  and _68394_ (_22789_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or _68395_ (_22790_, _22789_, _22787_);
  or _68396_ (_22791_, _22790_, _22785_);
  or _68397_ (_22792_, _22791_, _22780_);
  or _68398_ (_22793_, _22792_, _22769_);
  or _68399_ (_22794_, _22793_, _22746_);
  or _68400_ (_22795_, _22794_, _22701_);
  or _68401_ (_22796_, _22795_, _22604_);
  or _68402_ (_22797_, _22796_, _22408_);
  nor _68403_ (_22798_, _22032_, _22029_);
  nor _68404_ (_22799_, _22040_, _22036_);
  and _68405_ (_22800_, _22799_, _22798_);
  nor _68406_ (_22801_, _22055_, _22052_);
  nor _68407_ (_22802_, _22048_, _22045_);
  and _68408_ (_22803_, _22802_, _22801_);
  and _68409_ (_22804_, _22803_, _22800_);
  nor _68410_ (_22805_, _22006_, _21999_);
  nor _68411_ (_22806_, _21994_, _21989_);
  and _68412_ (_22807_, _22806_, _22805_);
  nor _68413_ (_22808_, _22016_, _22013_);
  nor _68414_ (_22809_, _22023_, _22020_);
  and _68415_ (_22810_, _22809_, _22808_);
  and _68416_ (_22811_, _22810_, _22807_);
  and _68417_ (_22812_, _22811_, _22804_);
  nor _68418_ (_22813_, _22070_, _22061_);
  nor _68419_ (_22814_, _22068_, _22063_);
  and _68420_ (_22815_, _22814_, _22813_);
  nor _68421_ (_22816_, _22081_, _22079_);
  nor _68422_ (_22817_, _22076_, _22074_);
  and _68423_ (_22818_, _22817_, _22816_);
  and _68424_ (_22819_, _22818_, _22815_);
  nor _68425_ (_22820_, _22099_, _22097_);
  nor _68426_ (_22821_, _22104_, _22102_);
  and _68427_ (_22822_, _22821_, _22820_);
  nor _68428_ (_22823_, _22088_, _22086_);
  nor _68429_ (_22824_, _22093_, _22091_);
  and _68430_ (_22825_, _22824_, _22823_);
  and _68431_ (_22826_, _22825_, _22822_);
  and _68432_ (_22827_, _22826_, _22819_);
  and _68433_ (_22828_, _22827_, _22812_);
  nor _68434_ (_22829_, _22154_, _22152_);
  nor _68435_ (_22830_, _22149_, _22147_);
  and _68436_ (_22831_, _22830_, _22829_);
  nor _68437_ (_22832_, _22136_, _22134_);
  nor _68438_ (_22833_, _22143_, _22141_);
  and _68439_ (_22834_, _22833_, _22832_);
  and _68440_ (_22835_, _22834_, _22831_);
  nor _68441_ (_22836_, _22129_, _22127_);
  nor _68442_ (_22837_, _22124_, _22122_);
  and _68443_ (_22838_, _22837_, _22836_);
  nor _68444_ (_22839_, _22118_, _22116_);
  nor _68445_ (_22840_, _22113_, _22111_);
  and _68446_ (_22841_, _22840_, _22839_);
  and _68447_ (_22842_, _22841_, _22838_);
  and _68448_ (_22843_, _22842_, _22835_);
  nor _68449_ (_22844_, _22196_, _22204_);
  nor _68450_ (_22845_, _22202_, _22194_);
  and _68451_ (_22846_, _22845_, _22844_);
  nor _68452_ (_22847_, _22185_, _22183_);
  nor _68453_ (_22848_, _22190_, _22188_);
  and _68454_ (_22849_, _22848_, _22847_);
  and _68455_ (_22850_, _22849_, _22846_);
  nor _68456_ (_22851_, _22178_, _22176_);
  nor _68457_ (_22852_, _22173_, _22171_);
  and _68458_ (_22853_, _22852_, _22851_);
  nor _68459_ (_22854_, _22167_, _22165_);
  nor _68460_ (_22855_, _22162_, _22160_);
  and _68461_ (_22856_, _22855_, _22854_);
  and _68462_ (_22857_, _22856_, _22853_);
  and _68463_ (_22858_, _22857_, _22850_);
  and _68464_ (_22859_, _22858_, _22843_);
  and _68465_ (_22860_, _22859_, _22828_);
  nor _68466_ (_22861_, _22231_, _22229_);
  nor _68467_ (_22862_, _22225_, _22223_);
  and _68468_ (_22863_, _22862_, _22861_);
  nor _68469_ (_22864_, _22214_, _22212_);
  nor _68470_ (_22865_, _22219_, _22217_);
  and _68471_ (_22866_, _22865_, _22864_);
  and _68472_ (_22867_, _22866_, _22863_);
  nor _68473_ (_22868_, _22249_, _22247_);
  nor _68474_ (_22869_, _22254_, _22252_);
  and _68475_ (_22870_, _22869_, _22868_);
  nor _68476_ (_22871_, _22243_, _22241_);
  nor _68477_ (_22872_, _22238_, _22236_);
  and _68478_ (_22873_, _22872_, _22871_);
  and _68479_ (_22874_, _22873_, _22870_);
  and _68480_ (_22875_, _22874_, _22867_);
  nor _68481_ (_22876_, _22296_, _22302_);
  nor _68482_ (_22877_, _22300_, _22294_);
  and _68483_ (_22878_, _22877_, _22876_);
  nor _68484_ (_22879_, _22285_, _22283_);
  nor _68485_ (_22880_, _22290_, _22288_);
  and _68486_ (_22881_, _22880_, _22879_);
  and _68487_ (_22882_, _22881_, _22878_);
  nor _68488_ (_22883_, _22273_, _22271_);
  nor _68489_ (_22884_, _22278_, _22276_);
  and _68490_ (_22885_, _22884_, _22883_);
  nor _68491_ (_22886_, _22267_, _22265_);
  nor _68492_ (_22887_, _22262_, _22260_);
  and _68493_ (_22888_, _22887_, _22886_);
  and _68494_ (_22889_, _22888_, _22885_);
  and _68495_ (_22890_, _22889_, _22882_);
  and _68496_ (_22891_, _22890_, _22875_);
  nor _68497_ (_22892_, _22335_, _22333_);
  nor _68498_ (_22893_, _22340_, _22338_);
  and _68499_ (_22894_, _22893_, _22892_);
  nor _68500_ (_22895_, _22351_, _22349_);
  nor _68501_ (_22896_, _22346_, _22344_);
  and _68502_ (_22897_, _22896_, _22895_);
  and _68503_ (_22898_, _22897_, _22894_);
  nor _68504_ (_22899_, _22317_, _22314_);
  nor _68505_ (_22900_, _22311_, _22309_);
  and _68506_ (_22901_, _22900_, _22899_);
  nor _68507_ (_22902_, _22323_, _22321_);
  nor _68508_ (_22903_, _22328_, _22326_);
  and _68509_ (_22904_, _22903_, _22902_);
  and _68510_ (_22905_, _22904_, _22901_);
  and _68511_ (_22906_, _22905_, _22898_);
  nor _68512_ (_22907_, _22384_, _22382_);
  nor _68513_ (_22908_, _22389_, _22387_);
  and _68514_ (_22909_, _22908_, _22907_);
  nor _68515_ (_22910_, _22400_, _22398_);
  nor _68516_ (_22911_, _22395_, _22393_);
  and _68517_ (_22912_, _22911_, _22910_);
  and _68518_ (_22913_, _22912_, _22909_);
  nor _68519_ (_22914_, _22366_, _22362_);
  nor _68520_ (_22915_, _22359_, _22357_);
  and _68521_ (_22916_, _22915_, _22914_);
  nor _68522_ (_22917_, _22372_, _22370_);
  nor _68523_ (_22918_, _22377_, _22375_);
  and _68524_ (_22919_, _22918_, _22917_);
  and _68525_ (_22920_, _22919_, _22916_);
  and _68526_ (_22921_, _22920_, _22913_);
  and _68527_ (_22922_, _22921_, _22906_);
  and _68528_ (_22923_, _22922_, _22891_);
  and _68529_ (_22924_, _22923_, _22860_);
  nor _68530_ (_22925_, _22428_, _22420_);
  nor _68531_ (_22926_, _22422_, _22426_);
  and _68532_ (_22927_, _22926_, _22925_);
  nor _68533_ (_22928_, _22416_, _22414_);
  nor _68534_ (_22929_, _22411_, _22409_);
  and _68535_ (_22930_, _22929_, _22928_);
  and _68536_ (_22931_, _22930_, _22927_);
  nor _68537_ (_22932_, _22440_, _22438_);
  nor _68538_ (_22933_, _22435_, _22433_);
  and _68539_ (_22934_, _22933_, _22932_);
  nor _68540_ (_22935_, _22446_, _22444_);
  nor _68541_ (_22936_, _22451_, _22449_);
  and _68542_ (_22937_, _22936_, _22935_);
  and _68543_ (_22938_, _22937_, _22934_);
  and _68544_ (_22939_, _22938_, _22931_);
  nor _68545_ (_22940_, _22493_, _22491_);
  nor _68546_ (_22941_, _22499_, _22496_);
  and _68547_ (_22942_, _22941_, _22940_);
  nor _68548_ (_22943_, _22487_, _22485_);
  nor _68549_ (_22944_, _22482_, _22480_);
  and _68550_ (_22945_, _22944_, _22943_);
  and _68551_ (_22946_, _22945_, _22942_);
  nor _68552_ (_22947_, _22470_, _22468_);
  nor _68553_ (_22948_, _22475_, _22473_);
  and _68554_ (_22949_, _22948_, _22947_);
  nor _68555_ (_22950_, _22459_, _22457_);
  nor _68556_ (_22951_, _22464_, _22462_);
  and _68557_ (_22952_, _22951_, _22950_);
  and _68558_ (_22953_, _22952_, _22949_);
  and _68559_ (_22954_, _22953_, _22946_);
  and _68560_ (_22955_, _22954_, _22939_);
  nor _68561_ (_22956_, _22519_, _22517_);
  nor _68562_ (_22957_, _22525_, _22522_);
  and _68563_ (_22958_, _22957_, _22956_);
  nor _68564_ (_22959_, _22508_, _22506_);
  nor _68565_ (_22960_, _22513_, _22511_);
  and _68566_ (_22961_, _22960_, _22959_);
  and _68567_ (_22962_, _22961_, _22958_);
  nor _68568_ (_22963_, _22548_, _22546_);
  nor _68569_ (_22964_, _22543_, _22541_);
  and _68570_ (_22965_, _22964_, _22963_);
  nor _68571_ (_22966_, _22532_, _22530_);
  nor _68572_ (_22967_, _22537_, _22535_);
  and _68573_ (_22968_, _22967_, _22966_);
  and _68574_ (_22969_, _22968_, _22965_);
  and _68575_ (_22970_, _22969_, _22962_);
  nor _68576_ (_22971_, _22563_, _22554_);
  nor _68577_ (_22972_, _22556_, _22561_);
  and _68578_ (_22973_, _22972_, _22971_);
  nor _68579_ (_22974_, _22574_, _22572_);
  nor _68580_ (_22975_, _22569_, _22567_);
  and _68581_ (_22976_, _22975_, _22974_);
  and _68582_ (_22977_, _22976_, _22973_);
  nor _68583_ (_22978_, _22592_, _22590_);
  nor _68584_ (_22979_, _22597_, _22595_);
  and _68585_ (_22980_, _22979_, _22978_);
  nor _68586_ (_22981_, _22581_, _22579_);
  nor _68587_ (_22982_, _22586_, _22584_);
  and _68588_ (_22983_, _22982_, _22981_);
  and _68589_ (_22984_, _22983_, _22980_);
  and _68590_ (_22985_, _22984_, _22977_);
  and _68591_ (_22986_, _22985_, _22970_);
  and _68592_ (_22987_, _22986_, _22955_);
  nor _68593_ (_22988_, _22644_, _22641_);
  nor _68594_ (_22989_, _22647_, _22639_);
  and _68595_ (_22990_, _22989_, _22988_);
  nor _68596_ (_22991_, _22635_, _22633_);
  nor _68597_ (_22992_, _22630_, _22628_);
  and _68598_ (_22993_, _22992_, _22991_);
  and _68599_ (_22994_, _22993_, _22990_);
  nor _68600_ (_22995_, _22607_, _22605_);
  nor _68601_ (_22996_, _22612_, _22610_);
  and _68602_ (_22997_, _22996_, _22995_);
  nor _68603_ (_22998_, _22618_, _22616_);
  nor _68604_ (_22999_, _22623_, _22621_);
  and _68605_ (_23000_, _22999_, _22998_);
  and _68606_ (_23001_, _23000_, _22997_);
  and _68607_ (_23002_, _23001_, _22994_);
  nor _68608_ (_23003_, _22695_, _22689_);
  nor _68609_ (_23004_, _22687_, _22693_);
  and _68610_ (_23005_, _23004_, _23003_);
  nor _68611_ (_23006_, _22678_, _22676_);
  nor _68612_ (_23007_, _22683_, _22681_);
  and _68613_ (_23008_, _23007_, _23006_);
  and _68614_ (_23009_, _23008_, _23005_);
  nor _68615_ (_23010_, _22671_, _22669_);
  nor _68616_ (_23011_, _22666_, _22664_);
  and _68617_ (_23012_, _23011_, _23010_);
  nor _68618_ (_23013_, _22655_, _22653_);
  nor _68619_ (_23014_, _22660_, _22658_);
  and _68620_ (_23015_, _23014_, _23013_);
  and _68621_ (_23016_, _23015_, _23012_);
  and _68622_ (_23017_, _23016_, _23009_);
  and _68623_ (_23018_, _23017_, _23002_);
  nor _68624_ (_23019_, _22788_, _22786_);
  nor _68625_ (_23020_, _22783_, _22781_);
  and _68626_ (_23021_, _23020_, _23019_);
  nor _68627_ (_23022_, _22772_, _22770_);
  nor _68628_ (_23023_, _22777_, _22775_);
  and _68629_ (_23024_, _23023_, _23022_);
  and _68630_ (_23025_, _23024_, _23021_);
  nor _68631_ (_23026_, _22754_, _22752_);
  nor _68632_ (_23027_, _22749_, _22747_);
  and _68633_ (_23028_, _23027_, _23026_);
  nor _68634_ (_23029_, _22765_, _22763_);
  nor _68635_ (_23030_, _22760_, _22758_);
  and _68636_ (_23031_, _23030_, _23029_);
  and _68637_ (_23032_, _23031_, _23028_);
  and _68638_ (_23033_, _23032_, _23025_);
  nor _68639_ (_23034_, _22012_, _22015_);
  nor _68640_ (_23035_, _22019_, _21986_);
  nand _68641_ (_23036_, _23035_, _23034_);
  nand _68642_ (_23037_, _23036_, _22702_);
  nor _68643_ (_23038_, _22725_, _22723_);
  nor _68644_ (_23039_, _22730_, _22728_);
  and _68645_ (_23040_, _23039_, _23038_);
  nor _68646_ (_23041_, _22741_, _22739_);
  nor _68647_ (_23042_, _22736_, _22734_);
  and _68648_ (_23043_, _23042_, _23041_);
  and _68649_ (_23044_, _23043_, _23040_);
  and _68650_ (_23045_, _23044_, _23037_);
  and _68651_ (_23046_, _23045_, _23033_);
  and _68652_ (_23047_, _23046_, _23018_);
  and _68653_ (_23048_, _23047_, _22987_);
  and _68654_ (_23049_, _23048_, _22924_);
  and _68655_ (_23050_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or _68656_ (_23051_, _23050_, _22797_);
  and _68657_ (_23052_, _23051_, _00006_);
  or _68658_ (_23053_, _23052_, _21944_);
  and _68659_ (_00003_[6], _23053_, _38997_);
  and _68660_ (_23054_, _15589_, iram_op1[5]);
  and _68661_ (_23055_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  and _68662_ (_23056_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or _68663_ (_23057_, _23056_, _23055_);
  and _68664_ (_23058_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and _68665_ (_23059_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or _68666_ (_23060_, _23059_, _23058_);
  or _68667_ (_23061_, _23060_, _23057_);
  and _68668_ (_23062_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  and _68669_ (_23063_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or _68670_ (_23064_, _23063_, _23062_);
  and _68671_ (_23065_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and _68672_ (_23066_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  or _68673_ (_23067_, _23066_, _23065_);
  or _68674_ (_23068_, _23067_, _23064_);
  or _68675_ (_23069_, _23068_, _23061_);
  and _68676_ (_23070_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and _68677_ (_23071_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  or _68678_ (_23072_, _23071_, _23070_);
  and _68679_ (_23073_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  and _68680_ (_23074_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or _68681_ (_23075_, _23074_, _23073_);
  or _68682_ (_23076_, _23075_, _23072_);
  and _68683_ (_23077_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and _68684_ (_23078_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  or _68685_ (_23079_, _23078_, _23077_);
  and _68686_ (_23080_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and _68687_ (_23081_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or _68688_ (_23082_, _23081_, _23080_);
  or _68689_ (_23083_, _23082_, _23079_);
  or _68690_ (_23084_, _23083_, _23076_);
  or _68691_ (_23085_, _23084_, _23069_);
  and _68692_ (_23086_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and _68693_ (_23087_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  or _68694_ (_23088_, _23087_, _23086_);
  and _68695_ (_23089_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  and _68696_ (_23090_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or _68697_ (_23091_, _23090_, _23089_);
  or _68698_ (_23092_, _23091_, _23088_);
  and _68699_ (_23093_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and _68700_ (_23094_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or _68701_ (_23095_, _23094_, _23093_);
  and _68702_ (_23096_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  and _68703_ (_23097_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or _68704_ (_23098_, _23097_, _23096_);
  or _68705_ (_23099_, _23098_, _23095_);
  or _68706_ (_23100_, _23099_, _23092_);
  and _68707_ (_23101_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  and _68708_ (_23102_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  or _68709_ (_23103_, _23102_, _23101_);
  and _68710_ (_23104_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  and _68711_ (_23105_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or _68712_ (_23106_, _23105_, _23104_);
  or _68713_ (_23107_, _23106_, _23103_);
  and _68714_ (_23108_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  and _68715_ (_23109_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or _68716_ (_23110_, _23109_, _23108_);
  and _68717_ (_23111_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and _68718_ (_23112_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or _68719_ (_23113_, _23112_, _23111_);
  or _68720_ (_23114_, _23113_, _23110_);
  or _68721_ (_23115_, _23114_, _23107_);
  or _68722_ (_23116_, _23115_, _23100_);
  or _68723_ (_23117_, _23116_, _23085_);
  and _68724_ (_23118_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and _68725_ (_23119_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  or _68726_ (_23120_, _23119_, _23118_);
  and _68727_ (_23121_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  and _68728_ (_23122_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or _68729_ (_23123_, _23122_, _23121_);
  or _68730_ (_23124_, _23123_, _23120_);
  and _68731_ (_23125_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and _68732_ (_23126_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  or _68733_ (_23127_, _23126_, _23125_);
  and _68734_ (_23128_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and _68735_ (_23129_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or _68736_ (_23130_, _23129_, _23128_);
  or _68737_ (_23131_, _23130_, _23127_);
  or _68738_ (_23132_, _23131_, _23124_);
  and _68739_ (_23133_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and _68740_ (_23134_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  or _68741_ (_23135_, _23134_, _23133_);
  and _68742_ (_23136_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  and _68743_ (_23137_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or _68744_ (_23138_, _23137_, _23136_);
  or _68745_ (_23139_, _23138_, _23135_);
  and _68746_ (_23140_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  and _68747_ (_23141_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or _68748_ (_23142_, _23141_, _23140_);
  and _68749_ (_23143_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and _68750_ (_23144_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or _68751_ (_23145_, _23144_, _23143_);
  or _68752_ (_23146_, _23145_, _23142_);
  or _68753_ (_23147_, _23146_, _23139_);
  or _68754_ (_23148_, _23147_, _23132_);
  and _68755_ (_23149_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  and _68756_ (_23150_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or _68757_ (_23151_, _23150_, _23149_);
  and _68758_ (_23152_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and _68759_ (_23153_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or _68760_ (_23154_, _23153_, _23152_);
  or _68761_ (_23155_, _23154_, _23151_);
  and _68762_ (_23156_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  and _68763_ (_23157_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or _68764_ (_23158_, _23157_, _23156_);
  and _68765_ (_23159_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and _68766_ (_23160_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or _68767_ (_23161_, _23160_, _23159_);
  or _68768_ (_23162_, _23161_, _23158_);
  or _68769_ (_23163_, _23162_, _23155_);
  and _68770_ (_23164_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and _68771_ (_23165_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or _68772_ (_23166_, _23165_, _23164_);
  and _68773_ (_23167_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  and _68774_ (_23168_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or _68775_ (_23169_, _23168_, _23167_);
  or _68776_ (_23170_, _23169_, _23166_);
  and _68777_ (_23171_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and _68778_ (_23172_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or _68779_ (_23173_, _23172_, _23171_);
  and _68780_ (_23174_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  and _68781_ (_23175_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or _68782_ (_23176_, _23175_, _23174_);
  or _68783_ (_23177_, _23176_, _23173_);
  or _68784_ (_23178_, _23177_, _23170_);
  or _68785_ (_23179_, _23178_, _23163_);
  or _68786_ (_23180_, _23179_, _23148_);
  or _68787_ (_23181_, _23180_, _23117_);
  and _68788_ (_23182_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and _68789_ (_23183_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or _68790_ (_23184_, _23183_, _23182_);
  and _68791_ (_23185_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  and _68792_ (_23186_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or _68793_ (_23187_, _23186_, _23185_);
  or _68794_ (_23188_, _23187_, _23184_);
  and _68795_ (_23189_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and _68796_ (_23190_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  or _68797_ (_23191_, _23190_, _23189_);
  and _68798_ (_23192_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and _68799_ (_23193_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or _68800_ (_23194_, _23193_, _23192_);
  or _68801_ (_23195_, _23194_, _23191_);
  or _68802_ (_23196_, _23195_, _23188_);
  and _68803_ (_23197_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  and _68804_ (_23198_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or _68805_ (_23199_, _23198_, _23197_);
  and _68806_ (_23200_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and _68807_ (_23201_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  or _68808_ (_23202_, _23201_, _23200_);
  or _68809_ (_23203_, _23202_, _23199_);
  and _68810_ (_23204_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and _68811_ (_23205_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or _68812_ (_23206_, _23205_, _23204_);
  and _68813_ (_23207_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  and _68814_ (_23208_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or _68815_ (_23209_, _23208_, _23207_);
  or _68816_ (_23210_, _23209_, _23206_);
  or _68817_ (_23211_, _23210_, _23203_);
  or _68818_ (_23212_, _23211_, _23196_);
  and _68819_ (_23213_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  and _68820_ (_23214_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or _68821_ (_23215_, _23214_, _23213_);
  and _68822_ (_23216_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and _68823_ (_23217_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  or _68824_ (_23218_, _23217_, _23216_);
  or _68825_ (_23219_, _23218_, _23215_);
  and _68826_ (_23220_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  and _68827_ (_23221_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or _68828_ (_23222_, _23221_, _23220_);
  and _68829_ (_23223_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and _68830_ (_23224_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or _68831_ (_23225_, _23224_, _23223_);
  or _68832_ (_23226_, _23225_, _23222_);
  or _68833_ (_23227_, _23226_, _23219_);
  and _68834_ (_23228_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and _68835_ (_23229_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  or _68836_ (_23230_, _23229_, _23228_);
  and _68837_ (_23231_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  and _68838_ (_23232_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or _68839_ (_23233_, _23232_, _23231_);
  or _68840_ (_23234_, _23233_, _23230_);
  and _68841_ (_23235_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and _68842_ (_23236_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  or _68843_ (_23237_, _23236_, _23235_);
  and _68844_ (_23238_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  and _68845_ (_23239_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or _68846_ (_23240_, _23239_, _23238_);
  or _68847_ (_23241_, _23240_, _23237_);
  or _68848_ (_23242_, _23241_, _23234_);
  or _68849_ (_23243_, _23242_, _23227_);
  or _68850_ (_23244_, _23243_, _23212_);
  and _68851_ (_23245_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  and _68852_ (_23246_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or _68853_ (_23247_, _23246_, _23245_);
  and _68854_ (_23248_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and _68855_ (_23249_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  or _68856_ (_23250_, _23249_, _23248_);
  or _68857_ (_23251_, _23250_, _23247_);
  and _68858_ (_23252_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and _68859_ (_23253_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  or _68860_ (_23254_, _23253_, _23252_);
  and _68861_ (_23255_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  and _68862_ (_23256_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or _68863_ (_23257_, _23256_, _23255_);
  or _68864_ (_23258_, _23257_, _23254_);
  or _68865_ (_23259_, _23258_, _23251_);
  and _68866_ (_23260_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and _68867_ (_23261_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  or _68868_ (_23262_, _23261_, _23260_);
  and _68869_ (_23263_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  and _68870_ (_23264_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or _68871_ (_23265_, _23264_, _23263_);
  or _68872_ (_23266_, _23265_, _23262_);
  and _68873_ (_23267_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and _68874_ (_23268_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  or _68875_ (_23269_, _23268_, _23267_);
  and _68876_ (_23270_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and _68877_ (_23271_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or _68878_ (_23272_, _23271_, _23270_);
  or _68879_ (_23273_, _23272_, _23269_);
  or _68880_ (_23274_, _23273_, _23266_);
  or _68881_ (_23275_, _23274_, _23259_);
  and _68882_ (_23276_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  and _68883_ (_23277_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or _68884_ (_23278_, _23277_, _23276_);
  and _68885_ (_23279_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  and _68886_ (_23280_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  or _68887_ (_23281_, _23280_, _23279_);
  or _68888_ (_23282_, _23281_, _23278_);
  and _68889_ (_23283_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and _68890_ (_23284_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  or _68891_ (_23285_, _23284_, _23283_);
  and _68892_ (_23286_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  and _68893_ (_23287_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or _68894_ (_23288_, _23287_, _23286_);
  or _68895_ (_23289_, _23288_, _23285_);
  or _68896_ (_23290_, _23289_, _23282_);
  and _68897_ (_23291_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and _68898_ (_23292_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  or _68899_ (_23293_, _23292_, _23291_);
  and _68900_ (_23294_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  and _68901_ (_23295_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or _68902_ (_23296_, _23295_, _23294_);
  or _68903_ (_23297_, _23296_, _23293_);
  and _68904_ (_23298_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and _68905_ (_23299_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  or _68906_ (_23300_, _23299_, _23298_);
  and _68907_ (_23301_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  and _68908_ (_23302_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or _68909_ (_23303_, _23302_, _23301_);
  or _68910_ (_23304_, _23303_, _23300_);
  or _68911_ (_23305_, _23304_, _23297_);
  or _68912_ (_23306_, _23305_, _23290_);
  or _68913_ (_23307_, _23306_, _23275_);
  or _68914_ (_23308_, _23307_, _23244_);
  or _68915_ (_23309_, _23308_, _23181_);
  and _68916_ (_23310_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  and _68917_ (_23311_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or _68918_ (_23312_, _23311_, _23310_);
  and _68919_ (_23313_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and _68920_ (_23314_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  or _68921_ (_23315_, _23314_, _23313_);
  or _68922_ (_23316_, _23315_, _23312_);
  and _68923_ (_23317_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  and _68924_ (_23318_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or _68925_ (_23319_, _23318_, _23317_);
  and _68926_ (_23320_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and _68927_ (_23321_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  or _68928_ (_23322_, _23321_, _23320_);
  or _68929_ (_23323_, _23322_, _23319_);
  or _68930_ (_23324_, _23323_, _23316_);
  and _68931_ (_23325_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and _68932_ (_23326_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  or _68933_ (_23327_, _23326_, _23325_);
  and _68934_ (_23328_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and _68935_ (_23329_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or _68936_ (_23330_, _23329_, _23328_);
  or _68937_ (_23331_, _23330_, _23327_);
  and _68938_ (_23332_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and _68939_ (_23333_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  or _68940_ (_23334_, _23333_, _23332_);
  and _68941_ (_23335_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  and _68942_ (_23336_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or _68943_ (_23337_, _23336_, _23335_);
  or _68944_ (_23338_, _23337_, _23334_);
  or _68945_ (_23339_, _23338_, _23331_);
  or _68946_ (_23340_, _23339_, _23324_);
  and _68947_ (_23341_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  and _68948_ (_23342_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or _68949_ (_23343_, _23342_, _23341_);
  and _68950_ (_23344_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and _68951_ (_23345_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or _68952_ (_23346_, _23345_, _23344_);
  or _68953_ (_23347_, _23346_, _23343_);
  and _68954_ (_23348_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  and _68955_ (_23349_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or _68956_ (_23350_, _23349_, _23348_);
  and _68957_ (_23351_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and _68958_ (_23352_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or _68959_ (_23353_, _23352_, _23351_);
  or _68960_ (_23354_, _23353_, _23350_);
  or _68961_ (_23355_, _23354_, _23347_);
  and _68962_ (_23356_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and _68963_ (_23357_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  or _68964_ (_23358_, _23357_, _23356_);
  and _68965_ (_23359_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  and _68966_ (_23360_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or _68967_ (_23361_, _23360_, _23359_);
  or _68968_ (_23362_, _23361_, _23358_);
  and _68969_ (_23363_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and _68970_ (_23364_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  or _68971_ (_23365_, _23364_, _23363_);
  and _68972_ (_23366_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  and _68973_ (_23367_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or _68974_ (_23368_, _23367_, _23366_);
  or _68975_ (_23369_, _23368_, _23365_);
  or _68976_ (_23370_, _23369_, _23362_);
  or _68977_ (_23371_, _23370_, _23355_);
  or _68978_ (_23372_, _23371_, _23340_);
  and _68979_ (_23373_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  and _68980_ (_23374_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or _68981_ (_23375_, _23374_, _23373_);
  and _68982_ (_23376_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and _68983_ (_23377_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or _68984_ (_23378_, _23377_, _23376_);
  or _68985_ (_23379_, _23378_, _23375_);
  and _68986_ (_23380_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  and _68987_ (_23381_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or _68988_ (_23382_, _23381_, _23380_);
  and _68989_ (_23383_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and _68990_ (_23384_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or _68991_ (_23385_, _23384_, _23383_);
  or _68992_ (_23386_, _23385_, _23382_);
  or _68993_ (_23387_, _23386_, _23379_);
  and _68994_ (_23388_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and _68995_ (_23389_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  or _68996_ (_23390_, _23389_, _23388_);
  and _68997_ (_23391_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  and _68998_ (_23392_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or _68999_ (_23393_, _23392_, _23391_);
  or _69000_ (_23394_, _23393_, _23390_);
  and _69001_ (_23395_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and _69002_ (_23396_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or _69003_ (_23397_, _23396_, _23395_);
  and _69004_ (_23398_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  and _69005_ (_23399_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or _69006_ (_23400_, _23399_, _23398_);
  or _69007_ (_23401_, _23400_, _23397_);
  or _69008_ (_23402_, _23401_, _23394_);
  or _69009_ (_23403_, _23402_, _23387_);
  and _69010_ (_23404_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  and _69011_ (_23405_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or _69012_ (_23406_, _23405_, _23404_);
  and _69013_ (_23407_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and _69014_ (_23408_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  or _69015_ (_23409_, _23408_, _23407_);
  or _69016_ (_23410_, _23409_, _23406_);
  and _69017_ (_23411_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  and _69018_ (_23412_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or _69019_ (_23413_, _23412_, _23411_);
  and _69020_ (_23414_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  and _69021_ (_23415_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or _69022_ (_23416_, _23415_, _23414_);
  or _69023_ (_23417_, _23416_, _23413_);
  or _69024_ (_23418_, _23417_, _23410_);
  and _69025_ (_23419_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and _69026_ (_23420_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or _69027_ (_23421_, _23420_, _23419_);
  and _69028_ (_23422_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  and _69029_ (_23423_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or _69030_ (_23424_, _23423_, _23422_);
  or _69031_ (_23425_, _23424_, _23421_);
  and _69032_ (_23426_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and _69033_ (_23427_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  or _69034_ (_23428_, _23427_, _23426_);
  and _69035_ (_23429_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  and _69036_ (_23430_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or _69037_ (_23431_, _23430_, _23429_);
  or _69038_ (_23432_, _23431_, _23428_);
  or _69039_ (_23433_, _23432_, _23425_);
  or _69040_ (_23434_, _23433_, _23418_);
  or _69041_ (_23435_, _23434_, _23403_);
  or _69042_ (_23436_, _23435_, _23372_);
  and _69043_ (_23437_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  and _69044_ (_23438_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or _69045_ (_23439_, _23438_, _23437_);
  and _69046_ (_23440_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and _69047_ (_23441_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or _69048_ (_23442_, _23441_, _23440_);
  or _69049_ (_23443_, _23442_, _23439_);
  and _69050_ (_23444_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  and _69051_ (_23445_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or _69052_ (_23446_, _23445_, _23444_);
  and _69053_ (_23447_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and _69054_ (_23448_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  or _69055_ (_23449_, _23448_, _23447_);
  or _69056_ (_23450_, _23449_, _23446_);
  or _69057_ (_23451_, _23450_, _23443_);
  and _69058_ (_23452_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and _69059_ (_23453_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  or _69060_ (_23454_, _23453_, _23452_);
  and _69061_ (_23455_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  and _69062_ (_23456_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or _69063_ (_23457_, _23456_, _23455_);
  or _69064_ (_23458_, _23457_, _23454_);
  and _69065_ (_23459_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and _69066_ (_23460_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  or _69067_ (_23461_, _23460_, _23459_);
  and _69068_ (_23462_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  and _69069_ (_23463_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  or _69070_ (_23464_, _23463_, _23462_);
  or _69071_ (_23465_, _23464_, _23461_);
  or _69072_ (_23466_, _23465_, _23458_);
  or _69073_ (_23467_, _23466_, _23451_);
  and _69074_ (_23468_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and _69075_ (_23469_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  or _69076_ (_23470_, _23469_, _23468_);
  and _69077_ (_23471_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  and _69078_ (_23472_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or _69079_ (_23473_, _23472_, _23471_);
  or _69080_ (_23474_, _23473_, _23470_);
  and _69081_ (_23475_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and _69082_ (_23476_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  or _69083_ (_23477_, _23476_, _23475_);
  and _69084_ (_23478_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  and _69085_ (_23479_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or _69086_ (_23480_, _23479_, _23478_);
  or _69087_ (_23481_, _23480_, _23477_);
  or _69088_ (_23482_, _23481_, _23474_);
  and _69089_ (_23483_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  and _69090_ (_23484_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or _69091_ (_23485_, _23484_, _23483_);
  and _69092_ (_23486_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and _69093_ (_23487_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or _69094_ (_23488_, _23487_, _23486_);
  or _69095_ (_23489_, _23488_, _23485_);
  and _69096_ (_23490_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  and _69097_ (_23491_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or _69098_ (_23492_, _23491_, _23490_);
  and _69099_ (_23493_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  and _69100_ (_23494_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  or _69101_ (_23495_, _23494_, _23493_);
  or _69102_ (_23496_, _23495_, _23492_);
  or _69103_ (_23497_, _23496_, _23489_);
  or _69104_ (_23498_, _23497_, _23482_);
  or _69105_ (_23499_, _23498_, _23467_);
  and _69106_ (_23500_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and _69107_ (_23501_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  or _69108_ (_23502_, _23501_, _23500_);
  and _69109_ (_23503_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  and _69110_ (_23504_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  or _69111_ (_23505_, _23504_, _23503_);
  or _69112_ (_23506_, _23505_, _23502_);
  and _69113_ (_23507_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and _69114_ (_23508_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  or _69115_ (_23509_, _23508_, _23507_);
  and _69116_ (_23510_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  and _69117_ (_23511_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or _69118_ (_23512_, _23511_, _23510_);
  or _69119_ (_23513_, _23512_, _23509_);
  or _69120_ (_23514_, _23513_, _23506_);
  and _69121_ (_23515_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  and _69122_ (_23516_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or _69123_ (_23517_, _23516_, _23515_);
  and _69124_ (_23518_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and _69125_ (_23519_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  or _69126_ (_23520_, _23519_, _23518_);
  or _69127_ (_23521_, _23520_, _23517_);
  and _69128_ (_23522_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  and _69129_ (_23523_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or _69130_ (_23524_, _23523_, _23522_);
  and _69131_ (_23525_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and _69132_ (_23526_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or _69133_ (_23527_, _23526_, _23525_);
  or _69134_ (_23528_, _23527_, _23524_);
  or _69135_ (_23529_, _23528_, _23521_);
  or _69136_ (_23530_, _23529_, _23514_);
  and _69137_ (_23531_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and _69138_ (_23532_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or _69139_ (_23533_, _23532_, _23531_);
  and _69140_ (_23534_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and _69141_ (_23535_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or _69142_ (_23536_, _23535_, _23534_);
  or _69143_ (_23537_, _23536_, _23533_);
  and _69144_ (_23538_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and _69145_ (_23539_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or _69146_ (_23540_, _23539_, _23538_);
  and _69147_ (_23541_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and _69148_ (_23542_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or _69149_ (_23543_, _23542_, _23541_);
  or _69150_ (_23544_, _23543_, _23540_);
  or _69151_ (_23545_, _23544_, _23537_);
  and _69152_ (_23546_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and _69153_ (_23547_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _69154_ (_23548_, _23547_, _23546_);
  and _69155_ (_23549_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and _69156_ (_23550_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or _69157_ (_23551_, _23550_, _23549_);
  or _69158_ (_23552_, _23551_, _23548_);
  and _69159_ (_23553_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and _69160_ (_23554_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and _69161_ (_23555_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or _69162_ (_23556_, _23555_, _23554_);
  or _69163_ (_23557_, _23556_, _23553_);
  or _69164_ (_23558_, _23557_, _23552_);
  or _69165_ (_23559_, _23558_, _23545_);
  or _69166_ (_23560_, _23559_, _23530_);
  or _69167_ (_23561_, _23560_, _23499_);
  or _69168_ (_23562_, _23561_, _23436_);
  or _69169_ (_23563_, _23562_, _23309_);
  and _69170_ (_23564_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or _69171_ (_23565_, _23564_, _23563_);
  and _69172_ (_23566_, _23565_, _00006_);
  or _69173_ (_23567_, _23566_, _23054_);
  and _69174_ (_00003_[5], _23567_, _38997_);
  and _69175_ (_23568_, _15589_, iram_op1[4]);
  and _69176_ (_23569_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  and _69177_ (_23570_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or _69178_ (_23571_, _23570_, _23569_);
  and _69179_ (_23572_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and _69180_ (_23573_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  or _69181_ (_23574_, _23573_, _23572_);
  or _69182_ (_23575_, _23574_, _23571_);
  and _69183_ (_23576_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  and _69184_ (_23577_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or _69185_ (_23578_, _23577_, _23576_);
  and _69186_ (_23579_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and _69187_ (_23580_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  or _69188_ (_23581_, _23580_, _23579_);
  or _69189_ (_23582_, _23581_, _23578_);
  or _69190_ (_23583_, _23582_, _23575_);
  and _69191_ (_23584_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and _69192_ (_23585_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  or _69193_ (_23586_, _23585_, _23584_);
  and _69194_ (_23587_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  and _69195_ (_23588_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or _69196_ (_23589_, _23588_, _23587_);
  or _69197_ (_23590_, _23589_, _23586_);
  and _69198_ (_23591_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and _69199_ (_23592_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  or _69200_ (_23593_, _23592_, _23591_);
  and _69201_ (_23594_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  and _69202_ (_23595_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  or _69203_ (_23596_, _23595_, _23594_);
  or _69204_ (_23597_, _23596_, _23593_);
  or _69205_ (_23598_, _23597_, _23590_);
  or _69206_ (_23599_, _23598_, _23583_);
  and _69207_ (_23600_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  and _69208_ (_23601_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or _69209_ (_23602_, _23601_, _23600_);
  and _69210_ (_23603_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and _69211_ (_23604_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  or _69212_ (_23605_, _23604_, _23603_);
  or _69213_ (_23606_, _23605_, _23602_);
  and _69214_ (_23607_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  and _69215_ (_23608_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or _69216_ (_23609_, _23608_, _23607_);
  and _69217_ (_23610_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and _69218_ (_23611_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or _69219_ (_23612_, _23611_, _23610_);
  or _69220_ (_23613_, _23612_, _23609_);
  or _69221_ (_23614_, _23613_, _23606_);
  and _69222_ (_23615_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and _69223_ (_23616_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  or _69224_ (_23617_, _23616_, _23615_);
  and _69225_ (_23618_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  and _69226_ (_23619_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or _69227_ (_23620_, _23619_, _23618_);
  or _69228_ (_23621_, _23620_, _23617_);
  and _69229_ (_23622_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and _69230_ (_23623_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  or _69231_ (_23624_, _23623_, _23622_);
  and _69232_ (_23625_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  and _69233_ (_23626_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or _69234_ (_23627_, _23626_, _23625_);
  or _69235_ (_23628_, _23627_, _23624_);
  or _69236_ (_23629_, _23628_, _23621_);
  or _69237_ (_23630_, _23629_, _23614_);
  or _69238_ (_23631_, _23630_, _23599_);
  and _69239_ (_23632_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and _69240_ (_23633_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  or _69241_ (_23634_, _23633_, _23632_);
  and _69242_ (_23635_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  and _69243_ (_23636_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or _69244_ (_23637_, _23636_, _23635_);
  or _69245_ (_23638_, _23637_, _23634_);
  and _69246_ (_23639_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and _69247_ (_23640_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  or _69248_ (_23641_, _23640_, _23639_);
  and _69249_ (_23642_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  and _69250_ (_23643_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or _69251_ (_23644_, _23643_, _23642_);
  or _69252_ (_23645_, _23644_, _23641_);
  or _69253_ (_23646_, _23645_, _23638_);
  and _69254_ (_23647_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  and _69255_ (_23648_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or _69256_ (_23649_, _23648_, _23647_);
  and _69257_ (_23650_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  and _69258_ (_23651_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  or _69259_ (_23652_, _23651_, _23650_);
  or _69260_ (_23653_, _23652_, _23649_);
  and _69261_ (_23654_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and _69262_ (_23655_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  or _69263_ (_23656_, _23655_, _23654_);
  and _69264_ (_23657_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  and _69265_ (_23658_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or _69266_ (_23659_, _23658_, _23657_);
  or _69267_ (_23660_, _23659_, _23656_);
  or _69268_ (_23661_, _23660_, _23653_);
  or _69269_ (_23662_, _23661_, _23646_);
  and _69270_ (_23663_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and _69271_ (_23664_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  or _69272_ (_23665_, _23664_, _23663_);
  and _69273_ (_23666_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  and _69274_ (_23667_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or _69275_ (_23668_, _23667_, _23666_);
  or _69276_ (_23669_, _23668_, _23665_);
  and _69277_ (_23670_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and _69278_ (_23671_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  or _69279_ (_23672_, _23671_, _23670_);
  and _69280_ (_23673_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  and _69281_ (_23674_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  or _69282_ (_23675_, _23674_, _23673_);
  or _69283_ (_23676_, _23675_, _23672_);
  or _69284_ (_23677_, _23676_, _23669_);
  and _69285_ (_23678_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  and _69286_ (_23679_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or _69287_ (_23680_, _23679_, _23678_);
  and _69288_ (_23681_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and _69289_ (_23682_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  or _69290_ (_23683_, _23682_, _23681_);
  or _69291_ (_23684_, _23683_, _23680_);
  and _69292_ (_23685_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  and _69293_ (_23686_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or _69294_ (_23687_, _23686_, _23685_);
  and _69295_ (_23688_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and _69296_ (_23689_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  or _69297_ (_23690_, _23689_, _23688_);
  or _69298_ (_23691_, _23690_, _23687_);
  or _69299_ (_23692_, _23691_, _23684_);
  or _69300_ (_23693_, _23692_, _23677_);
  or _69301_ (_23694_, _23693_, _23662_);
  or _69302_ (_23695_, _23694_, _23631_);
  and _69303_ (_23696_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and _69304_ (_23697_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  or _69305_ (_23698_, _23697_, _23696_);
  and _69306_ (_23699_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  and _69307_ (_23700_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or _69308_ (_23701_, _23700_, _23699_);
  or _69309_ (_23702_, _23701_, _23698_);
  and _69310_ (_23703_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and _69311_ (_23704_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  or _69312_ (_23705_, _23704_, _23703_);
  and _69313_ (_23706_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  and _69314_ (_23707_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  or _69315_ (_23708_, _23707_, _23706_);
  or _69316_ (_23709_, _23708_, _23705_);
  or _69317_ (_23710_, _23709_, _23702_);
  and _69318_ (_23711_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  and _69319_ (_23712_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or _69320_ (_23713_, _23712_, _23711_);
  and _69321_ (_23714_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and _69322_ (_23715_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  or _69323_ (_23716_, _23715_, _23714_);
  or _69324_ (_23717_, _23716_, _23713_);
  and _69325_ (_23718_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  and _69326_ (_23719_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or _69327_ (_23720_, _23719_, _23718_);
  and _69328_ (_23721_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and _69329_ (_23722_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  or _69330_ (_23723_, _23722_, _23721_);
  or _69331_ (_23724_, _23723_, _23720_);
  or _69332_ (_23725_, _23724_, _23717_);
  or _69333_ (_23726_, _23725_, _23710_);
  and _69334_ (_23727_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  and _69335_ (_23728_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or _69336_ (_23729_, _23728_, _23727_);
  and _69337_ (_23730_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and _69338_ (_23731_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  or _69339_ (_23732_, _23731_, _23730_);
  or _69340_ (_23733_, _23732_, _23729_);
  and _69341_ (_23734_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  and _69342_ (_23735_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or _69343_ (_23736_, _23735_, _23734_);
  and _69344_ (_23737_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  and _69345_ (_23738_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  or _69346_ (_23739_, _23738_, _23737_);
  or _69347_ (_23740_, _23739_, _23736_);
  or _69348_ (_23741_, _23740_, _23733_);
  and _69349_ (_23742_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  and _69350_ (_23743_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or _69351_ (_23744_, _23743_, _23742_);
  and _69352_ (_23745_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and _69353_ (_23746_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  or _69354_ (_23747_, _23746_, _23745_);
  or _69355_ (_23748_, _23747_, _23744_);
  and _69356_ (_23749_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and _69357_ (_23750_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  or _69358_ (_23751_, _23750_, _23749_);
  and _69359_ (_23752_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  and _69360_ (_23753_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or _69361_ (_23754_, _23753_, _23752_);
  or _69362_ (_23755_, _23754_, _23751_);
  or _69363_ (_23756_, _23755_, _23748_);
  or _69364_ (_23757_, _23756_, _23741_);
  or _69365_ (_23758_, _23757_, _23726_);
  and _69366_ (_23759_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  and _69367_ (_23760_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or _69368_ (_23761_, _23760_, _23759_);
  and _69369_ (_23762_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and _69370_ (_23763_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  or _69371_ (_23764_, _23763_, _23762_);
  or _69372_ (_23765_, _23764_, _23761_);
  and _69373_ (_23766_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  and _69374_ (_23767_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or _69375_ (_23768_, _23767_, _23766_);
  and _69376_ (_23769_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and _69377_ (_23770_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  or _69378_ (_23771_, _23770_, _23769_);
  or _69379_ (_23772_, _23771_, _23768_);
  or _69380_ (_23773_, _23772_, _23765_);
  and _69381_ (_23774_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and _69382_ (_23775_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  or _69383_ (_23776_, _23775_, _23774_);
  and _69384_ (_23777_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  and _69385_ (_23778_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or _69386_ (_23779_, _23778_, _23777_);
  or _69387_ (_23780_, _23779_, _23776_);
  and _69388_ (_23781_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and _69389_ (_23782_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  or _69390_ (_23783_, _23782_, _23781_);
  and _69391_ (_23784_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and _69392_ (_23785_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or _69393_ (_23786_, _23785_, _23784_);
  or _69394_ (_23787_, _23786_, _23783_);
  or _69395_ (_23788_, _23787_, _23780_);
  or _69396_ (_23789_, _23788_, _23773_);
  and _69397_ (_23790_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  and _69398_ (_23791_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or _69399_ (_23792_, _23791_, _23790_);
  and _69400_ (_23793_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  and _69401_ (_23794_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  or _69402_ (_23795_, _23794_, _23793_);
  or _69403_ (_23796_, _23795_, _23792_);
  and _69404_ (_23797_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  and _69405_ (_23798_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or _69406_ (_23799_, _23798_, _23797_);
  and _69407_ (_23800_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and _69408_ (_23801_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  or _69409_ (_23802_, _23801_, _23800_);
  or _69410_ (_23803_, _23802_, _23799_);
  or _69411_ (_23804_, _23803_, _23796_);
  and _69412_ (_23805_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and _69413_ (_23806_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  or _69414_ (_23807_, _23806_, _23805_);
  and _69415_ (_23808_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  and _69416_ (_23809_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or _69417_ (_23810_, _23809_, _23808_);
  or _69418_ (_23811_, _23810_, _23807_);
  and _69419_ (_23812_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and _69420_ (_23813_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  or _69421_ (_23814_, _23813_, _23812_);
  and _69422_ (_23815_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  and _69423_ (_23816_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or _69424_ (_23817_, _23816_, _23815_);
  or _69425_ (_23818_, _23817_, _23814_);
  or _69426_ (_23819_, _23818_, _23811_);
  or _69427_ (_23820_, _23819_, _23804_);
  or _69428_ (_23821_, _23820_, _23789_);
  or _69429_ (_23822_, _23821_, _23758_);
  or _69430_ (_23823_, _23822_, _23695_);
  and _69431_ (_23824_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  and _69432_ (_23825_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or _69433_ (_23826_, _23825_, _23824_);
  and _69434_ (_23827_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and _69435_ (_23828_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  or _69436_ (_23829_, _23828_, _23827_);
  or _69437_ (_23830_, _23829_, _23826_);
  and _69438_ (_23831_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  and _69439_ (_23832_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or _69440_ (_23833_, _23832_, _23831_);
  and _69441_ (_23834_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and _69442_ (_23835_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  or _69443_ (_23836_, _23835_, _23834_);
  or _69444_ (_23837_, _23836_, _23833_);
  or _69445_ (_23838_, _23837_, _23830_);
  and _69446_ (_23839_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and _69447_ (_23840_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  or _69448_ (_23841_, _23840_, _23839_);
  and _69449_ (_23842_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and _69450_ (_23843_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or _69451_ (_23844_, _23843_, _23842_);
  or _69452_ (_23845_, _23844_, _23841_);
  and _69453_ (_23846_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and _69454_ (_23847_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  or _69455_ (_23848_, _23847_, _23846_);
  and _69456_ (_23849_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  and _69457_ (_23850_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or _69458_ (_23851_, _23850_, _23849_);
  or _69459_ (_23852_, _23851_, _23848_);
  or _69460_ (_23853_, _23852_, _23845_);
  or _69461_ (_23854_, _23853_, _23838_);
  and _69462_ (_23855_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  and _69463_ (_23856_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or _69464_ (_23857_, _23856_, _23855_);
  and _69465_ (_23858_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and _69466_ (_23859_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  or _69467_ (_23860_, _23859_, _23858_);
  or _69468_ (_23861_, _23860_, _23857_);
  and _69469_ (_23862_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  and _69470_ (_23863_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or _69471_ (_23864_, _23863_, _23862_);
  and _69472_ (_23865_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and _69473_ (_23866_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or _69474_ (_23867_, _23866_, _23865_);
  or _69475_ (_23868_, _23867_, _23864_);
  or _69476_ (_23869_, _23868_, _23861_);
  and _69477_ (_23870_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and _69478_ (_23871_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  or _69479_ (_23872_, _23871_, _23870_);
  and _69480_ (_23873_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  and _69481_ (_23874_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or _69482_ (_23875_, _23874_, _23873_);
  or _69483_ (_23876_, _23875_, _23872_);
  and _69484_ (_23877_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and _69485_ (_23878_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  or _69486_ (_23879_, _23878_, _23877_);
  and _69487_ (_23880_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  and _69488_ (_23881_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or _69489_ (_23882_, _23881_, _23880_);
  or _69490_ (_23883_, _23882_, _23879_);
  or _69491_ (_23884_, _23883_, _23876_);
  or _69492_ (_23885_, _23884_, _23869_);
  or _69493_ (_23886_, _23885_, _23854_);
  and _69494_ (_23887_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and _69495_ (_23888_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  or _69496_ (_23889_, _23888_, _23887_);
  and _69497_ (_23890_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and _69498_ (_23891_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or _69499_ (_23892_, _23891_, _23890_);
  or _69500_ (_23893_, _23892_, _23889_);
  and _69501_ (_23894_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and _69502_ (_23895_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  or _69503_ (_23896_, _23895_, _23894_);
  and _69504_ (_23897_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  and _69505_ (_23898_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or _69506_ (_23899_, _23898_, _23897_);
  or _69507_ (_23900_, _23899_, _23896_);
  or _69508_ (_23901_, _23900_, _23893_);
  and _69509_ (_23902_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  and _69510_ (_23903_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or _69511_ (_23904_, _23903_, _23902_);
  and _69512_ (_23905_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and _69513_ (_23906_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  or _69514_ (_23907_, _23906_, _23905_);
  or _69515_ (_23908_, _23907_, _23904_);
  and _69516_ (_23909_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  and _69517_ (_23910_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or _69518_ (_23911_, _23910_, _23909_);
  and _69519_ (_23912_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and _69520_ (_23913_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or _69521_ (_23914_, _23913_, _23912_);
  or _69522_ (_23915_, _23914_, _23911_);
  or _69523_ (_23916_, _23915_, _23908_);
  or _69524_ (_23917_, _23916_, _23901_);
  and _69525_ (_23918_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and _69526_ (_23919_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or _69527_ (_23920_, _23919_, _23918_);
  and _69528_ (_23921_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  and _69529_ (_23922_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or _69530_ (_23923_, _23922_, _23921_);
  or _69531_ (_23924_, _23923_, _23920_);
  and _69532_ (_23925_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  and _69533_ (_23926_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or _69534_ (_23927_, _23926_, _23925_);
  and _69535_ (_23928_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and _69536_ (_23929_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or _69537_ (_23930_, _23929_, _23928_);
  or _69538_ (_23931_, _23930_, _23927_);
  or _69539_ (_23932_, _23931_, _23924_);
  and _69540_ (_23933_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  and _69541_ (_23934_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or _69542_ (_23935_, _23934_, _23933_);
  and _69543_ (_23936_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  and _69544_ (_23937_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or _69545_ (_23938_, _23937_, _23936_);
  or _69546_ (_23939_, _23938_, _23935_);
  and _69547_ (_23940_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  and _69548_ (_23941_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or _69549_ (_23942_, _23941_, _23940_);
  and _69550_ (_23943_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and _69551_ (_23944_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or _69552_ (_23945_, _23944_, _23943_);
  or _69553_ (_23946_, _23945_, _23942_);
  or _69554_ (_23947_, _23946_, _23939_);
  or _69555_ (_23948_, _23947_, _23932_);
  or _69556_ (_23949_, _23948_, _23917_);
  or _69557_ (_23950_, _23949_, _23886_);
  and _69558_ (_23951_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  and _69559_ (_23952_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or _69560_ (_23953_, _23952_, _23951_);
  and _69561_ (_23954_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and _69562_ (_23955_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  or _69563_ (_23956_, _23955_, _23954_);
  or _69564_ (_23957_, _23956_, _23953_);
  and _69565_ (_23958_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  and _69566_ (_23959_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or _69567_ (_23960_, _23959_, _23958_);
  and _69568_ (_23961_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and _69569_ (_23962_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or _69570_ (_23963_, _23962_, _23961_);
  or _69571_ (_23964_, _23963_, _23960_);
  or _69572_ (_23965_, _23964_, _23957_);
  and _69573_ (_23966_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and _69574_ (_23967_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  or _69575_ (_23968_, _23967_, _23966_);
  and _69576_ (_23969_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  and _69577_ (_23970_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or _69578_ (_23971_, _23970_, _23969_);
  or _69579_ (_23972_, _23971_, _23968_);
  and _69580_ (_23973_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and _69581_ (_23974_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  or _69582_ (_23975_, _23974_, _23973_);
  and _69583_ (_23976_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  and _69584_ (_23977_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or _69585_ (_23978_, _23977_, _23976_);
  or _69586_ (_23979_, _23978_, _23975_);
  or _69587_ (_23980_, _23979_, _23972_);
  or _69588_ (_23981_, _23980_, _23965_);
  and _69589_ (_23982_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and _69590_ (_23983_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  or _69591_ (_23984_, _23983_, _23982_);
  and _69592_ (_23985_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  and _69593_ (_23986_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or _69594_ (_23987_, _23986_, _23985_);
  or _69595_ (_23988_, _23987_, _23984_);
  and _69596_ (_23989_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and _69597_ (_23990_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  or _69598_ (_23991_, _23990_, _23989_);
  and _69599_ (_23992_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  and _69600_ (_23993_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  or _69601_ (_23994_, _23993_, _23992_);
  or _69602_ (_23995_, _23994_, _23991_);
  or _69603_ (_23996_, _23995_, _23988_);
  and _69604_ (_23997_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and _69605_ (_23998_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  or _69606_ (_23999_, _23998_, _23997_);
  and _69607_ (_24000_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  and _69608_ (_24001_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or _69609_ (_24002_, _24001_, _24000_);
  or _69610_ (_24003_, _24002_, _23999_);
  and _69611_ (_24004_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and _69612_ (_24005_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  or _69613_ (_24006_, _24005_, _24004_);
  and _69614_ (_24007_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  and _69615_ (_24008_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or _69616_ (_24009_, _24008_, _24007_);
  or _69617_ (_24010_, _24009_, _24006_);
  or _69618_ (_24011_, _24010_, _24003_);
  or _69619_ (_24012_, _24011_, _23996_);
  or _69620_ (_24013_, _24012_, _23981_);
  and _69621_ (_24014_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and _69622_ (_24015_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  or _69623_ (_24016_, _24015_, _24014_);
  and _69624_ (_24017_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  and _69625_ (_24018_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or _69626_ (_24019_, _24018_, _24017_);
  or _69627_ (_24020_, _24019_, _24016_);
  and _69628_ (_24021_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and _69629_ (_24022_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  or _69630_ (_24023_, _24022_, _24021_);
  and _69631_ (_24024_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and _69632_ (_24025_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or _69633_ (_24026_, _24025_, _24024_);
  or _69634_ (_24027_, _24026_, _24023_);
  or _69635_ (_24028_, _24027_, _24020_);
  and _69636_ (_24029_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  and _69637_ (_24030_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or _69638_ (_24031_, _24030_, _24029_);
  and _69639_ (_24032_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and _69640_ (_24033_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or _69641_ (_24034_, _24033_, _24032_);
  or _69642_ (_24035_, _24034_, _24031_);
  and _69643_ (_24036_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  and _69644_ (_24037_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or _69645_ (_24038_, _24037_, _24036_);
  and _69646_ (_24039_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and _69647_ (_24040_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  or _69648_ (_24041_, _24040_, _24039_);
  or _69649_ (_24042_, _24041_, _24038_);
  or _69650_ (_24043_, _24042_, _24035_);
  or _69651_ (_24044_, _24043_, _24028_);
  and _69652_ (_24045_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and _69653_ (_24046_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and _69654_ (_24047_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or _69655_ (_24048_, _24047_, _24046_);
  or _69656_ (_24049_, _24048_, _24045_);
  and _69657_ (_24050_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and _69658_ (_24051_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or _69659_ (_24052_, _24051_, _24050_);
  and _69660_ (_24053_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and _69661_ (_24054_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _69662_ (_24055_, _24054_, _24053_);
  or _69663_ (_24056_, _24055_, _24052_);
  or _69664_ (_24057_, _24056_, _24049_);
  and _69665_ (_24058_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and _69666_ (_24059_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _69667_ (_24060_, _24059_, _24058_);
  and _69668_ (_24061_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and _69669_ (_24062_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or _69670_ (_24063_, _24062_, _24061_);
  or _69671_ (_24064_, _24063_, _24060_);
  and _69672_ (_24065_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and _69673_ (_24066_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _69674_ (_24067_, _24066_, _24065_);
  and _69675_ (_24068_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and _69676_ (_24069_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or _69677_ (_24070_, _24069_, _24068_);
  or _69678_ (_24071_, _24070_, _24067_);
  or _69679_ (_24072_, _24071_, _24064_);
  or _69680_ (_24073_, _24072_, _24057_);
  or _69681_ (_24074_, _24073_, _24044_);
  or _69682_ (_24075_, _24074_, _24013_);
  or _69683_ (_24076_, _24075_, _23950_);
  or _69684_ (_24077_, _24076_, _23823_);
  and _69685_ (_24078_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or _69686_ (_24079_, _24078_, _24077_);
  and _69687_ (_24080_, _24079_, _00006_);
  or _69688_ (_24081_, _24080_, _23568_);
  and _69689_ (_00003_[4], _24081_, _38997_);
  and _69690_ (_24082_, _15589_, iram_op1[3]);
  and _69691_ (_24083_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and _69692_ (_24084_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  or _69693_ (_24085_, _24084_, _24083_);
  and _69694_ (_24086_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  and _69695_ (_24087_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or _69696_ (_24088_, _24087_, _24086_);
  or _69697_ (_24089_, _24088_, _24085_);
  and _69698_ (_24090_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and _69699_ (_24091_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  or _69700_ (_24092_, _24091_, _24090_);
  and _69701_ (_24093_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and _69702_ (_24094_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or _69703_ (_24095_, _24094_, _24093_);
  or _69704_ (_24096_, _24095_, _24092_);
  or _69705_ (_24097_, _24096_, _24089_);
  and _69706_ (_24098_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  and _69707_ (_24099_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or _69708_ (_24100_, _24099_, _24098_);
  and _69709_ (_24101_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and _69710_ (_24102_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  or _69711_ (_24103_, _24102_, _24101_);
  or _69712_ (_24104_, _24103_, _24100_);
  and _69713_ (_24105_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  and _69714_ (_24106_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or _69715_ (_24107_, _24106_, _24105_);
  and _69716_ (_24108_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and _69717_ (_24109_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  or _69718_ (_24110_, _24109_, _24108_);
  or _69719_ (_24111_, _24110_, _24107_);
  or _69720_ (_24112_, _24111_, _24104_);
  or _69721_ (_24113_, _24112_, _24097_);
  and _69722_ (_24114_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  and _69723_ (_24115_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or _69724_ (_24116_, _24115_, _24114_);
  and _69725_ (_24117_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  and _69726_ (_24118_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  or _69727_ (_24119_, _24118_, _24117_);
  or _69728_ (_24120_, _24119_, _24116_);
  and _69729_ (_24121_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  and _69730_ (_24122_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or _69731_ (_24123_, _24122_, _24121_);
  and _69732_ (_24124_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and _69733_ (_24125_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  or _69734_ (_24126_, _24125_, _24124_);
  or _69735_ (_24127_, _24126_, _24123_);
  or _69736_ (_24128_, _24127_, _24120_);
  and _69737_ (_24129_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and _69738_ (_24130_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  or _69739_ (_24131_, _24130_, _24129_);
  and _69740_ (_24132_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  and _69741_ (_24133_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or _69742_ (_24134_, _24133_, _24132_);
  or _69743_ (_24135_, _24134_, _24131_);
  and _69744_ (_24136_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and _69745_ (_24137_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  or _69746_ (_24138_, _24137_, _24136_);
  and _69747_ (_24139_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  and _69748_ (_24140_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or _69749_ (_24141_, _24140_, _24139_);
  or _69750_ (_24142_, _24141_, _24138_);
  or _69751_ (_24143_, _24142_, _24135_);
  or _69752_ (_24144_, _24143_, _24128_);
  or _69753_ (_24145_, _24144_, _24113_);
  and _69754_ (_24146_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and _69755_ (_24147_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  or _69756_ (_24148_, _24147_, _24146_);
  and _69757_ (_24149_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  and _69758_ (_24150_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or _69759_ (_24151_, _24150_, _24149_);
  or _69760_ (_24152_, _24151_, _24148_);
  and _69761_ (_24153_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and _69762_ (_24154_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  or _69763_ (_24155_, _24154_, _24153_);
  and _69764_ (_24156_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  and _69765_ (_24157_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  or _69766_ (_24158_, _24157_, _24156_);
  or _69767_ (_24159_, _24158_, _24155_);
  or _69768_ (_24160_, _24159_, _24152_);
  and _69769_ (_24161_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and _69770_ (_24162_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  or _69771_ (_24163_, _24162_, _24161_);
  and _69772_ (_24164_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  and _69773_ (_24165_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or _69774_ (_24166_, _24165_, _24164_);
  or _69775_ (_24167_, _24166_, _24163_);
  and _69776_ (_24168_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  and _69777_ (_24169_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or _69778_ (_24170_, _24169_, _24168_);
  and _69779_ (_24171_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and _69780_ (_24172_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  or _69781_ (_24173_, _24172_, _24171_);
  or _69782_ (_24174_, _24173_, _24170_);
  or _69783_ (_24175_, _24174_, _24167_);
  or _69784_ (_24176_, _24175_, _24160_);
  and _69785_ (_24177_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and _69786_ (_24178_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  or _69787_ (_24179_, _24178_, _24177_);
  and _69788_ (_24180_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  and _69789_ (_24181_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or _69790_ (_24182_, _24181_, _24180_);
  or _69791_ (_24183_, _24182_, _24179_);
  and _69792_ (_24184_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and _69793_ (_24185_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  or _69794_ (_24186_, _24185_, _24184_);
  and _69795_ (_24187_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  and _69796_ (_24188_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or _69797_ (_24189_, _24188_, _24187_);
  or _69798_ (_24190_, _24189_, _24186_);
  or _69799_ (_24191_, _24190_, _24183_);
  and _69800_ (_24192_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  and _69801_ (_24193_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or _69802_ (_24194_, _24193_, _24192_);
  and _69803_ (_24195_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and _69804_ (_24196_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or _69805_ (_24197_, _24196_, _24195_);
  or _69806_ (_24198_, _24197_, _24194_);
  and _69807_ (_24199_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  and _69808_ (_24200_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or _69809_ (_24201_, _24200_, _24199_);
  and _69810_ (_24202_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and _69811_ (_24203_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  or _69812_ (_24204_, _24203_, _24202_);
  or _69813_ (_24205_, _24204_, _24201_);
  or _69814_ (_24206_, _24205_, _24198_);
  or _69815_ (_24207_, _24206_, _24191_);
  or _69816_ (_24208_, _24207_, _24176_);
  or _69817_ (_24209_, _24208_, _24145_);
  and _69818_ (_24210_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and _69819_ (_24211_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  or _69820_ (_24212_, _24211_, _24210_);
  and _69821_ (_24213_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  and _69822_ (_24214_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or _69823_ (_24215_, _24214_, _24213_);
  or _69824_ (_24216_, _24215_, _24212_);
  and _69825_ (_24217_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and _69826_ (_24218_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  or _69827_ (_24219_, _24218_, _24217_);
  and _69828_ (_24220_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and _69829_ (_24221_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or _69830_ (_24222_, _24221_, _24220_);
  or _69831_ (_24223_, _24222_, _24219_);
  or _69832_ (_24224_, _24223_, _24216_);
  and _69833_ (_24225_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  and _69834_ (_24226_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or _69835_ (_24227_, _24226_, _24225_);
  and _69836_ (_24228_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and _69837_ (_24229_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  or _69838_ (_24230_, _24229_, _24228_);
  or _69839_ (_24231_, _24230_, _24227_);
  and _69840_ (_24232_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and _69841_ (_24233_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  or _69842_ (_24234_, _24233_, _24232_);
  and _69843_ (_24235_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  and _69844_ (_24236_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or _69845_ (_24237_, _24236_, _24235_);
  or _69846_ (_24238_, _24237_, _24234_);
  or _69847_ (_24239_, _24238_, _24231_);
  or _69848_ (_24240_, _24239_, _24224_);
  and _69849_ (_24241_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  and _69850_ (_24242_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or _69851_ (_24243_, _24242_, _24241_);
  and _69852_ (_24244_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and _69853_ (_24245_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  or _69854_ (_24246_, _24245_, _24244_);
  or _69855_ (_24247_, _24246_, _24243_);
  and _69856_ (_24248_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  and _69857_ (_24249_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or _69858_ (_24250_, _24249_, _24248_);
  and _69859_ (_24251_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and _69860_ (_24252_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or _69861_ (_24253_, _24252_, _24251_);
  or _69862_ (_24254_, _24253_, _24250_);
  or _69863_ (_24255_, _24254_, _24247_);
  and _69864_ (_24256_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and _69865_ (_24257_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  or _69866_ (_24258_, _24257_, _24256_);
  and _69867_ (_24259_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  and _69868_ (_24260_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or _69869_ (_24261_, _24260_, _24259_);
  or _69870_ (_24262_, _24261_, _24258_);
  and _69871_ (_24263_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and _69872_ (_24264_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  or _69873_ (_24265_, _24264_, _24263_);
  and _69874_ (_24266_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  and _69875_ (_24267_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or _69876_ (_24268_, _24267_, _24266_);
  or _69877_ (_24269_, _24268_, _24265_);
  or _69878_ (_24270_, _24269_, _24262_);
  or _69879_ (_24271_, _24270_, _24255_);
  or _69880_ (_24272_, _24271_, _24240_);
  and _69881_ (_24273_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and _69882_ (_24274_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or _69883_ (_24275_, _24274_, _24273_);
  and _69884_ (_24276_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and _69885_ (_24277_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  or _69886_ (_24278_, _24277_, _24276_);
  or _69887_ (_24279_, _24278_, _24275_);
  and _69888_ (_24280_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and _69889_ (_24281_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  or _69890_ (_24282_, _24281_, _24280_);
  and _69891_ (_24283_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  and _69892_ (_24284_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or _69893_ (_24285_, _24284_, _24283_);
  or _69894_ (_24286_, _24285_, _24282_);
  or _69895_ (_24287_, _24286_, _24279_);
  and _69896_ (_24288_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  and _69897_ (_24289_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or _69898_ (_24290_, _24289_, _24288_);
  and _69899_ (_24291_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and _69900_ (_24292_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  or _69901_ (_24293_, _24292_, _24291_);
  or _69902_ (_24294_, _24293_, _24290_);
  and _69903_ (_24295_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  and _69904_ (_24296_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or _69905_ (_24297_, _24296_, _24295_);
  and _69906_ (_24298_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and _69907_ (_24299_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  or _69908_ (_24300_, _24299_, _24298_);
  or _69909_ (_24301_, _24300_, _24297_);
  or _69910_ (_24302_, _24301_, _24294_);
  or _69911_ (_24303_, _24302_, _24287_);
  and _69912_ (_24304_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  and _69913_ (_24305_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or _69914_ (_24306_, _24305_, _24304_);
  and _69915_ (_24307_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and _69916_ (_24308_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or _69917_ (_24309_, _24308_, _24307_);
  or _69918_ (_24310_, _24309_, _24306_);
  and _69919_ (_24311_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  and _69920_ (_24312_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or _69921_ (_24313_, _24312_, _24311_);
  and _69922_ (_24314_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and _69923_ (_24315_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  or _69924_ (_24316_, _24315_, _24314_);
  or _69925_ (_24317_, _24316_, _24313_);
  or _69926_ (_24318_, _24317_, _24310_);
  and _69927_ (_24319_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and _69928_ (_24320_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  or _69929_ (_24321_, _24320_, _24319_);
  and _69930_ (_24322_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  and _69931_ (_24323_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or _69932_ (_24324_, _24323_, _24322_);
  or _69933_ (_24325_, _24324_, _24321_);
  and _69934_ (_24326_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and _69935_ (_24327_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  or _69936_ (_24328_, _24327_, _24326_);
  and _69937_ (_24329_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  and _69938_ (_24330_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or _69939_ (_24331_, _24330_, _24329_);
  or _69940_ (_24332_, _24331_, _24328_);
  or _69941_ (_24333_, _24332_, _24325_);
  or _69942_ (_24334_, _24333_, _24318_);
  or _69943_ (_24335_, _24334_, _24303_);
  or _69944_ (_24336_, _24335_, _24272_);
  or _69945_ (_24337_, _24336_, _24209_);
  and _69946_ (_24338_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  and _69947_ (_24339_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or _69948_ (_24340_, _24339_, _24338_);
  and _69949_ (_24341_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and _69950_ (_24342_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  or _69951_ (_24343_, _24342_, _24341_);
  or _69952_ (_24344_, _24343_, _24340_);
  and _69953_ (_24345_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  and _69954_ (_24346_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or _69955_ (_24347_, _24346_, _24345_);
  and _69956_ (_24348_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and _69957_ (_24349_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  or _69958_ (_24350_, _24349_, _24348_);
  or _69959_ (_24351_, _24350_, _24347_);
  or _69960_ (_24352_, _24351_, _24344_);
  and _69961_ (_24353_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and _69962_ (_24354_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  or _69963_ (_24355_, _24354_, _24353_);
  and _69964_ (_24356_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and _69965_ (_24357_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or _69966_ (_24358_, _24357_, _24356_);
  or _69967_ (_24359_, _24358_, _24355_);
  and _69968_ (_24360_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and _69969_ (_24361_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  or _69970_ (_24362_, _24361_, _24360_);
  and _69971_ (_24363_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  and _69972_ (_24364_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or _69973_ (_24365_, _24364_, _24363_);
  or _69974_ (_24366_, _24365_, _24362_);
  or _69975_ (_24367_, _24366_, _24359_);
  or _69976_ (_24368_, _24367_, _24352_);
  and _69977_ (_24369_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  and _69978_ (_24370_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or _69979_ (_24371_, _24370_, _24369_);
  and _69980_ (_24372_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and _69981_ (_24373_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  or _69982_ (_24374_, _24373_, _24372_);
  or _69983_ (_24375_, _24374_, _24371_);
  and _69984_ (_24376_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  and _69985_ (_24377_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or _69986_ (_24378_, _24377_, _24376_);
  and _69987_ (_24379_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  and _69988_ (_24380_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  or _69989_ (_24381_, _24380_, _24379_);
  or _69990_ (_24382_, _24381_, _24378_);
  or _69991_ (_24383_, _24382_, _24375_);
  and _69992_ (_24384_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and _69993_ (_24385_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  or _69994_ (_24386_, _24385_, _24384_);
  and _69995_ (_24387_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  and _69996_ (_24388_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or _69997_ (_24389_, _24388_, _24387_);
  or _69998_ (_24390_, _24389_, _24386_);
  and _69999_ (_24391_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and _70000_ (_24392_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  or _70001_ (_24393_, _24392_, _24391_);
  and _70002_ (_24394_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  and _70003_ (_24395_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or _70004_ (_24396_, _24395_, _24394_);
  or _70005_ (_24397_, _24396_, _24393_);
  or _70006_ (_24398_, _24397_, _24390_);
  or _70007_ (_24399_, _24398_, _24383_);
  or _70008_ (_24400_, _24399_, _24368_);
  and _70009_ (_24401_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  and _70010_ (_24402_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  or _70011_ (_24403_, _24402_, _24401_);
  and _70012_ (_24404_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and _70013_ (_24405_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  or _70014_ (_24406_, _24405_, _24404_);
  or _70015_ (_24407_, _24406_, _24403_);
  and _70016_ (_24408_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and _70017_ (_24409_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  or _70018_ (_24410_, _24409_, _24408_);
  and _70019_ (_24411_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  and _70020_ (_24412_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or _70021_ (_24413_, _24412_, _24411_);
  or _70022_ (_24414_, _24413_, _24410_);
  or _70023_ (_24415_, _24414_, _24407_);
  and _70024_ (_24416_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  and _70025_ (_24417_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or _70026_ (_24418_, _24417_, _24416_);
  and _70027_ (_24419_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and _70028_ (_24420_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  or _70029_ (_24421_, _24420_, _24419_);
  or _70030_ (_24422_, _24421_, _24418_);
  and _70031_ (_24423_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  and _70032_ (_24424_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or _70033_ (_24425_, _24424_, _24423_);
  and _70034_ (_24426_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and _70035_ (_24427_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or _70036_ (_24428_, _24427_, _24426_);
  or _70037_ (_24429_, _24428_, _24425_);
  or _70038_ (_24430_, _24429_, _24422_);
  or _70039_ (_24431_, _24430_, _24415_);
  and _70040_ (_24432_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and _70041_ (_24433_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or _70042_ (_24434_, _24433_, _24432_);
  and _70043_ (_24435_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  and _70044_ (_24436_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or _70045_ (_24437_, _24436_, _24435_);
  or _70046_ (_24438_, _24437_, _24434_);
  and _70047_ (_24439_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and _70048_ (_24440_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or _70049_ (_24441_, _24440_, _24439_);
  and _70050_ (_24442_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  and _70051_ (_24443_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or _70052_ (_24444_, _24443_, _24442_);
  or _70053_ (_24445_, _24444_, _24441_);
  or _70054_ (_24446_, _24445_, _24438_);
  and _70055_ (_24447_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and _70056_ (_24448_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or _70057_ (_24449_, _24448_, _24447_);
  and _70058_ (_24450_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  and _70059_ (_24451_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or _70060_ (_24452_, _24451_, _24450_);
  or _70061_ (_24453_, _24452_, _24449_);
  and _70062_ (_24454_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  and _70063_ (_24455_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or _70064_ (_24456_, _24455_, _24454_);
  and _70065_ (_24457_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  and _70066_ (_24458_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or _70067_ (_24459_, _24458_, _24457_);
  or _70068_ (_24460_, _24459_, _24456_);
  or _70069_ (_24461_, _24460_, _24453_);
  or _70070_ (_24462_, _24461_, _24446_);
  or _70071_ (_24463_, _24462_, _24431_);
  or _70072_ (_24464_, _24463_, _24400_);
  and _70073_ (_24465_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  and _70074_ (_24466_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or _70075_ (_24467_, _24466_, _24465_);
  and _70076_ (_24468_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and _70077_ (_24469_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  or _70078_ (_24470_, _24469_, _24468_);
  or _70079_ (_24471_, _24470_, _24467_);
  and _70080_ (_24472_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  and _70081_ (_24473_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or _70082_ (_24474_, _24473_, _24472_);
  and _70083_ (_24475_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and _70084_ (_24476_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  or _70085_ (_24477_, _24476_, _24475_);
  or _70086_ (_24478_, _24477_, _24474_);
  or _70087_ (_24479_, _24478_, _24471_);
  and _70088_ (_24480_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and _70089_ (_24481_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  or _70090_ (_24482_, _24481_, _24480_);
  and _70091_ (_24483_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  and _70092_ (_24484_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or _70093_ (_24485_, _24484_, _24483_);
  or _70094_ (_24486_, _24485_, _24482_);
  and _70095_ (_24487_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and _70096_ (_24488_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  or _70097_ (_24489_, _24488_, _24487_);
  and _70098_ (_24490_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  and _70099_ (_24491_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  or _70100_ (_24492_, _24491_, _24490_);
  or _70101_ (_24493_, _24492_, _24489_);
  or _70102_ (_24494_, _24493_, _24486_);
  or _70103_ (_24495_, _24494_, _24479_);
  and _70104_ (_24496_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  and _70105_ (_24497_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or _70106_ (_24498_, _24497_, _24496_);
  and _70107_ (_24499_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and _70108_ (_24500_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  or _70109_ (_24501_, _24500_, _24499_);
  or _70110_ (_24502_, _24501_, _24498_);
  and _70111_ (_24503_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  and _70112_ (_24504_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or _70113_ (_24505_, _24504_, _24503_);
  and _70114_ (_24506_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and _70115_ (_24507_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or _70116_ (_24508_, _24507_, _24506_);
  or _70117_ (_24509_, _24508_, _24505_);
  or _70118_ (_24510_, _24509_, _24502_);
  and _70119_ (_24511_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and _70120_ (_24512_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  or _70121_ (_24513_, _24512_, _24511_);
  and _70122_ (_24514_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  and _70123_ (_24515_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or _70124_ (_24516_, _24515_, _24514_);
  or _70125_ (_24517_, _24516_, _24513_);
  and _70126_ (_24518_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and _70127_ (_24519_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  or _70128_ (_24520_, _24519_, _24518_);
  and _70129_ (_24521_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  and _70130_ (_24522_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or _70131_ (_24523_, _24522_, _24521_);
  or _70132_ (_24524_, _24523_, _24520_);
  or _70133_ (_24525_, _24524_, _24517_);
  or _70134_ (_24526_, _24525_, _24510_);
  or _70135_ (_24527_, _24526_, _24495_);
  and _70136_ (_24528_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  and _70137_ (_24529_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or _70138_ (_24530_, _24529_, _24528_);
  and _70139_ (_24531_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and _70140_ (_24532_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or _70141_ (_24533_, _24532_, _24531_);
  or _70142_ (_24534_, _24533_, _24530_);
  and _70143_ (_24535_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  and _70144_ (_24536_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or _70145_ (_24537_, _24536_, _24535_);
  and _70146_ (_24538_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and _70147_ (_24539_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  or _70148_ (_24540_, _24539_, _24538_);
  or _70149_ (_24541_, _24540_, _24537_);
  or _70150_ (_24542_, _24541_, _24534_);
  and _70151_ (_24543_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and _70152_ (_24544_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  or _70153_ (_24545_, _24544_, _24543_);
  and _70154_ (_24546_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  and _70155_ (_24547_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  or _70156_ (_24548_, _24547_, _24546_);
  or _70157_ (_24549_, _24548_, _24545_);
  and _70158_ (_24550_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and _70159_ (_24551_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  or _70160_ (_24552_, _24551_, _24550_);
  and _70161_ (_24553_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  and _70162_ (_24554_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or _70163_ (_24555_, _24554_, _24553_);
  or _70164_ (_24556_, _24555_, _24552_);
  or _70165_ (_24557_, _24556_, _24549_);
  or _70166_ (_24558_, _24557_, _24542_);
  and _70167_ (_24559_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and _70168_ (_24560_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or _70169_ (_24561_, _24560_, _24559_);
  and _70170_ (_24562_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and _70171_ (_24563_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or _70172_ (_24564_, _24563_, _24562_);
  or _70173_ (_24565_, _24564_, _24561_);
  and _70174_ (_24566_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and _70175_ (_24567_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or _70176_ (_24568_, _24567_, _24566_);
  and _70177_ (_24569_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and _70178_ (_24570_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or _70179_ (_24571_, _24570_, _24569_);
  or _70180_ (_24572_, _24571_, _24568_);
  or _70181_ (_24573_, _24572_, _24565_);
  and _70182_ (_24574_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and _70183_ (_24575_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or _70184_ (_24576_, _24575_, _24574_);
  and _70185_ (_24577_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and _70186_ (_24578_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _70187_ (_24579_, _24578_, _24577_);
  or _70188_ (_24580_, _24579_, _24576_);
  and _70189_ (_24581_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and _70190_ (_24582_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and _70191_ (_24583_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _70192_ (_24584_, _24583_, _24582_);
  or _70193_ (_24585_, _24584_, _24581_);
  or _70194_ (_24586_, _24585_, _24580_);
  or _70195_ (_24587_, _24586_, _24573_);
  or _70196_ (_24588_, _24587_, _24558_);
  or _70197_ (_24589_, _24588_, _24527_);
  or _70198_ (_24590_, _24589_, _24464_);
  or _70199_ (_24591_, _24590_, _24337_);
  and _70200_ (_24592_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or _70201_ (_24593_, _24592_, _24591_);
  and _70202_ (_24594_, _24593_, _00006_);
  or _70203_ (_24595_, _24594_, _24082_);
  and _70204_ (_00003_[3], _24595_, _38997_);
  and _70205_ (_24596_, _15589_, iram_op1[2]);
  and _70206_ (_24597_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and _70207_ (_24598_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  or _70208_ (_24599_, _24598_, _24597_);
  and _70209_ (_24600_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and _70210_ (_24601_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or _70211_ (_24602_, _24601_, _24600_);
  or _70212_ (_24603_, _24602_, _24599_);
  and _70213_ (_24604_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and _70214_ (_24605_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  or _70215_ (_24606_, _24605_, _24604_);
  and _70216_ (_24607_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  and _70217_ (_24608_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or _70218_ (_24609_, _24608_, _24607_);
  or _70219_ (_24610_, _24609_, _24606_);
  or _70220_ (_24611_, _24610_, _24603_);
  and _70221_ (_24612_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  and _70222_ (_24613_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or _70223_ (_24614_, _24613_, _24612_);
  and _70224_ (_24615_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and _70225_ (_24616_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  or _70226_ (_24617_, _24616_, _24615_);
  or _70227_ (_24618_, _24617_, _24614_);
  and _70228_ (_24619_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  and _70229_ (_24620_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or _70230_ (_24621_, _24620_, _24619_);
  and _70231_ (_24622_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and _70232_ (_24623_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  or _70233_ (_24624_, _24623_, _24622_);
  or _70234_ (_24625_, _24624_, _24621_);
  or _70235_ (_24626_, _24625_, _24618_);
  or _70236_ (_24627_, _24626_, _24611_);
  and _70237_ (_24628_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  and _70238_ (_24629_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or _70239_ (_24630_, _24629_, _24628_);
  and _70240_ (_24631_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and _70241_ (_24632_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or _70242_ (_24633_, _24632_, _24631_);
  or _70243_ (_24634_, _24633_, _24630_);
  and _70244_ (_24635_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  and _70245_ (_24636_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or _70246_ (_24637_, _24636_, _24635_);
  and _70247_ (_24638_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and _70248_ (_24639_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  or _70249_ (_24640_, _24639_, _24638_);
  or _70250_ (_24641_, _24640_, _24637_);
  or _70251_ (_24642_, _24641_, _24634_);
  and _70252_ (_24643_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and _70253_ (_24644_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  or _70254_ (_24645_, _24644_, _24643_);
  and _70255_ (_24646_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  and _70256_ (_24647_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or _70257_ (_24648_, _24647_, _24646_);
  or _70258_ (_24649_, _24648_, _24645_);
  and _70259_ (_24650_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and _70260_ (_24651_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  or _70261_ (_24652_, _24651_, _24650_);
  and _70262_ (_24653_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  and _70263_ (_24654_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or _70264_ (_24655_, _24654_, _24653_);
  or _70265_ (_24656_, _24655_, _24652_);
  or _70266_ (_24657_, _24656_, _24649_);
  or _70267_ (_24658_, _24657_, _24642_);
  or _70268_ (_24659_, _24658_, _24627_);
  and _70269_ (_24660_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and _70270_ (_24661_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  or _70271_ (_24662_, _24661_, _24660_);
  and _70272_ (_24663_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  and _70273_ (_24664_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or _70274_ (_24665_, _24664_, _24663_);
  or _70275_ (_24666_, _24665_, _24662_);
  and _70276_ (_24667_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and _70277_ (_24668_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  or _70278_ (_24669_, _24668_, _24667_);
  and _70279_ (_24670_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  and _70280_ (_24671_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  or _70281_ (_24672_, _24671_, _24670_);
  or _70282_ (_24673_, _24672_, _24669_);
  or _70283_ (_24674_, _24673_, _24666_);
  and _70284_ (_24675_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  and _70285_ (_24676_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or _70286_ (_24677_, _24676_, _24675_);
  and _70287_ (_24678_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and _70288_ (_24679_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  or _70289_ (_24680_, _24679_, _24678_);
  or _70290_ (_24681_, _24680_, _24677_);
  and _70291_ (_24682_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  and _70292_ (_24683_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or _70293_ (_24684_, _24683_, _24682_);
  and _70294_ (_24685_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and _70295_ (_24686_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  or _70296_ (_24687_, _24686_, _24685_);
  or _70297_ (_24688_, _24687_, _24684_);
  or _70298_ (_24689_, _24688_, _24681_);
  or _70299_ (_24690_, _24689_, _24674_);
  and _70300_ (_24691_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and _70301_ (_24692_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or _70302_ (_24693_, _24692_, _24691_);
  and _70303_ (_24694_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  and _70304_ (_24695_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or _70305_ (_24696_, _24695_, _24694_);
  or _70306_ (_24697_, _24696_, _24693_);
  and _70307_ (_24698_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  and _70308_ (_24699_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or _70309_ (_24700_, _24699_, _24698_);
  and _70310_ (_24701_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and _70311_ (_24702_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  or _70312_ (_24703_, _24702_, _24701_);
  or _70313_ (_24704_, _24703_, _24700_);
  or _70314_ (_24705_, _24704_, _24697_);
  and _70315_ (_24706_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and _70316_ (_24707_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  or _70317_ (_24708_, _24707_, _24706_);
  and _70318_ (_24709_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  and _70319_ (_24710_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or _70320_ (_24711_, _24710_, _24709_);
  or _70321_ (_24712_, _24711_, _24708_);
  and _70322_ (_24713_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and _70323_ (_24714_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  or _70324_ (_24715_, _24714_, _24713_);
  and _70325_ (_24716_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  and _70326_ (_24717_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or _70327_ (_24718_, _24717_, _24716_);
  or _70328_ (_24719_, _24718_, _24715_);
  or _70329_ (_24720_, _24719_, _24712_);
  or _70330_ (_24721_, _24720_, _24705_);
  or _70331_ (_24722_, _24721_, _24690_);
  or _70332_ (_24723_, _24722_, _24659_);
  and _70333_ (_24724_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and _70334_ (_24725_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  or _70335_ (_24726_, _24725_, _24724_);
  and _70336_ (_24727_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  and _70337_ (_24728_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or _70338_ (_24729_, _24728_, _24727_);
  or _70339_ (_24730_, _24729_, _24726_);
  and _70340_ (_24731_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and _70341_ (_24732_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  or _70342_ (_24733_, _24732_, _24731_);
  and _70343_ (_24734_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  and _70344_ (_24735_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  or _70345_ (_24736_, _24735_, _24734_);
  or _70346_ (_24737_, _24736_, _24733_);
  or _70347_ (_24738_, _24737_, _24730_);
  and _70348_ (_24739_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  and _70349_ (_24740_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or _70350_ (_24741_, _24740_, _24739_);
  and _70351_ (_24742_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and _70352_ (_24743_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  or _70353_ (_24744_, _24743_, _24742_);
  or _70354_ (_24745_, _24744_, _24741_);
  and _70355_ (_24746_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  and _70356_ (_24747_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or _70357_ (_24748_, _24747_, _24746_);
  and _70358_ (_24749_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and _70359_ (_24750_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  or _70360_ (_24751_, _24750_, _24749_);
  or _70361_ (_24752_, _24751_, _24748_);
  or _70362_ (_24753_, _24752_, _24745_);
  or _70363_ (_24754_, _24753_, _24738_);
  and _70364_ (_24755_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  and _70365_ (_24756_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or _70366_ (_24757_, _24756_, _24755_);
  and _70367_ (_24758_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and _70368_ (_24759_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  or _70369_ (_24760_, _24759_, _24758_);
  or _70370_ (_24761_, _24760_, _24757_);
  and _70371_ (_24762_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  and _70372_ (_24763_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or _70373_ (_24764_, _24763_, _24762_);
  and _70374_ (_24765_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and _70375_ (_24766_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or _70376_ (_24767_, _24766_, _24765_);
  or _70377_ (_24768_, _24767_, _24764_);
  or _70378_ (_24769_, _24768_, _24761_);
  and _70379_ (_24770_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and _70380_ (_24771_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  or _70381_ (_24772_, _24771_, _24770_);
  and _70382_ (_24773_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  and _70383_ (_24774_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or _70384_ (_24775_, _24774_, _24773_);
  or _70385_ (_24776_, _24775_, _24772_);
  and _70386_ (_24777_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and _70387_ (_24778_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  or _70388_ (_24779_, _24778_, _24777_);
  and _70389_ (_24780_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  and _70390_ (_24781_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or _70391_ (_24782_, _24781_, _24780_);
  or _70392_ (_24783_, _24782_, _24779_);
  or _70393_ (_24784_, _24783_, _24776_);
  or _70394_ (_24785_, _24784_, _24769_);
  or _70395_ (_24786_, _24785_, _24754_);
  and _70396_ (_24787_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and _70397_ (_24788_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  or _70398_ (_24789_, _24788_, _24787_);
  and _70399_ (_24790_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  and _70400_ (_24791_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or _70401_ (_24792_, _24791_, _24790_);
  or _70402_ (_24793_, _24792_, _24789_);
  and _70403_ (_24794_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and _70404_ (_24795_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  or _70405_ (_24796_, _24795_, _24794_);
  and _70406_ (_24797_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  and _70407_ (_24798_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  or _70408_ (_24799_, _24798_, _24797_);
  or _70409_ (_24800_, _24799_, _24796_);
  or _70410_ (_24801_, _24800_, _24793_);
  and _70411_ (_24802_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  and _70412_ (_24803_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or _70413_ (_24804_, _24803_, _24802_);
  and _70414_ (_24805_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and _70415_ (_24806_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  or _70416_ (_24807_, _24806_, _24805_);
  or _70417_ (_24808_, _24807_, _24804_);
  and _70418_ (_24809_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  and _70419_ (_24810_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or _70420_ (_24811_, _24810_, _24809_);
  and _70421_ (_24812_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and _70422_ (_24813_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  or _70423_ (_24814_, _24813_, _24812_);
  or _70424_ (_24815_, _24814_, _24811_);
  or _70425_ (_24816_, _24815_, _24808_);
  or _70426_ (_24817_, _24816_, _24801_);
  and _70427_ (_24818_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  and _70428_ (_24819_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or _70429_ (_24820_, _24819_, _24818_);
  and _70430_ (_24821_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and _70431_ (_24822_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  or _70432_ (_24823_, _24822_, _24821_);
  or _70433_ (_24824_, _24823_, _24820_);
  and _70434_ (_24825_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  and _70435_ (_24826_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or _70436_ (_24827_, _24826_, _24825_);
  and _70437_ (_24828_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  and _70438_ (_24829_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  or _70439_ (_24830_, _24829_, _24828_);
  or _70440_ (_24831_, _24830_, _24827_);
  or _70441_ (_24832_, _24831_, _24824_);
  and _70442_ (_24833_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and _70443_ (_24834_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  or _70444_ (_24835_, _24834_, _24833_);
  and _70445_ (_24836_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  and _70446_ (_24837_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or _70447_ (_24838_, _24837_, _24836_);
  or _70448_ (_24839_, _24838_, _24835_);
  and _70449_ (_24840_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and _70450_ (_24841_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  or _70451_ (_24842_, _24841_, _24840_);
  and _70452_ (_24843_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  and _70453_ (_24844_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or _70454_ (_24845_, _24844_, _24843_);
  or _70455_ (_24846_, _24845_, _24842_);
  or _70456_ (_24847_, _24846_, _24839_);
  or _70457_ (_24848_, _24847_, _24832_);
  or _70458_ (_24849_, _24848_, _24817_);
  or _70459_ (_24850_, _24849_, _24786_);
  or _70460_ (_24851_, _24850_, _24723_);
  and _70461_ (_24852_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and _70462_ (_24853_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  or _70463_ (_24854_, _24853_, _24852_);
  and _70464_ (_24855_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  and _70465_ (_24856_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or _70466_ (_24857_, _24856_, _24855_);
  or _70467_ (_24858_, _24857_, _24854_);
  and _70468_ (_24859_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and _70469_ (_24860_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  or _70470_ (_24861_, _24860_, _24859_);
  and _70471_ (_24862_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and _70472_ (_24863_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or _70473_ (_24864_, _24863_, _24862_);
  or _70474_ (_24865_, _24864_, _24861_);
  or _70475_ (_24866_, _24865_, _24858_);
  and _70476_ (_24867_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  and _70477_ (_24868_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or _70478_ (_24869_, _24868_, _24867_);
  and _70479_ (_24870_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and _70480_ (_24871_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  or _70481_ (_24872_, _24871_, _24870_);
  or _70482_ (_24873_, _24872_, _24869_);
  and _70483_ (_24874_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and _70484_ (_24875_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  or _70485_ (_24876_, _24875_, _24874_);
  and _70486_ (_24877_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  and _70487_ (_24878_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or _70488_ (_24879_, _24878_, _24877_);
  or _70489_ (_24880_, _24879_, _24876_);
  or _70490_ (_24881_, _24880_, _24873_);
  or _70491_ (_24882_, _24881_, _24866_);
  and _70492_ (_24883_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  and _70493_ (_24884_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or _70494_ (_24885_, _24884_, _24883_);
  and _70495_ (_24886_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and _70496_ (_24887_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  or _70497_ (_24888_, _24887_, _24886_);
  or _70498_ (_24889_, _24888_, _24885_);
  and _70499_ (_24890_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  and _70500_ (_24891_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or _70501_ (_24892_, _24891_, _24890_);
  and _70502_ (_24893_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  and _70503_ (_24894_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  or _70504_ (_24895_, _24894_, _24893_);
  or _70505_ (_24896_, _24895_, _24892_);
  or _70506_ (_24897_, _24896_, _24889_);
  and _70507_ (_24898_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and _70508_ (_24899_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  or _70509_ (_24900_, _24899_, _24898_);
  and _70510_ (_24901_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  and _70511_ (_24902_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or _70512_ (_24903_, _24902_, _24901_);
  or _70513_ (_24904_, _24903_, _24900_);
  and _70514_ (_24905_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and _70515_ (_24906_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  or _70516_ (_24907_, _24906_, _24905_);
  and _70517_ (_24908_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  and _70518_ (_24909_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or _70519_ (_24910_, _24909_, _24908_);
  or _70520_ (_24911_, _24910_, _24907_);
  or _70521_ (_24912_, _24911_, _24904_);
  or _70522_ (_24913_, _24912_, _24897_);
  or _70523_ (_24914_, _24913_, _24882_);
  and _70524_ (_24915_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and _70525_ (_24916_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  or _70526_ (_24917_, _24916_, _24915_);
  and _70527_ (_24918_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  and _70528_ (_24919_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or _70529_ (_24920_, _24919_, _24918_);
  or _70530_ (_24921_, _24920_, _24917_);
  and _70531_ (_24922_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and _70532_ (_24923_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  or _70533_ (_24924_, _24923_, _24922_);
  and _70534_ (_24925_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  and _70535_ (_24926_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  or _70536_ (_24927_, _24926_, _24925_);
  or _70537_ (_24928_, _24927_, _24924_);
  or _70538_ (_24929_, _24928_, _24921_);
  and _70539_ (_24930_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and _70540_ (_24931_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  or _70541_ (_24932_, _24931_, _24930_);
  and _70542_ (_24933_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  and _70543_ (_24934_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or _70544_ (_24935_, _24934_, _24933_);
  or _70545_ (_24936_, _24935_, _24932_);
  and _70546_ (_24937_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  and _70547_ (_24938_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or _70548_ (_24939_, _24938_, _24937_);
  and _70549_ (_24940_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and _70550_ (_24941_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or _70551_ (_24942_, _24941_, _24940_);
  or _70552_ (_24943_, _24942_, _24939_);
  or _70553_ (_24944_, _24943_, _24936_);
  or _70554_ (_24945_, _24944_, _24929_);
  and _70555_ (_24946_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  and _70556_ (_24947_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or _70557_ (_24948_, _24947_, _24946_);
  and _70558_ (_24949_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and _70559_ (_24950_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or _70560_ (_24951_, _24950_, _24949_);
  or _70561_ (_24952_, _24951_, _24948_);
  and _70562_ (_24953_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  and _70563_ (_24954_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or _70564_ (_24955_, _24954_, _24953_);
  and _70565_ (_24956_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and _70566_ (_24957_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or _70567_ (_24958_, _24957_, _24956_);
  or _70568_ (_24959_, _24958_, _24955_);
  or _70569_ (_24960_, _24959_, _24952_);
  and _70570_ (_24961_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and _70571_ (_24962_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or _70572_ (_24963_, _24962_, _24961_);
  and _70573_ (_24964_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  and _70574_ (_24965_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or _70575_ (_24966_, _24965_, _24964_);
  or _70576_ (_24967_, _24966_, _24963_);
  and _70577_ (_24968_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and _70578_ (_24969_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or _70579_ (_24970_, _24969_, _24968_);
  and _70580_ (_24971_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  and _70581_ (_24972_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or _70582_ (_24973_, _24972_, _24971_);
  or _70583_ (_24974_, _24973_, _24970_);
  or _70584_ (_24975_, _24974_, _24967_);
  or _70585_ (_24976_, _24975_, _24960_);
  or _70586_ (_24977_, _24976_, _24945_);
  or _70587_ (_24978_, _24977_, _24914_);
  and _70588_ (_24979_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  and _70589_ (_24980_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or _70590_ (_24981_, _24980_, _24979_);
  and _70591_ (_24982_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and _70592_ (_24983_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  or _70593_ (_24984_, _24983_, _24982_);
  or _70594_ (_24985_, _24984_, _24981_);
  and _70595_ (_24986_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and _70596_ (_24987_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  or _70597_ (_24988_, _24987_, _24986_);
  and _70598_ (_24989_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  and _70599_ (_24990_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or _70600_ (_24991_, _24990_, _24989_);
  or _70601_ (_24992_, _24991_, _24988_);
  or _70602_ (_24993_, _24992_, _24985_);
  and _70603_ (_24994_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and _70604_ (_24995_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  or _70605_ (_24996_, _24995_, _24994_);
  and _70606_ (_24997_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  and _70607_ (_24998_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or _70608_ (_24999_, _24998_, _24997_);
  or _70609_ (_25000_, _24999_, _24996_);
  and _70610_ (_25001_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and _70611_ (_25002_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  or _70612_ (_25003_, _25002_, _25001_);
  and _70613_ (_25004_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  and _70614_ (_25005_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  or _70615_ (_25006_, _25005_, _25004_);
  or _70616_ (_25007_, _25006_, _25003_);
  or _70617_ (_25008_, _25007_, _25000_);
  or _70618_ (_25009_, _25008_, _24993_);
  and _70619_ (_25010_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  and _70620_ (_25011_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or _70621_ (_25012_, _25011_, _25010_);
  and _70622_ (_25013_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  and _70623_ (_25014_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  or _70624_ (_25015_, _25014_, _25013_);
  or _70625_ (_25016_, _25015_, _25012_);
  and _70626_ (_25017_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  and _70627_ (_25018_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or _70628_ (_25019_, _25018_, _25017_);
  and _70629_ (_25020_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and _70630_ (_25021_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  or _70631_ (_25022_, _25021_, _25020_);
  or _70632_ (_25023_, _25022_, _25019_);
  or _70633_ (_25024_, _25023_, _25016_);
  and _70634_ (_25025_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and _70635_ (_25026_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  or _70636_ (_25027_, _25026_, _25025_);
  and _70637_ (_25028_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  and _70638_ (_25029_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or _70639_ (_25030_, _25029_, _25028_);
  or _70640_ (_25031_, _25030_, _25027_);
  and _70641_ (_25032_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and _70642_ (_25033_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  or _70643_ (_25034_, _25033_, _25032_);
  and _70644_ (_25035_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  and _70645_ (_25036_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or _70646_ (_25037_, _25036_, _25035_);
  or _70647_ (_25038_, _25037_, _25034_);
  or _70648_ (_25039_, _25038_, _25031_);
  or _70649_ (_25040_, _25039_, _25024_);
  or _70650_ (_25041_, _25040_, _25009_);
  and _70651_ (_25042_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and _70652_ (_25043_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  or _70653_ (_25044_, _25043_, _25042_);
  and _70654_ (_25045_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  and _70655_ (_25046_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or _70656_ (_25047_, _25046_, _25045_);
  or _70657_ (_25048_, _25047_, _25044_);
  and _70658_ (_25049_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and _70659_ (_25050_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  or _70660_ (_25051_, _25050_, _25049_);
  and _70661_ (_25052_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and _70662_ (_25053_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or _70663_ (_25054_, _25053_, _25052_);
  or _70664_ (_25055_, _25054_, _25051_);
  or _70665_ (_25056_, _25055_, _25048_);
  and _70666_ (_25057_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  and _70667_ (_25058_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or _70668_ (_25059_, _25058_, _25057_);
  and _70669_ (_25060_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and _70670_ (_25061_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or _70671_ (_25062_, _25061_, _25060_);
  or _70672_ (_25063_, _25062_, _25059_);
  and _70673_ (_25064_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  and _70674_ (_25065_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or _70675_ (_25066_, _25065_, _25064_);
  and _70676_ (_25067_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and _70677_ (_25068_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  or _70678_ (_25069_, _25068_, _25067_);
  or _70679_ (_25070_, _25069_, _25066_);
  or _70680_ (_25071_, _25070_, _25063_);
  or _70681_ (_25072_, _25071_, _25056_);
  and _70682_ (_25073_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  and _70683_ (_25074_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or _70684_ (_25075_, _25074_, _25073_);
  and _70685_ (_25076_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and _70686_ (_25077_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _70687_ (_25078_, _25077_, _25076_);
  or _70688_ (_25079_, _25078_, _25075_);
  and _70689_ (_25080_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and _70690_ (_25081_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and _70691_ (_25082_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or _70692_ (_25083_, _25082_, _25081_);
  or _70693_ (_25084_, _25083_, _25080_);
  or _70694_ (_25085_, _25084_, _25079_);
  and _70695_ (_25086_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _70696_ (_25087_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or _70697_ (_25088_, _25087_, _25086_);
  and _70698_ (_25089_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and _70699_ (_25090_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or _70700_ (_25091_, _25090_, _25089_);
  or _70701_ (_25092_, _25091_, _25088_);
  and _70702_ (_25093_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and _70703_ (_25094_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or _70704_ (_25095_, _25094_, _25093_);
  and _70705_ (_25096_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and _70706_ (_25097_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or _70707_ (_25098_, _25097_, _25096_);
  or _70708_ (_25099_, _25098_, _25095_);
  or _70709_ (_25100_, _25099_, _25092_);
  or _70710_ (_25101_, _25100_, _25085_);
  or _70711_ (_25102_, _25101_, _25072_);
  or _70712_ (_25103_, _25102_, _25041_);
  or _70713_ (_25104_, _25103_, _24978_);
  or _70714_ (_25105_, _25104_, _24851_);
  and _70715_ (_25106_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or _70716_ (_25107_, _25106_, _25105_);
  and _70717_ (_25108_, _25107_, _00006_);
  or _70718_ (_25109_, _25108_, _24596_);
  and _70719_ (_00003_[2], _25109_, _38997_);
  and _70720_ (_25110_, _15589_, iram_op1[1]);
  and _70721_ (_25111_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  and _70722_ (_25112_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or _70723_ (_25113_, _25112_, _25111_);
  and _70724_ (_25114_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and _70725_ (_25115_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  or _70726_ (_25116_, _25115_, _25114_);
  or _70727_ (_25117_, _25116_, _25113_);
  and _70728_ (_25118_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  and _70729_ (_25119_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or _70730_ (_25120_, _25119_, _25118_);
  and _70731_ (_25121_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and _70732_ (_25122_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  or _70733_ (_25123_, _25122_, _25121_);
  or _70734_ (_25124_, _25123_, _25120_);
  or _70735_ (_25125_, _25124_, _25117_);
  and _70736_ (_25126_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and _70737_ (_25127_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  or _70738_ (_25128_, _25127_, _25126_);
  and _70739_ (_25129_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  and _70740_ (_25130_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or _70741_ (_25131_, _25130_, _25129_);
  or _70742_ (_25132_, _25131_, _25128_);
  and _70743_ (_25133_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and _70744_ (_25134_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  or _70745_ (_25135_, _25134_, _25133_);
  and _70746_ (_25136_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and _70747_ (_25137_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or _70748_ (_25138_, _25137_, _25136_);
  or _70749_ (_25139_, _25138_, _25135_);
  or _70750_ (_25140_, _25139_, _25132_);
  or _70751_ (_25141_, _25140_, _25125_);
  and _70752_ (_25142_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  and _70753_ (_25143_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or _70754_ (_25144_, _25143_, _25142_);
  and _70755_ (_25145_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and _70756_ (_25146_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  or _70757_ (_25147_, _25146_, _25145_);
  or _70758_ (_25148_, _25147_, _25144_);
  and _70759_ (_25149_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  and _70760_ (_25150_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or _70761_ (_25151_, _25150_, _25149_);
  and _70762_ (_25152_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and _70763_ (_25153_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or _70764_ (_25154_, _25153_, _25152_);
  or _70765_ (_25155_, _25154_, _25151_);
  or _70766_ (_25156_, _25155_, _25148_);
  and _70767_ (_25157_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and _70768_ (_25158_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  or _70769_ (_25159_, _25158_, _25157_);
  and _70770_ (_25160_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  and _70771_ (_25161_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or _70772_ (_25162_, _25161_, _25160_);
  or _70773_ (_25163_, _25162_, _25159_);
  and _70774_ (_25164_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and _70775_ (_25165_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  or _70776_ (_25166_, _25165_, _25164_);
  and _70777_ (_25167_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  and _70778_ (_25168_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or _70779_ (_25169_, _25168_, _25167_);
  or _70780_ (_25170_, _25169_, _25166_);
  or _70781_ (_25171_, _25170_, _25163_);
  or _70782_ (_25172_, _25171_, _25156_);
  or _70783_ (_25173_, _25172_, _25141_);
  and _70784_ (_25174_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and _70785_ (_25175_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  or _70786_ (_25176_, _25175_, _25174_);
  and _70787_ (_25177_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  and _70788_ (_25178_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or _70789_ (_25179_, _25178_, _25177_);
  or _70790_ (_25180_, _25179_, _25176_);
  and _70791_ (_25181_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and _70792_ (_25182_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  or _70793_ (_25183_, _25182_, _25181_);
  and _70794_ (_25184_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and _70795_ (_25185_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or _70796_ (_25186_, _25185_, _25184_);
  or _70797_ (_25187_, _25186_, _25183_);
  or _70798_ (_25188_, _25187_, _25180_);
  and _70799_ (_25189_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  and _70800_ (_25190_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or _70801_ (_25191_, _25190_, _25189_);
  and _70802_ (_25192_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and _70803_ (_25193_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  or _70804_ (_25194_, _25193_, _25192_);
  or _70805_ (_25195_, _25194_, _25191_);
  and _70806_ (_25196_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  and _70807_ (_25197_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or _70808_ (_25198_, _25197_, _25196_);
  and _70809_ (_25199_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and _70810_ (_25200_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  or _70811_ (_25201_, _25200_, _25199_);
  or _70812_ (_25202_, _25201_, _25198_);
  or _70813_ (_25203_, _25202_, _25195_);
  or _70814_ (_25204_, _25203_, _25188_);
  and _70815_ (_25205_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  and _70816_ (_25206_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or _70817_ (_25207_, _25206_, _25205_);
  and _70818_ (_25208_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and _70819_ (_25209_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  or _70820_ (_25210_, _25209_, _25208_);
  or _70821_ (_25211_, _25210_, _25207_);
  and _70822_ (_25212_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  and _70823_ (_25213_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or _70824_ (_25214_, _25213_, _25212_);
  and _70825_ (_25215_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and _70826_ (_25216_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or _70827_ (_25217_, _25216_, _25215_);
  or _70828_ (_25218_, _25217_, _25214_);
  or _70829_ (_25219_, _25218_, _25211_);
  and _70830_ (_25220_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and _70831_ (_25221_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  or _70832_ (_25222_, _25221_, _25220_);
  and _70833_ (_25223_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  and _70834_ (_25224_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or _70835_ (_25225_, _25224_, _25223_);
  or _70836_ (_25226_, _25225_, _25222_);
  and _70837_ (_25227_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and _70838_ (_25228_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  or _70839_ (_25229_, _25228_, _25227_);
  and _70840_ (_25230_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  and _70841_ (_25231_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or _70842_ (_25232_, _25231_, _25230_);
  or _70843_ (_25233_, _25232_, _25229_);
  or _70844_ (_25234_, _25233_, _25226_);
  or _70845_ (_25235_, _25234_, _25219_);
  or _70846_ (_25236_, _25235_, _25204_);
  or _70847_ (_25237_, _25236_, _25173_);
  and _70848_ (_25238_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  and _70849_ (_25239_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or _70850_ (_25240_, _25239_, _25238_);
  and _70851_ (_25241_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and _70852_ (_25242_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  or _70853_ (_25243_, _25242_, _25241_);
  or _70854_ (_25244_, _25243_, _25240_);
  and _70855_ (_25245_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  and _70856_ (_25246_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or _70857_ (_25247_, _25246_, _25245_);
  and _70858_ (_25248_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and _70859_ (_25249_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  or _70860_ (_25250_, _25249_, _25248_);
  or _70861_ (_25251_, _25250_, _25247_);
  or _70862_ (_25252_, _25251_, _25244_);
  and _70863_ (_25253_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and _70864_ (_25254_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  or _70865_ (_25255_, _25254_, _25253_);
  and _70866_ (_25256_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  and _70867_ (_25257_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  or _70868_ (_25258_, _25257_, _25256_);
  or _70869_ (_25259_, _25258_, _25255_);
  and _70870_ (_25260_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and _70871_ (_25261_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  or _70872_ (_25262_, _25261_, _25260_);
  and _70873_ (_25263_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  and _70874_ (_25264_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or _70875_ (_25265_, _25264_, _25263_);
  or _70876_ (_25266_, _25265_, _25262_);
  or _70877_ (_25267_, _25266_, _25259_);
  or _70878_ (_25268_, _25267_, _25252_);
  and _70879_ (_25269_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  and _70880_ (_25270_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or _70881_ (_25271_, _25270_, _25269_);
  and _70882_ (_25272_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and _70883_ (_25273_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  or _70884_ (_25274_, _25273_, _25272_);
  or _70885_ (_25275_, _25274_, _25271_);
  and _70886_ (_25276_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  and _70887_ (_25277_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or _70888_ (_25278_, _25277_, _25276_);
  and _70889_ (_25279_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and _70890_ (_25280_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or _70891_ (_25281_, _25280_, _25279_);
  or _70892_ (_25282_, _25281_, _25278_);
  or _70893_ (_25283_, _25282_, _25275_);
  and _70894_ (_25284_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and _70895_ (_25285_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  or _70896_ (_25286_, _25285_, _25284_);
  and _70897_ (_25287_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  and _70898_ (_25288_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or _70899_ (_25289_, _25288_, _25287_);
  or _70900_ (_25290_, _25289_, _25286_);
  and _70901_ (_25291_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and _70902_ (_25292_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  or _70903_ (_25293_, _25292_, _25291_);
  and _70904_ (_25294_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  and _70905_ (_25295_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or _70906_ (_25296_, _25295_, _25294_);
  or _70907_ (_25297_, _25296_, _25293_);
  or _70908_ (_25298_, _25297_, _25290_);
  or _70909_ (_25299_, _25298_, _25283_);
  or _70910_ (_25300_, _25299_, _25268_);
  and _70911_ (_25301_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  and _70912_ (_25302_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or _70913_ (_25303_, _25302_, _25301_);
  and _70914_ (_25304_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and _70915_ (_25305_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  or _70916_ (_25306_, _25305_, _25304_);
  or _70917_ (_25307_, _25306_, _25303_);
  and _70918_ (_25308_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  and _70919_ (_25309_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or _70920_ (_25310_, _25309_, _25308_);
  and _70921_ (_25311_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and _70922_ (_25312_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or _70923_ (_25313_, _25312_, _25311_);
  or _70924_ (_25314_, _25313_, _25310_);
  or _70925_ (_25315_, _25314_, _25307_);
  and _70926_ (_25316_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and _70927_ (_25317_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  or _70928_ (_25318_, _25317_, _25316_);
  and _70929_ (_25319_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  and _70930_ (_25320_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or _70931_ (_25321_, _25320_, _25319_);
  or _70932_ (_25322_, _25321_, _25318_);
  and _70933_ (_25323_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and _70934_ (_25324_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  or _70935_ (_25325_, _25324_, _25323_);
  and _70936_ (_25326_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  and _70937_ (_25327_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or _70938_ (_25328_, _25327_, _25326_);
  or _70939_ (_25329_, _25328_, _25325_);
  or _70940_ (_25330_, _25329_, _25322_);
  or _70941_ (_25331_, _25330_, _25315_);
  and _70942_ (_25332_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and _70943_ (_25333_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  or _70944_ (_25334_, _25333_, _25332_);
  and _70945_ (_25335_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  and _70946_ (_25336_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or _70947_ (_25337_, _25336_, _25335_);
  or _70948_ (_25338_, _25337_, _25334_);
  and _70949_ (_25339_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and _70950_ (_25340_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  or _70951_ (_25341_, _25340_, _25339_);
  and _70952_ (_25342_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  and _70953_ (_25343_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  or _70954_ (_25344_, _25343_, _25342_);
  or _70955_ (_25345_, _25344_, _25341_);
  or _70956_ (_25346_, _25345_, _25338_);
  and _70957_ (_25347_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  and _70958_ (_25348_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or _70959_ (_25349_, _25348_, _25347_);
  and _70960_ (_25350_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and _70961_ (_25351_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  or _70962_ (_25352_, _25351_, _25350_);
  or _70963_ (_25353_, _25352_, _25349_);
  and _70964_ (_25354_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  and _70965_ (_25355_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or _70966_ (_25356_, _25355_, _25354_);
  and _70967_ (_25357_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and _70968_ (_25358_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  or _70969_ (_25359_, _25358_, _25357_);
  or _70970_ (_25360_, _25359_, _25356_);
  or _70971_ (_25361_, _25360_, _25353_);
  or _70972_ (_25362_, _25361_, _25346_);
  or _70973_ (_25363_, _25362_, _25331_);
  or _70974_ (_25364_, _25363_, _25300_);
  or _70975_ (_25365_, _25364_, _25237_);
  and _70976_ (_25366_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  and _70977_ (_25367_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or _70978_ (_25368_, _25367_, _25366_);
  and _70979_ (_25369_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and _70980_ (_25370_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  or _70981_ (_25371_, _25370_, _25369_);
  or _70982_ (_25372_, _25371_, _25368_);
  and _70983_ (_25373_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  and _70984_ (_25374_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or _70985_ (_25375_, _25374_, _25373_);
  and _70986_ (_25376_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and _70987_ (_25377_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  or _70988_ (_25378_, _25377_, _25376_);
  or _70989_ (_25379_, _25378_, _25375_);
  or _70990_ (_25380_, _25379_, _25372_);
  and _70991_ (_25381_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and _70992_ (_25382_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  or _70993_ (_25383_, _25382_, _25381_);
  and _70994_ (_25384_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  and _70995_ (_25385_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  or _70996_ (_25386_, _25385_, _25384_);
  or _70997_ (_25387_, _25386_, _25383_);
  and _70998_ (_25388_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and _70999_ (_25389_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  or _71000_ (_25390_, _25389_, _25388_);
  and _71001_ (_25391_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  and _71002_ (_25392_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or _71003_ (_25393_, _25392_, _25391_);
  or _71004_ (_25394_, _25393_, _25390_);
  or _71005_ (_25395_, _25394_, _25387_);
  or _71006_ (_25396_, _25395_, _25380_);
  and _71007_ (_25397_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  and _71008_ (_25398_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or _71009_ (_25399_, _25398_, _25397_);
  and _71010_ (_25400_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and _71011_ (_25401_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  or _71012_ (_25402_, _25401_, _25400_);
  or _71013_ (_25403_, _25402_, _25399_);
  and _71014_ (_25404_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  and _71015_ (_25405_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or _71016_ (_25406_, _25405_, _25404_);
  and _71017_ (_25407_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and _71018_ (_25408_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or _71019_ (_25409_, _25408_, _25407_);
  or _71020_ (_25410_, _25409_, _25406_);
  or _71021_ (_25411_, _25410_, _25403_);
  and _71022_ (_25412_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and _71023_ (_25413_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  or _71024_ (_25414_, _25413_, _25412_);
  and _71025_ (_25415_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  and _71026_ (_25416_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or _71027_ (_25417_, _25416_, _25415_);
  or _71028_ (_25418_, _25417_, _25414_);
  and _71029_ (_25419_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and _71030_ (_25420_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  or _71031_ (_25421_, _25420_, _25419_);
  and _71032_ (_25422_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  and _71033_ (_25423_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or _71034_ (_25424_, _25423_, _25422_);
  or _71035_ (_25425_, _25424_, _25421_);
  or _71036_ (_25426_, _25425_, _25418_);
  or _71037_ (_25427_, _25426_, _25411_);
  or _71038_ (_25428_, _25427_, _25396_);
  and _71039_ (_25429_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  and _71040_ (_25430_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or _71041_ (_25431_, _25430_, _25429_);
  and _71042_ (_25432_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  and _71043_ (_25433_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  or _71044_ (_25434_, _25433_, _25432_);
  or _71045_ (_25435_, _25434_, _25431_);
  and _71046_ (_25436_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  and _71047_ (_25437_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or _71048_ (_25438_, _25437_, _25436_);
  and _71049_ (_25439_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and _71050_ (_25440_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  or _71051_ (_25441_, _25440_, _25439_);
  or _71052_ (_25442_, _25441_, _25438_);
  or _71053_ (_25443_, _25442_, _25435_);
  and _71054_ (_25444_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and _71055_ (_25445_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  or _71056_ (_25446_, _25445_, _25444_);
  and _71057_ (_25447_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  and _71058_ (_25448_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or _71059_ (_25449_, _25448_, _25447_);
  or _71060_ (_25450_, _25449_, _25446_);
  and _71061_ (_25451_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and _71062_ (_25452_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  or _71063_ (_25453_, _25452_, _25451_);
  and _71064_ (_25454_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  and _71065_ (_25455_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  or _71066_ (_25456_, _25455_, _25454_);
  or _71067_ (_25457_, _25456_, _25453_);
  or _71068_ (_25458_, _25457_, _25450_);
  or _71069_ (_25459_, _25458_, _25443_);
  and _71070_ (_25460_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  and _71071_ (_25461_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or _71072_ (_25462_, _25461_, _25460_);
  and _71073_ (_25463_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and _71074_ (_25464_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or _71075_ (_25465_, _25464_, _25463_);
  or _71076_ (_25466_, _25465_, _25462_);
  and _71077_ (_25467_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  and _71078_ (_25468_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or _71079_ (_25469_, _25468_, _25467_);
  and _71080_ (_25470_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  and _71081_ (_25471_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or _71082_ (_25472_, _25471_, _25470_);
  or _71083_ (_25473_, _25472_, _25469_);
  or _71084_ (_25474_, _25473_, _25466_);
  and _71085_ (_25475_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  and _71086_ (_25476_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or _71087_ (_25477_, _25476_, _25475_);
  and _71088_ (_25478_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  and _71089_ (_25479_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or _71090_ (_25480_, _25479_, _25478_);
  or _71091_ (_25481_, _25480_, _25477_);
  and _71092_ (_25482_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and _71093_ (_25483_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or _71094_ (_25484_, _25483_, _25482_);
  and _71095_ (_25485_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  and _71096_ (_25486_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or _71097_ (_25487_, _25486_, _25485_);
  or _71098_ (_25488_, _25487_, _25484_);
  or _71099_ (_25489_, _25488_, _25481_);
  or _71100_ (_25490_, _25489_, _25474_);
  or _71101_ (_25491_, _25490_, _25459_);
  or _71102_ (_25492_, _25491_, _25428_);
  and _71103_ (_25493_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and _71104_ (_25494_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  or _71105_ (_25495_, _25494_, _25493_);
  and _71106_ (_25496_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  and _71107_ (_25497_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  or _71108_ (_25498_, _25497_, _25496_);
  or _71109_ (_25499_, _25498_, _25495_);
  and _71110_ (_25500_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and _71111_ (_25501_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  or _71112_ (_25502_, _25501_, _25500_);
  and _71113_ (_25503_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  and _71114_ (_25504_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or _71115_ (_25505_, _25504_, _25503_);
  or _71116_ (_25506_, _25505_, _25502_);
  or _71117_ (_25507_, _25506_, _25499_);
  and _71118_ (_25508_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  and _71119_ (_25509_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or _71120_ (_25510_, _25509_, _25508_);
  and _71121_ (_25511_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and _71122_ (_25512_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  or _71123_ (_25513_, _25512_, _25511_);
  or _71124_ (_25514_, _25513_, _25510_);
  and _71125_ (_25515_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  and _71126_ (_25516_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or _71127_ (_25517_, _25516_, _25515_);
  and _71128_ (_25518_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and _71129_ (_25519_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  or _71130_ (_25520_, _25519_, _25518_);
  or _71131_ (_25521_, _25520_, _25517_);
  or _71132_ (_25522_, _25521_, _25514_);
  or _71133_ (_25523_, _25522_, _25507_);
  and _71134_ (_25524_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  and _71135_ (_25525_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or _71136_ (_25526_, _25525_, _25524_);
  and _71137_ (_25527_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and _71138_ (_25528_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  or _71139_ (_25529_, _25528_, _25527_);
  or _71140_ (_25530_, _25529_, _25526_);
  and _71141_ (_25531_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  and _71142_ (_25532_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or _71143_ (_25533_, _25532_, _25531_);
  and _71144_ (_25534_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and _71145_ (_25535_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or _71146_ (_25536_, _25535_, _25534_);
  or _71147_ (_25537_, _25536_, _25533_);
  or _71148_ (_25538_, _25537_, _25530_);
  and _71149_ (_25539_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and _71150_ (_25540_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  or _71151_ (_25541_, _25540_, _25539_);
  and _71152_ (_25542_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  and _71153_ (_25543_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or _71154_ (_25544_, _25543_, _25542_);
  or _71155_ (_25545_, _25544_, _25541_);
  and _71156_ (_25546_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and _71157_ (_25547_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  or _71158_ (_25548_, _25547_, _25546_);
  and _71159_ (_25549_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  and _71160_ (_25550_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or _71161_ (_25551_, _25550_, _25549_);
  or _71162_ (_25552_, _25551_, _25548_);
  or _71163_ (_25553_, _25552_, _25545_);
  or _71164_ (_25554_, _25553_, _25538_);
  or _71165_ (_25555_, _25554_, _25523_);
  and _71166_ (_25556_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  and _71167_ (_25557_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or _71168_ (_25558_, _25557_, _25556_);
  and _71169_ (_25559_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and _71170_ (_25560_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  or _71171_ (_25561_, _25560_, _25559_);
  or _71172_ (_25562_, _25561_, _25558_);
  and _71173_ (_25563_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  and _71174_ (_25564_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or _71175_ (_25565_, _25564_, _25563_);
  and _71176_ (_25566_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and _71177_ (_25567_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  or _71178_ (_25568_, _25567_, _25566_);
  or _71179_ (_25569_, _25568_, _25565_);
  or _71180_ (_25570_, _25569_, _25562_);
  and _71181_ (_25571_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and _71182_ (_25572_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  or _71183_ (_25573_, _25572_, _25571_);
  and _71184_ (_25574_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  and _71185_ (_25575_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  or _71186_ (_25576_, _25575_, _25574_);
  or _71187_ (_25577_, _25576_, _25573_);
  and _71188_ (_25578_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and _71189_ (_25579_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  or _71190_ (_25580_, _25579_, _25578_);
  and _71191_ (_25581_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  and _71192_ (_25582_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or _71193_ (_25583_, _25582_, _25581_);
  or _71194_ (_25584_, _25583_, _25580_);
  or _71195_ (_25585_, _25584_, _25577_);
  or _71196_ (_25586_, _25585_, _25570_);
  and _71197_ (_25587_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _71198_ (_25588_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or _71199_ (_25589_, _25588_, _25587_);
  and _71200_ (_25590_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and _71201_ (_25591_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or _71202_ (_25592_, _25591_, _25590_);
  or _71203_ (_25593_, _25592_, _25589_);
  and _71204_ (_25594_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and _71205_ (_25595_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or _71206_ (_25596_, _25595_, _25594_);
  and _71207_ (_25597_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and _71208_ (_25598_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or _71209_ (_25599_, _25598_, _25597_);
  or _71210_ (_25600_, _25599_, _25596_);
  or _71211_ (_25601_, _25600_, _25593_);
  and _71212_ (_25602_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and _71213_ (_25603_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or _71214_ (_25604_, _25603_, _25602_);
  and _71215_ (_25605_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and _71216_ (_25606_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or _71217_ (_25607_, _25606_, _25605_);
  or _71218_ (_25608_, _25607_, _25604_);
  and _71219_ (_25609_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and _71220_ (_25610_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and _71221_ (_25611_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _71222_ (_25612_, _25611_, _25610_);
  or _71223_ (_25613_, _25612_, _25609_);
  or _71224_ (_25614_, _25613_, _25608_);
  or _71225_ (_25615_, _25614_, _25601_);
  or _71226_ (_25616_, _25615_, _25586_);
  or _71227_ (_25617_, _25616_, _25555_);
  or _71228_ (_25618_, _25617_, _25492_);
  or _71229_ (_25619_, _25618_, _25365_);
  and _71230_ (_25620_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or _71231_ (_25621_, _25620_, _25619_);
  and _71232_ (_25622_, _25621_, _00006_);
  or _71233_ (_25623_, _25622_, _25110_);
  and _71234_ (_00003_[1], _25623_, _38997_);
  and _71235_ (_25624_, _15589_, iram_op1[0]);
  and _71236_ (_25625_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and _71237_ (_25626_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  or _71238_ (_25627_, _25626_, _25625_);
  and _71239_ (_25628_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  and _71240_ (_25629_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or _71241_ (_25630_, _25629_, _25628_);
  or _71242_ (_25631_, _25630_, _25627_);
  and _71243_ (_25632_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and _71244_ (_25633_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  or _71245_ (_25634_, _25633_, _25632_);
  and _71246_ (_25635_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  and _71247_ (_25636_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or _71248_ (_25637_, _25636_, _25635_);
  or _71249_ (_25638_, _25637_, _25634_);
  or _71250_ (_25639_, _25638_, _25631_);
  and _71251_ (_25640_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  and _71252_ (_25641_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or _71253_ (_25642_, _25641_, _25640_);
  and _71254_ (_25643_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and _71255_ (_25644_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or _71256_ (_25645_, _25644_, _25643_);
  or _71257_ (_25646_, _25645_, _25642_);
  and _71258_ (_25647_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  and _71259_ (_25648_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or _71260_ (_25649_, _25648_, _25647_);
  and _71261_ (_25650_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and _71262_ (_25651_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  or _71263_ (_25652_, _25651_, _25650_);
  or _71264_ (_25653_, _25652_, _25649_);
  or _71265_ (_25654_, _25653_, _25646_);
  or _71266_ (_25655_, _25654_, _25639_);
  and _71267_ (_25656_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and _71268_ (_25657_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  or _71269_ (_25658_, _25657_, _25656_);
  and _71270_ (_25659_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  and _71271_ (_25660_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or _71272_ (_25661_, _25660_, _25659_);
  or _71273_ (_25662_, _25661_, _25658_);
  and _71274_ (_25663_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and _71275_ (_25664_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  or _71276_ (_25665_, _25664_, _25663_);
  and _71277_ (_25666_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  and _71278_ (_25667_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  or _71279_ (_25668_, _25667_, _25666_);
  or _71280_ (_25669_, _25668_, _25665_);
  or _71281_ (_25670_, _25669_, _25662_);
  and _71282_ (_25671_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  and _71283_ (_25672_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or _71284_ (_25673_, _25672_, _25671_);
  and _71285_ (_25674_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and _71286_ (_25675_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  or _71287_ (_25676_, _25675_, _25674_);
  or _71288_ (_25677_, _25676_, _25673_);
  and _71289_ (_25678_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  and _71290_ (_25679_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or _71291_ (_25680_, _25679_, _25678_);
  and _71292_ (_25681_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and _71293_ (_25682_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  or _71294_ (_25683_, _25682_, _25681_);
  or _71295_ (_25684_, _25683_, _25680_);
  or _71296_ (_25685_, _25684_, _25677_);
  or _71297_ (_25686_, _25685_, _25670_);
  or _71298_ (_25687_, _25686_, _25655_);
  and _71299_ (_25688_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and _71300_ (_25689_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  or _71301_ (_25690_, _25689_, _25688_);
  and _71302_ (_25691_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and _71303_ (_25692_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or _71304_ (_25693_, _25692_, _25691_);
  or _71305_ (_25694_, _25693_, _25690_);
  and _71306_ (_25695_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and _71307_ (_25696_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  or _71308_ (_25697_, _25696_, _25695_);
  and _71309_ (_25698_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  and _71310_ (_25699_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or _71311_ (_25700_, _25699_, _25698_);
  or _71312_ (_25701_, _25700_, _25697_);
  or _71313_ (_25702_, _25701_, _25694_);
  and _71314_ (_25703_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  and _71315_ (_25704_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or _71316_ (_25705_, _25704_, _25703_);
  and _71317_ (_25706_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and _71318_ (_25707_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  or _71319_ (_25708_, _25707_, _25706_);
  or _71320_ (_25709_, _25708_, _25705_);
  and _71321_ (_25710_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  and _71322_ (_25711_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or _71323_ (_25712_, _25711_, _25710_);
  and _71324_ (_25713_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and _71325_ (_25714_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or _71326_ (_25715_, _25714_, _25713_);
  or _71327_ (_25716_, _25715_, _25712_);
  or _71328_ (_25717_, _25716_, _25709_);
  or _71329_ (_25718_, _25717_, _25702_);
  and _71330_ (_25719_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  and _71331_ (_25720_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or _71332_ (_25721_, _25720_, _25719_);
  and _71333_ (_25722_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  and _71334_ (_25723_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or _71335_ (_25724_, _25723_, _25722_);
  or _71336_ (_25725_, _25724_, _25721_);
  and _71337_ (_25726_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and _71338_ (_25727_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or _71339_ (_25728_, _25727_, _25726_);
  and _71340_ (_25729_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  and _71341_ (_25730_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or _71342_ (_25731_, _25730_, _25729_);
  or _71343_ (_25732_, _25731_, _25728_);
  or _71344_ (_25733_, _25732_, _25725_);
  and _71345_ (_25734_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  and _71346_ (_25735_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or _71347_ (_25736_, _25735_, _25734_);
  and _71348_ (_25737_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  and _71349_ (_25738_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or _71350_ (_25739_, _25738_, _25737_);
  or _71351_ (_25740_, _25739_, _25736_);
  and _71352_ (_25741_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  and _71353_ (_25742_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or _71354_ (_25743_, _25742_, _25741_);
  and _71355_ (_25744_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and _71356_ (_25745_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or _71357_ (_25746_, _25745_, _25744_);
  or _71358_ (_25747_, _25746_, _25743_);
  or _71359_ (_25748_, _25747_, _25740_);
  or _71360_ (_25749_, _25748_, _25733_);
  or _71361_ (_25750_, _25749_, _25718_);
  or _71362_ (_25751_, _25750_, _25687_);
  and _71363_ (_25752_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  and _71364_ (_25753_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or _71365_ (_25754_, _25753_, _25752_);
  and _71366_ (_25755_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and _71367_ (_25756_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  or _71368_ (_25757_, _25756_, _25755_);
  or _71369_ (_25758_, _25757_, _25754_);
  and _71370_ (_25759_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  and _71371_ (_25760_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or _71372_ (_25761_, _25760_, _25759_);
  and _71373_ (_25762_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and _71374_ (_25763_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  or _71375_ (_25764_, _25763_, _25762_);
  or _71376_ (_25765_, _25764_, _25761_);
  or _71377_ (_25766_, _25765_, _25758_);
  and _71378_ (_25767_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and _71379_ (_25768_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  or _71380_ (_25769_, _25768_, _25767_);
  and _71381_ (_25770_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  and _71382_ (_25771_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  or _71383_ (_25772_, _25771_, _25770_);
  or _71384_ (_25773_, _25772_, _25769_);
  and _71385_ (_25774_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and _71386_ (_25775_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  or _71387_ (_25776_, _25775_, _25774_);
  and _71388_ (_25777_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  and _71389_ (_25778_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or _71390_ (_25779_, _25778_, _25777_);
  or _71391_ (_25780_, _25779_, _25776_);
  or _71392_ (_25781_, _25780_, _25773_);
  or _71393_ (_25782_, _25781_, _25766_);
  and _71394_ (_25783_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  and _71395_ (_25784_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or _71396_ (_25785_, _25784_, _25783_);
  and _71397_ (_25786_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and _71398_ (_25787_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  or _71399_ (_25788_, _25787_, _25786_);
  or _71400_ (_25789_, _25788_, _25785_);
  and _71401_ (_25790_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and _71402_ (_25791_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or _71403_ (_25792_, _25791_, _25790_);
  and _71404_ (_25793_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and _71405_ (_25794_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or _71406_ (_25795_, _25794_, _25793_);
  or _71407_ (_25796_, _25795_, _25792_);
  or _71408_ (_25797_, _25796_, _25789_);
  and _71409_ (_25798_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and _71410_ (_25799_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  or _71411_ (_25800_, _25799_, _25798_);
  and _71412_ (_25801_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and _71413_ (_25802_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or _71414_ (_25803_, _25802_, _25801_);
  or _71415_ (_25804_, _25803_, _25800_);
  and _71416_ (_25805_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and _71417_ (_25806_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  or _71418_ (_25807_, _25806_, _25805_);
  and _71419_ (_25808_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  and _71420_ (_25809_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or _71421_ (_25810_, _25809_, _25808_);
  or _71422_ (_25811_, _25810_, _25807_);
  or _71423_ (_25812_, _25811_, _25804_);
  or _71424_ (_25813_, _25812_, _25797_);
  or _71425_ (_25814_, _25813_, _25782_);
  and _71426_ (_25815_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  and _71427_ (_25816_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or _71428_ (_25817_, _25816_, _25815_);
  and _71429_ (_25818_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and _71430_ (_25819_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  or _71431_ (_25820_, _25819_, _25818_);
  or _71432_ (_25821_, _25820_, _25817_);
  and _71433_ (_25822_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  and _71434_ (_25823_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or _71435_ (_25824_, _25823_, _25822_);
  and _71436_ (_25825_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and _71437_ (_25826_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  or _71438_ (_25827_, _25826_, _25825_);
  or _71439_ (_25828_, _25827_, _25824_);
  or _71440_ (_25829_, _25828_, _25821_);
  and _71441_ (_25830_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and _71442_ (_25831_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  or _71443_ (_25832_, _25831_, _25830_);
  and _71444_ (_25833_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  and _71445_ (_25834_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or _71446_ (_25835_, _25834_, _25833_);
  or _71447_ (_25836_, _25835_, _25832_);
  and _71448_ (_25837_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and _71449_ (_25838_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  or _71450_ (_25839_, _25838_, _25837_);
  and _71451_ (_25840_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  and _71452_ (_25841_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  or _71453_ (_25842_, _25841_, _25840_);
  or _71454_ (_25843_, _25842_, _25839_);
  or _71455_ (_25844_, _25843_, _25836_);
  or _71456_ (_25845_, _25844_, _25829_);
  and _71457_ (_25846_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and _71458_ (_25847_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  or _71459_ (_25848_, _25847_, _25846_);
  and _71460_ (_25849_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  and _71461_ (_25850_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or _71462_ (_25851_, _25850_, _25849_);
  or _71463_ (_25852_, _25851_, _25848_);
  and _71464_ (_25853_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and _71465_ (_25854_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  or _71466_ (_25855_, _25854_, _25853_);
  and _71467_ (_25856_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  and _71468_ (_25857_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or _71469_ (_25858_, _25857_, _25856_);
  or _71470_ (_25859_, _25858_, _25855_);
  or _71471_ (_25860_, _25859_, _25852_);
  and _71472_ (_25861_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  and _71473_ (_25862_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or _71474_ (_25863_, _25862_, _25861_);
  and _71475_ (_25864_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and _71476_ (_25865_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  or _71477_ (_25866_, _25865_, _25864_);
  or _71478_ (_25867_, _25866_, _25863_);
  and _71479_ (_25868_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  and _71480_ (_25869_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or _71481_ (_25870_, _25869_, _25868_);
  and _71482_ (_25871_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and _71483_ (_25872_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or _71484_ (_25873_, _25872_, _25871_);
  or _71485_ (_25874_, _25873_, _25870_);
  or _71486_ (_25875_, _25874_, _25867_);
  or _71487_ (_25876_, _25875_, _25860_);
  or _71488_ (_25877_, _25876_, _25845_);
  or _71489_ (_25878_, _25877_, _25814_);
  or _71490_ (_25879_, _25878_, _25751_);
  and _71491_ (_25880_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and _71492_ (_25881_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  or _71493_ (_25882_, _25881_, _25880_);
  and _71494_ (_25883_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  and _71495_ (_25884_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or _71496_ (_25885_, _25884_, _25883_);
  or _71497_ (_25886_, _25885_, _25882_);
  and _71498_ (_25887_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and _71499_ (_25888_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  or _71500_ (_25889_, _25888_, _25887_);
  and _71501_ (_25890_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and _71502_ (_25891_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or _71503_ (_25892_, _25891_, _25890_);
  or _71504_ (_25893_, _25892_, _25889_);
  or _71505_ (_25894_, _25893_, _25886_);
  and _71506_ (_25895_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  and _71507_ (_25896_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or _71508_ (_25897_, _25896_, _25895_);
  and _71509_ (_25898_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and _71510_ (_25899_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  or _71511_ (_25900_, _25899_, _25898_);
  or _71512_ (_25901_, _25900_, _25897_);
  and _71513_ (_25902_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  and _71514_ (_25903_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or _71515_ (_25904_, _25903_, _25902_);
  and _71516_ (_25905_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and _71517_ (_25906_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  or _71518_ (_25907_, _25906_, _25905_);
  or _71519_ (_25908_, _25907_, _25904_);
  or _71520_ (_25909_, _25908_, _25901_);
  or _71521_ (_25910_, _25909_, _25894_);
  and _71522_ (_25911_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  and _71523_ (_25912_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or _71524_ (_25913_, _25912_, _25911_);
  and _71525_ (_25914_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and _71526_ (_25915_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  or _71527_ (_25916_, _25915_, _25914_);
  or _71528_ (_25917_, _25916_, _25913_);
  and _71529_ (_25918_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  and _71530_ (_25919_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or _71531_ (_25920_, _25919_, _25918_);
  and _71532_ (_25921_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and _71533_ (_25922_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or _71534_ (_25923_, _25922_, _25921_);
  or _71535_ (_25924_, _25923_, _25920_);
  or _71536_ (_25925_, _25924_, _25917_);
  and _71537_ (_25926_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and _71538_ (_25927_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  or _71539_ (_25928_, _25927_, _25926_);
  and _71540_ (_25929_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  and _71541_ (_25930_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or _71542_ (_25931_, _25930_, _25929_);
  or _71543_ (_25932_, _25931_, _25928_);
  and _71544_ (_25933_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and _71545_ (_25934_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  or _71546_ (_25935_, _25934_, _25933_);
  and _71547_ (_25936_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  and _71548_ (_25937_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or _71549_ (_25938_, _25937_, _25936_);
  or _71550_ (_25939_, _25938_, _25935_);
  or _71551_ (_25940_, _25939_, _25932_);
  or _71552_ (_25941_, _25940_, _25925_);
  or _71553_ (_25942_, _25941_, _25910_);
  and _71554_ (_25943_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and _71555_ (_25944_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  or _71556_ (_25945_, _25944_, _25943_);
  and _71557_ (_25946_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  and _71558_ (_25947_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or _71559_ (_25948_, _25947_, _25946_);
  or _71560_ (_25949_, _25948_, _25945_);
  and _71561_ (_25950_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and _71562_ (_25951_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  or _71563_ (_25952_, _25951_, _25950_);
  and _71564_ (_25953_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and _71565_ (_25954_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or _71566_ (_25955_, _25954_, _25953_);
  or _71567_ (_25956_, _25955_, _25952_);
  or _71568_ (_25957_, _25956_, _25949_);
  and _71569_ (_25958_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  and _71570_ (_25959_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or _71571_ (_25960_, _25959_, _25958_);
  and _71572_ (_25961_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and _71573_ (_25962_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  or _71574_ (_25963_, _25962_, _25961_);
  or _71575_ (_25964_, _25963_, _25960_);
  and _71576_ (_25965_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  and _71577_ (_25966_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or _71578_ (_25967_, _25966_, _25965_);
  and _71579_ (_25968_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and _71580_ (_25969_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  or _71581_ (_25970_, _25969_, _25968_);
  or _71582_ (_25971_, _25970_, _25967_);
  or _71583_ (_25972_, _25971_, _25964_);
  or _71584_ (_25973_, _25972_, _25957_);
  and _71585_ (_25974_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  and _71586_ (_25975_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or _71587_ (_25976_, _25975_, _25974_);
  and _71588_ (_25977_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and _71589_ (_25978_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  or _71590_ (_25979_, _25978_, _25977_);
  or _71591_ (_25980_, _25979_, _25976_);
  and _71592_ (_25981_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  and _71593_ (_25982_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or _71594_ (_25983_, _25982_, _25981_);
  and _71595_ (_25984_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  and _71596_ (_25985_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  or _71597_ (_25986_, _25985_, _25984_);
  or _71598_ (_25987_, _25986_, _25983_);
  or _71599_ (_25988_, _25987_, _25980_);
  and _71600_ (_25989_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and _71601_ (_25990_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  or _71602_ (_25991_, _25990_, _25989_);
  and _71603_ (_25992_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  and _71604_ (_25993_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or _71605_ (_25994_, _25993_, _25992_);
  or _71606_ (_25995_, _25994_, _25991_);
  and _71607_ (_25996_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and _71608_ (_25997_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  or _71609_ (_25998_, _25997_, _25996_);
  and _71610_ (_25999_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  and _71611_ (_26000_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or _71612_ (_26001_, _26000_, _25999_);
  or _71613_ (_26002_, _26001_, _25998_);
  or _71614_ (_26003_, _26002_, _25995_);
  or _71615_ (_26004_, _26003_, _25988_);
  or _71616_ (_26005_, _26004_, _25973_);
  or _71617_ (_26006_, _26005_, _25942_);
  and _71618_ (_26007_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and _71619_ (_26008_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  or _71620_ (_26009_, _26008_, _26007_);
  and _71621_ (_26010_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and _71622_ (_26011_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or _71623_ (_26012_, _26011_, _26010_);
  or _71624_ (_26013_, _26012_, _26009_);
  and _71625_ (_26014_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and _71626_ (_26015_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  or _71627_ (_26016_, _26015_, _26014_);
  and _71628_ (_26017_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  and _71629_ (_26018_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or _71630_ (_26019_, _26018_, _26017_);
  or _71631_ (_26020_, _26019_, _26016_);
  or _71632_ (_26021_, _26020_, _26013_);
  and _71633_ (_26022_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  and _71634_ (_26023_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or _71635_ (_26024_, _26023_, _26022_);
  and _71636_ (_26025_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and _71637_ (_26026_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  or _71638_ (_26027_, _26026_, _26025_);
  or _71639_ (_26028_, _26027_, _26024_);
  and _71640_ (_26029_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  and _71641_ (_26030_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or _71642_ (_26031_, _26030_, _26029_);
  and _71643_ (_26032_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and _71644_ (_26033_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  or _71645_ (_26034_, _26033_, _26032_);
  or _71646_ (_26035_, _26034_, _26031_);
  or _71647_ (_26036_, _26035_, _26028_);
  or _71648_ (_26037_, _26036_, _26021_);
  and _71649_ (_26038_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  and _71650_ (_26039_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or _71651_ (_26040_, _26039_, _26038_);
  and _71652_ (_26041_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  and _71653_ (_26042_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  or _71654_ (_26043_, _26042_, _26041_);
  or _71655_ (_26044_, _26043_, _26040_);
  and _71656_ (_26045_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  and _71657_ (_26046_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or _71658_ (_26047_, _26046_, _26045_);
  and _71659_ (_26048_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and _71660_ (_26049_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  or _71661_ (_26050_, _26049_, _26048_);
  or _71662_ (_26051_, _26050_, _26047_);
  or _71663_ (_26052_, _26051_, _26044_);
  and _71664_ (_26053_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and _71665_ (_26054_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  or _71666_ (_26055_, _26054_, _26053_);
  and _71667_ (_26056_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  and _71668_ (_26057_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or _71669_ (_26058_, _26057_, _26056_);
  or _71670_ (_26059_, _26058_, _26055_);
  and _71671_ (_26060_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and _71672_ (_26061_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  or _71673_ (_26062_, _26061_, _26060_);
  and _71674_ (_26063_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  and _71675_ (_26064_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or _71676_ (_26065_, _26064_, _26063_);
  or _71677_ (_26066_, _26065_, _26062_);
  or _71678_ (_26067_, _26066_, _26059_);
  or _71679_ (_26068_, _26067_, _26052_);
  or _71680_ (_26069_, _26068_, _26037_);
  and _71681_ (_26070_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and _71682_ (_26071_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and _71683_ (_26072_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or _71684_ (_26073_, _26072_, _26071_);
  or _71685_ (_26074_, _26073_, _26070_);
  and _71686_ (_26075_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and _71687_ (_26076_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or _71688_ (_26077_, _26076_, _26075_);
  and _71689_ (_26078_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and _71690_ (_26079_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or _71691_ (_26080_, _26079_, _26078_);
  or _71692_ (_26081_, _26080_, _26077_);
  or _71693_ (_26082_, _26081_, _26074_);
  and _71694_ (_26083_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _71695_ (_26084_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or _71696_ (_26085_, _26084_, _26083_);
  and _71697_ (_26086_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and _71698_ (_26087_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or _71699_ (_26088_, _26087_, _26086_);
  or _71700_ (_26089_, _26088_, _26085_);
  and _71701_ (_26090_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and _71702_ (_26091_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or _71703_ (_26092_, _26091_, _26090_);
  and _71704_ (_26093_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and _71705_ (_26094_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or _71706_ (_26095_, _26094_, _26093_);
  or _71707_ (_26096_, _26095_, _26092_);
  or _71708_ (_26097_, _26096_, _26089_);
  or _71709_ (_26098_, _26097_, _26082_);
  and _71710_ (_26099_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and _71711_ (_26100_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  or _71712_ (_26101_, _26100_, _26099_);
  and _71713_ (_26102_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  and _71714_ (_26103_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or _71715_ (_26104_, _26103_, _26102_);
  or _71716_ (_26105_, _26104_, _26101_);
  and _71717_ (_26106_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and _71718_ (_26107_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  or _71719_ (_26108_, _26107_, _26106_);
  and _71720_ (_26109_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and _71721_ (_26110_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or _71722_ (_26111_, _26110_, _26109_);
  or _71723_ (_26112_, _26111_, _26108_);
  or _71724_ (_26113_, _26112_, _26105_);
  and _71725_ (_26114_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  and _71726_ (_26115_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or _71727_ (_26116_, _26115_, _26114_);
  and _71728_ (_26117_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and _71729_ (_26118_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  or _71730_ (_26119_, _26118_, _26117_);
  or _71731_ (_26120_, _26119_, _26116_);
  and _71732_ (_26121_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  and _71733_ (_26122_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or _71734_ (_26123_, _26122_, _26121_);
  and _71735_ (_26124_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and _71736_ (_26125_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or _71737_ (_26126_, _26125_, _26124_);
  or _71738_ (_26127_, _26126_, _26123_);
  or _71739_ (_26128_, _26127_, _26120_);
  or _71740_ (_26129_, _26128_, _26113_);
  or _71741_ (_26130_, _26129_, _26098_);
  or _71742_ (_26131_, _26130_, _26069_);
  or _71743_ (_26132_, _26131_, _26006_);
  or _71744_ (_26133_, _26132_, _25879_);
  and _71745_ (_26134_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or _71746_ (_26135_, _26134_, _26133_);
  and _71747_ (_26136_, _26135_, _00006_);
  or _71748_ (_26137_, _26136_, _25624_);
  and _71749_ (_00003_[0], _26137_, _38997_);
  not _71750_ (_26138_, first_instr);
  nor _71751_ (_26139_, _15585_, _26138_);
  or _71752_ (_00002_, _26139_, rst);
  and _71753_ (_26140_, _15585_, iram_op1[7]);
  and _71754_ (_26141_, _15589_, iram_op1_reg[7]);
  or _71755_ (_26142_, _26141_, _26140_);
  and _71756_ (_00004_[7], _26142_, _38997_);
  and _71757_ (_26143_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _71758_ (_26144_, _21574_, acc_reg[7]);
  or _71759_ (_26145_, _26144_, _26143_);
  and _71760_ (_00000_[7], _26145_, _38997_);
  and _71761_ (_26146_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _71762_ (_26147_, cy_reg, _21574_);
  or _71763_ (_26148_, _26147_, _26146_);
  and _71764_ (_00001_, _26148_, _38997_);
  and _71765_ (_26149_, _18651_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _71766_ (_26150_, _26149_, _21683_);
  nor _71767_ (_26151_, _26150_, _16198_);
  nor _71768_ (_26152_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _71769_ (_26153_, _18646_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _71770_ (_26154_, _26153_, _26152_);
  nor _71771_ (_26155_, _26154_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _71772_ (_26156_, _26155_, _26151_);
  and _71773_ (_26157_, _26156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _71774_ (_26158_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _71775_ (_26159_, \oc8051_symbolic_cxrom1.regvalid [8], _16202_);
  nor _71776_ (_26160_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _71777_ (_26161_, _26160_, _26159_);
  and _71778_ (_26162_, _26161_, _26158_);
  and _71779_ (_26163_, _18663_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _71780_ (_26164_, _26163_, _21675_);
  and _71781_ (_26165_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], _16194_);
  and _71782_ (_26166_, _26165_, _26164_);
  or _71783_ (_26167_, _26166_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _71784_ (_26168_, _26167_, _26162_);
  nor _71785_ (_26169_, _26168_, _26157_);
  and _71786_ (_26170_, _18622_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _71787_ (_26171_, _26170_);
  nor _71788_ (_26172_, _21670_, _16198_);
  and _71789_ (_26173_, _26172_, _26171_);
  nor _71790_ (_26174_, \oc8051_symbolic_cxrom1.regvalid [11], _16202_);
  nor _71791_ (_26175_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _71792_ (_26176_, _26175_, _26174_);
  and _71793_ (_26177_, _26176_, _16198_);
  nor _71794_ (_26178_, _26177_, _26173_);
  nor _71795_ (_26179_, _26178_, _16194_);
  and _71796_ (_26180_, _18885_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _71797_ (_26181_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _71798_ (_26182_, _26181_, _26180_);
  and _71799_ (_26183_, _26182_, _26158_);
  and _71800_ (_26184_, _18630_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _71801_ (_26185_, _26184_, _21679_);
  and _71802_ (_26186_, _26185_, _26165_);
  or _71803_ (_26187_, _26186_, _16190_);
  or _71804_ (_26188_, _26187_, _26183_);
  nor _71805_ (_26189_, _26188_, _26179_);
  nor _71806_ (_26190_, _26189_, _26169_);
  nor _71807_ (_26191_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71808_ (_26192_, _20612_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71809_ (_26193_, _26192_, _26191_);
  and _71810_ (_26194_, _26193_, _26165_);
  not _71811_ (_26195_, _26194_);
  and _71812_ (_26196_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _71813_ (_26197_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71814_ (_26198_, _19705_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71815_ (_26199_, _26198_, _26197_);
  and _71816_ (_26200_, _26199_, _26196_);
  nor _71817_ (_26201_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71818_ (_26202_, _20606_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71819_ (_26203_, _26202_, _26201_);
  and _71820_ (_26204_, _26203_, _26158_);
  nor _71821_ (_26205_, _26204_, _26200_);
  and _71822_ (_26206_, _26205_, _26195_);
  nor _71823_ (_26207_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71824_ (_26208_, _20621_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71825_ (_26209_, _26208_, _26207_);
  and _71826_ (_26210_, _16198_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _71827_ (_26211_, _26210_, _26209_);
  nor _71828_ (_26212_, _26211_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _71829_ (_26213_, _26212_, _26206_);
  nor _71830_ (_26214_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71831_ (_26215_, _20318_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71832_ (_26216_, _26215_, _26214_);
  and _71833_ (_26217_, _26216_, _26165_);
  not _71834_ (_26218_, _26217_);
  nor _71835_ (_26219_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71836_ (_26220_, _20521_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71837_ (_26221_, _26220_, _26219_);
  and _71838_ (_26222_, _26221_, _26196_);
  nor _71839_ (_26223_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71840_ (_26224_, _19913_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71841_ (_26225_, _26224_, _26223_);
  and _71842_ (_26226_, _26225_, _26158_);
  nor _71843_ (_26227_, _26226_, _26222_);
  and _71844_ (_26228_, _26227_, _26218_);
  nor _71845_ (_26229_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71846_ (_26230_, _20116_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71847_ (_26231_, _26230_, _26229_);
  and _71848_ (_26232_, _26231_, _26210_);
  nor _71849_ (_26233_, _26232_, _16202_);
  and _71850_ (_26234_, _26233_, _26228_);
  nor _71851_ (_26235_, _26234_, _26213_);
  and _71852_ (_26236_, _26235_, _26190_);
  nor _71853_ (_26237_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71854_ (_26238_, _20704_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71855_ (_26239_, _26238_, _26237_);
  and _71856_ (_26240_, _26239_, _26165_);
  not _71857_ (_26241_, _26240_);
  nor _71858_ (_26242_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71859_ (_26243_, _19735_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71860_ (_26244_, _26243_, _26242_);
  and _71861_ (_26245_, _26244_, _26196_);
  nor _71862_ (_26246_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71863_ (_26247_, _20698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71864_ (_26248_, _26247_, _26246_);
  and _71865_ (_26249_, _26248_, _26158_);
  nor _71866_ (_26250_, _26249_, _26245_);
  and _71867_ (_26251_, _26250_, _26241_);
  nor _71868_ (_26252_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71869_ (_26253_, _20713_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71870_ (_26254_, _26253_, _26252_);
  and _71871_ (_26255_, _26254_, _26210_);
  nor _71872_ (_26256_, _26255_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _71873_ (_26257_, _26256_, _26251_);
  nor _71874_ (_26258_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71875_ (_26259_, _20346_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71876_ (_26260_, _26259_, _26258_);
  and _71877_ (_26261_, _26260_, _26165_);
  not _71878_ (_26262_, _26261_);
  nor _71879_ (_26263_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71880_ (_26264_, _20547_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71881_ (_26265_, _26264_, _26263_);
  and _71882_ (_26266_, _26265_, _26196_);
  nor _71883_ (_26267_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71884_ (_26268_, _19937_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71885_ (_26269_, _26268_, _26267_);
  and _71886_ (_26270_, _26269_, _26158_);
  nor _71887_ (_26271_, _26270_, _26266_);
  and _71888_ (_26272_, _26271_, _26262_);
  nor _71889_ (_26273_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71890_ (_26274_, _20142_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71891_ (_26275_, _26274_, _26273_);
  and _71892_ (_26276_, _26275_, _26210_);
  nor _71893_ (_26277_, _26276_, _16202_);
  and _71894_ (_26278_, _26277_, _26272_);
  nor _71895_ (_26279_, _26278_, _26257_);
  and _71896_ (_26280_, _26279_, _26190_);
  nor _71897_ (_26281_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71898_ (_26282_, _20658_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71899_ (_26283_, _26282_, _26281_);
  and _71900_ (_26284_, _26283_, _26165_);
  not _71901_ (_26285_, _26284_);
  nor _71902_ (_26286_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71903_ (_26287_, _19721_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71904_ (_26288_, _26287_, _26286_);
  and _71905_ (_26289_, _26288_, _26196_);
  nor _71906_ (_26290_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71907_ (_26291_, _20652_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71908_ (_26292_, _26291_, _26290_);
  and _71909_ (_26293_, _26292_, _26158_);
  nor _71910_ (_26294_, _26293_, _26289_);
  and _71911_ (_26295_, _26294_, _26285_);
  nor _71912_ (_26296_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71913_ (_26297_, _20667_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71914_ (_26298_, _26297_, _26296_);
  and _71915_ (_26299_, _26298_, _26210_);
  nor _71916_ (_26300_, _26299_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _71917_ (_26301_, _26300_, _26295_);
  nor _71918_ (_26302_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71919_ (_26303_, _20334_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71920_ (_26304_, _26303_, _26302_);
  and _71921_ (_26305_, _26304_, _26165_);
  not _71922_ (_26306_, _26305_);
  nor _71923_ (_26307_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71924_ (_26308_, _20534_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71925_ (_26309_, _26308_, _26307_);
  and _71926_ (_26310_, _26309_, _26196_);
  nor _71927_ (_26311_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71928_ (_26312_, _19925_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71929_ (_26313_, _26312_, _26311_);
  and _71930_ (_26314_, _26313_, _26158_);
  nor _71931_ (_26315_, _26314_, _26310_);
  and _71932_ (_26316_, _26315_, _26306_);
  nor _71933_ (_26317_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71934_ (_26318_, _20127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71935_ (_26319_, _26318_, _26317_);
  and _71936_ (_26320_, _26319_, _26210_);
  nor _71937_ (_26321_, _26320_, _16202_);
  and _71938_ (_26322_, _26321_, _26316_);
  nor _71939_ (_26323_, _26322_, _26301_);
  nor _71940_ (_26324_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71941_ (_26325_, _20750_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71942_ (_26326_, _26325_, _26324_);
  and _71943_ (_26327_, _26326_, _26165_);
  not _71944_ (_26328_, _26327_);
  nor _71945_ (_26329_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71946_ (_26330_, _19745_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71947_ (_26331_, _26330_, _26329_);
  and _71948_ (_26332_, _26331_, _26196_);
  nor _71949_ (_26333_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71950_ (_26334_, _20744_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71951_ (_26335_, _26334_, _26333_);
  and _71952_ (_26336_, _26335_, _26158_);
  nor _71953_ (_26337_, _26336_, _26332_);
  and _71954_ (_26338_, _26337_, _26328_);
  nor _71955_ (_26339_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71956_ (_26340_, _20759_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71957_ (_26341_, _26340_, _26339_);
  and _71958_ (_26342_, _26341_, _26210_);
  nor _71959_ (_26343_, _26342_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _71960_ (_26344_, _26343_, _26338_);
  nor _71961_ (_26345_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71962_ (_26346_, _20359_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71963_ (_26347_, _26346_, _26345_);
  and _71964_ (_26348_, _26347_, _26165_);
  not _71965_ (_26349_, _26348_);
  nor _71966_ (_26350_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71967_ (_26351_, _20559_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71968_ (_26352_, _26351_, _26350_);
  and _71969_ (_26353_, _26352_, _26196_);
  nor _71970_ (_26354_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71971_ (_26355_, _19951_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71972_ (_26356_, _26355_, _26354_);
  and _71973_ (_26357_, _26356_, _26158_);
  nor _71974_ (_26358_, _26357_, _26353_);
  and _71975_ (_26359_, _26358_, _26349_);
  nor _71976_ (_26360_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71977_ (_26361_, _20154_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71978_ (_26362_, _26361_, _26360_);
  and _71979_ (_26363_, _26362_, _26210_);
  nor _71980_ (_26364_, _26363_, _16202_);
  and _71981_ (_26365_, _26364_, _26359_);
  nor _71982_ (_26366_, _26365_, _26344_);
  nor _71983_ (_26367_, _26366_, _26323_);
  and _71984_ (_26368_, _26367_, _26280_);
  and _71985_ (_26369_, _26368_, _26236_);
  nor _71986_ (_26370_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71987_ (_26371_, _20888_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71988_ (_26372_, _26371_, _26370_);
  and _71989_ (_26373_, _26372_, _26165_);
  not _71990_ (_26374_, _26373_);
  nor _71991_ (_26375_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71992_ (_26376_, _19782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71993_ (_26377_, _26376_, _26375_);
  and _71994_ (_26378_, _26377_, _26196_);
  nor _71995_ (_26379_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _71996_ (_26380_, _20882_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _71997_ (_26381_, _26380_, _26379_);
  and _71998_ (_26382_, _26381_, _26158_);
  nor _71999_ (_26383_, _26382_, _26378_);
  and _72000_ (_26384_, _26383_, _26374_);
  nor _72001_ (_26385_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72002_ (_26386_, _20897_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72003_ (_26387_, _26386_, _26385_);
  and _72004_ (_26388_, _26387_, _26210_);
  nor _72005_ (_26389_, _26388_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _72006_ (_26390_, _26389_, _26384_);
  nor _72007_ (_26391_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72008_ (_26392_, _20395_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72009_ (_26393_, _26392_, _26391_);
  and _72010_ (_26394_, _26393_, _26165_);
  not _72011_ (_26395_, _26394_);
  nor _72012_ (_26396_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72013_ (_26397_, _20593_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72014_ (_26398_, _26397_, _26396_);
  and _72015_ (_26399_, _26398_, _26196_);
  nor _72016_ (_26400_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72017_ (_26401_, _19988_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72018_ (_26402_, _26401_, _26400_);
  and _72019_ (_26403_, _26402_, _26158_);
  nor _72020_ (_26404_, _26403_, _26399_);
  and _72021_ (_26405_, _26404_, _26395_);
  nor _72022_ (_26406_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72023_ (_26407_, _20190_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72024_ (_26408_, _26407_, _26406_);
  and _72025_ (_26409_, _26408_, _26210_);
  nor _72026_ (_26410_, _26409_, _16202_);
  and _72027_ (_26411_, _26410_, _26405_);
  nor _72028_ (_26412_, _26411_, _26390_);
  and _72029_ (_26413_, _26412_, _26190_);
  nor _72030_ (_26414_, \oc8051_symbolic_cxrom1.regarray[4] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72031_ (_26415_, _18457_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72032_ (_26416_, _26415_, _26414_);
  and _72033_ (_26417_, _26416_, _26165_);
  not _72034_ (_26418_, _26417_);
  nor _72035_ (_26419_, \oc8051_symbolic_cxrom1.regarray[6] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72036_ (_26420_, _18451_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72037_ (_26421_, _26420_, _26419_);
  and _72038_ (_26422_, _26421_, _26196_);
  nor _72039_ (_26423_, \oc8051_symbolic_cxrom1.regarray[0] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72040_ (_26424_, _18443_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72041_ (_26425_, _26424_, _26423_);
  and _72042_ (_26426_, _26425_, _26158_);
  nor _72043_ (_26427_, _26426_, _26422_);
  and _72044_ (_26428_, _26427_, _26418_);
  nor _72045_ (_26429_, \oc8051_symbolic_cxrom1.regarray[2] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72046_ (_26430_, _18462_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72047_ (_26431_, _26430_, _26429_);
  and _72048_ (_26432_, _26431_, _26210_);
  nor _72049_ (_26433_, _26432_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _72050_ (_26434_, _26433_, _26428_);
  nor _72051_ (_26435_, \oc8051_symbolic_cxrom1.regarray[12] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72052_ (_26436_, _18478_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72053_ (_26437_, _26436_, _26435_);
  and _72054_ (_26438_, _26437_, _26165_);
  not _72055_ (_26439_, _26438_);
  nor _72056_ (_26440_, \oc8051_symbolic_cxrom1.regarray[14] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72057_ (_26441_, _18483_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72058_ (_26442_, _26441_, _26440_);
  and _72059_ (_26443_, _26442_, _26196_);
  nor _72060_ (_26444_, \oc8051_symbolic_cxrom1.regarray[8] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72061_ (_26445_, _18472_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72062_ (_26446_, _26445_, _26444_);
  and _72063_ (_26447_, _26446_, _26158_);
  nor _72064_ (_26448_, _26447_, _26443_);
  and _72065_ (_26449_, _26448_, _26439_);
  nor _72066_ (_26450_, \oc8051_symbolic_cxrom1.regarray[10] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72067_ (_26451_, _18489_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72068_ (_26452_, _26451_, _26450_);
  and _72069_ (_26453_, _26452_, _26210_);
  nor _72070_ (_26454_, _26453_, _16202_);
  and _72071_ (_26455_, _26454_, _26449_);
  nor _72072_ (_26456_, _26455_, _26434_);
  and _72073_ (_26457_, _26456_, _26190_);
  nor _72074_ (_26458_, _26457_, _26413_);
  nor _72075_ (_26459_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72076_ (_26460_, _20796_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72077_ (_26461_, _26460_, _26459_);
  and _72078_ (_26462_, _26461_, _26165_);
  not _72079_ (_26463_, _26462_);
  nor _72080_ (_26464_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72081_ (_26465_, _19759_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72082_ (_26466_, _26465_, _26464_);
  and _72083_ (_26467_, _26466_, _26196_);
  nor _72084_ (_26468_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72085_ (_26469_, _20790_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72086_ (_26470_, _26469_, _26468_);
  and _72087_ (_26471_, _26470_, _26158_);
  nor _72088_ (_26472_, _26471_, _26467_);
  and _72089_ (_26473_, _26472_, _26463_);
  nor _72090_ (_26474_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72091_ (_26475_, _20805_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72092_ (_26476_, _26475_, _26474_);
  and _72093_ (_26477_, _26476_, _26210_);
  nor _72094_ (_26478_, _26477_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _72095_ (_26479_, _26478_, _26473_);
  nor _72096_ (_26480_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72097_ (_26481_, _20372_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72098_ (_26482_, _26481_, _26480_);
  and _72099_ (_26483_, _26482_, _26165_);
  not _72100_ (_26484_, _26483_);
  nor _72101_ (_26485_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72102_ (_26486_, _20571_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72103_ (_26487_, _26486_, _26485_);
  and _72104_ (_26488_, _26487_, _26196_);
  nor _72105_ (_26489_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72106_ (_26490_, _19963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72107_ (_26491_, _26490_, _26489_);
  and _72108_ (_26492_, _26491_, _26158_);
  nor _72109_ (_26493_, _26492_, _26488_);
  and _72110_ (_26494_, _26493_, _26484_);
  nor _72111_ (_26495_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72112_ (_26496_, _20165_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72113_ (_26497_, _26496_, _26495_);
  and _72114_ (_26498_, _26497_, _26210_);
  nor _72115_ (_26499_, _26498_, _16202_);
  and _72116_ (_26500_, _26499_, _26494_);
  nor _72117_ (_26501_, _26500_, _26479_);
  and _72118_ (_26502_, _26501_, _26190_);
  nor _72119_ (_26503_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72120_ (_26504_, _20842_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72121_ (_26505_, _26504_, _26503_);
  and _72122_ (_26506_, _26505_, _26165_);
  not _72123_ (_26507_, _26506_);
  nor _72124_ (_26508_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72125_ (_26509_, _19770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72126_ (_26510_, _26509_, _26508_);
  and _72127_ (_26511_, _26510_, _26196_);
  nor _72128_ (_26512_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72129_ (_26513_, _20836_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72130_ (_26514_, _26513_, _26512_);
  and _72131_ (_26515_, _26514_, _26158_);
  nor _72132_ (_26516_, _26515_, _26511_);
  and _72133_ (_26517_, _26516_, _26507_);
  nor _72134_ (_26518_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72135_ (_26519_, _20851_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72136_ (_26520_, _26519_, _26518_);
  and _72137_ (_26521_, _26520_, _26210_);
  nor _72138_ (_26522_, _26521_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _72139_ (_26523_, _26522_, _26517_);
  nor _72140_ (_26524_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72141_ (_26525_, _20382_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72142_ (_26526_, _26525_, _26524_);
  and _72143_ (_26527_, _26526_, _26165_);
  not _72144_ (_26528_, _26527_);
  nor _72145_ (_26529_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72146_ (_26530_, _20584_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72147_ (_26531_, _26530_, _26529_);
  and _72148_ (_26532_, _26531_, _26196_);
  nor _72149_ (_26533_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72150_ (_26534_, _19975_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72151_ (_26535_, _26534_, _26533_);
  and _72152_ (_26536_, _26535_, _26158_);
  nor _72153_ (_26537_, _26536_, _26532_);
  and _72154_ (_26538_, _26537_, _26528_);
  nor _72155_ (_26539_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _72156_ (_26540_, _20178_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72157_ (_26541_, _26540_, _26539_);
  and _72158_ (_26542_, _26541_, _26210_);
  nor _72159_ (_26543_, _26542_, _16202_);
  and _72160_ (_26544_, _26543_, _26538_);
  nor _72161_ (_26545_, _26544_, _26523_);
  and _72162_ (_26546_, _26545_, _26190_);
  nor _72163_ (_26547_, _26546_, _26502_);
  and _72164_ (_26548_, _26547_, _26458_);
  and _72165_ (_26549_, _26548_, _38997_);
  and _72166_ (_00008_, _26549_, _26369_);
  not _72167_ (_26550_, _26236_);
  and _72168_ (_26551_, _26368_, _26550_);
  and _72169_ (_00007_, _26551_, _26549_);
  or _72170_ (_26552_, _21983_, _15589_);
  or _72171_ (_26553_, _15585_, op1_out_r[7]);
  and _72172_ (_26554_, _26553_, _38997_);
  and _72173_ (_00005_[7], _26554_, _26552_);
  and _72174_ (_26555_, _15589_, iram_op1[7]);
  and _72175_ (_26556_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  and _72176_ (_26557_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or _72177_ (_26558_, _26557_, _26556_);
  and _72178_ (_26559_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and _72179_ (_26560_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  or _72180_ (_26561_, _26560_, _26559_);
  or _72181_ (_26562_, _26561_, _26558_);
  and _72182_ (_26563_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  and _72183_ (_26564_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or _72184_ (_26565_, _26564_, _26563_);
  and _72185_ (_26566_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and _72186_ (_26567_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  or _72187_ (_26568_, _26567_, _26566_);
  or _72188_ (_26569_, _26568_, _26565_);
  or _72189_ (_26570_, _26569_, _26562_);
  and _72190_ (_26571_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and _72191_ (_26572_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  or _72192_ (_26573_, _26572_, _26571_);
  and _72193_ (_26574_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  and _72194_ (_26575_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or _72195_ (_26576_, _26575_, _26574_);
  or _72196_ (_26577_, _26576_, _26573_);
  and _72197_ (_26578_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and _72198_ (_26579_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  or _72199_ (_26580_, _26579_, _26578_);
  and _72200_ (_26581_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  and _72201_ (_26582_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  or _72202_ (_26583_, _26582_, _26581_);
  or _72203_ (_26584_, _26583_, _26580_);
  or _72204_ (_26585_, _26584_, _26577_);
  or _72205_ (_26586_, _26585_, _26570_);
  and _72206_ (_26587_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and _72207_ (_26588_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or _72208_ (_26589_, _26588_, _26587_);
  and _72209_ (_26590_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  and _72210_ (_26591_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or _72211_ (_26592_, _26591_, _26590_);
  or _72212_ (_26593_, _26592_, _26589_);
  and _72213_ (_26594_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and _72214_ (_26595_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  or _72215_ (_26596_, _26595_, _26594_);
  and _72216_ (_26597_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  and _72217_ (_26598_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or _72218_ (_26599_, _26598_, _26597_);
  or _72219_ (_26600_, _26599_, _26596_);
  or _72220_ (_26601_, _26600_, _26593_);
  and _72221_ (_26602_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  and _72222_ (_26603_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or _72223_ (_26604_, _26603_, _26602_);
  and _72224_ (_26605_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and _72225_ (_26606_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or _72226_ (_26607_, _26606_, _26605_);
  or _72227_ (_26608_, _26607_, _26604_);
  and _72228_ (_26609_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  and _72229_ (_26610_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or _72230_ (_26611_, _26610_, _26609_);
  and _72231_ (_26612_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  and _72232_ (_26613_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or _72233_ (_26614_, _26613_, _26612_);
  or _72234_ (_26615_, _26614_, _26611_);
  or _72235_ (_26616_, _26615_, _26608_);
  or _72236_ (_26617_, _26616_, _26601_);
  or _72237_ (_26618_, _26617_, _26586_);
  and _72238_ (_26619_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and _72239_ (_26620_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  or _72240_ (_26621_, _26620_, _26619_);
  and _72241_ (_26622_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  and _72242_ (_26623_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or _72243_ (_26624_, _26623_, _26622_);
  or _72244_ (_26625_, _26624_, _26621_);
  and _72245_ (_26626_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and _72246_ (_26627_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  or _72247_ (_26628_, _26627_, _26626_);
  and _72248_ (_26629_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  and _72249_ (_26630_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or _72250_ (_26631_, _26630_, _26629_);
  or _72251_ (_26632_, _26631_, _26628_);
  or _72252_ (_26633_, _26632_, _26625_);
  and _72253_ (_26634_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  and _72254_ (_26635_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or _72255_ (_26636_, _26635_, _26634_);
  and _72256_ (_26637_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  and _72257_ (_26638_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or _72258_ (_26639_, _26638_, _26637_);
  or _72259_ (_26640_, _26639_, _26636_);
  and _72260_ (_26641_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  and _72261_ (_26642_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or _72262_ (_26643_, _26642_, _26641_);
  and _72263_ (_26644_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and _72264_ (_26645_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  or _72265_ (_26646_, _26645_, _26644_);
  or _72266_ (_26647_, _26646_, _26643_);
  or _72267_ (_26648_, _26647_, _26640_);
  or _72268_ (_26649_, _26648_, _26633_);
  and _72269_ (_26650_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and _72270_ (_26651_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  or _72271_ (_26652_, _26651_, _26650_);
  and _72272_ (_26653_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  and _72273_ (_26654_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or _72274_ (_26655_, _26654_, _26653_);
  or _72275_ (_26656_, _26655_, _26652_);
  and _72276_ (_26657_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and _72277_ (_26658_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  or _72278_ (_26659_, _26658_, _26657_);
  and _72279_ (_26660_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and _72280_ (_26661_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or _72281_ (_26662_, _26661_, _26660_);
  or _72282_ (_26663_, _26662_, _26659_);
  or _72283_ (_26664_, _26663_, _26656_);
  and _72284_ (_26665_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  and _72285_ (_26666_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or _72286_ (_26667_, _26666_, _26665_);
  and _72287_ (_26668_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and _72288_ (_26669_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  or _72289_ (_26670_, _26669_, _26668_);
  or _72290_ (_26671_, _26670_, _26667_);
  and _72291_ (_26672_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  and _72292_ (_26673_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or _72293_ (_26674_, _26673_, _26672_);
  and _72294_ (_26675_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and _72295_ (_26676_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  or _72296_ (_26677_, _26676_, _26675_);
  or _72297_ (_26678_, _26677_, _26674_);
  or _72298_ (_26679_, _26678_, _26671_);
  or _72299_ (_26680_, _26679_, _26664_);
  or _72300_ (_26681_, _26680_, _26649_);
  or _72301_ (_26682_, _26681_, _26618_);
  and _72302_ (_26683_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  and _72303_ (_26684_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or _72304_ (_26685_, _26684_, _26683_);
  and _72305_ (_26686_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and _72306_ (_26687_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or _72307_ (_26688_, _26687_, _26686_);
  or _72308_ (_26689_, _26688_, _26685_);
  and _72309_ (_26690_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  and _72310_ (_26691_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or _72311_ (_26692_, _26691_, _26690_);
  and _72312_ (_26693_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and _72313_ (_26694_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  or _72314_ (_26695_, _26694_, _26693_);
  or _72315_ (_26696_, _26695_, _26692_);
  or _72316_ (_26697_, _26696_, _26689_);
  and _72317_ (_26698_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and _72318_ (_26699_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or _72319_ (_26700_, _26699_, _26698_);
  and _72320_ (_26701_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  and _72321_ (_26702_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or _72322_ (_26703_, _26702_, _26701_);
  or _72323_ (_26704_, _26703_, _26700_);
  and _72324_ (_26705_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and _72325_ (_26706_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or _72326_ (_26707_, _26706_, _26705_);
  and _72327_ (_26708_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  and _72328_ (_26709_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or _72329_ (_26710_, _26709_, _26708_);
  or _72330_ (_26711_, _26710_, _26707_);
  or _72331_ (_26712_, _26711_, _26704_);
  or _72332_ (_26713_, _26712_, _26697_);
  and _72333_ (_26714_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  and _72334_ (_26715_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or _72335_ (_26716_, _26715_, _26714_);
  and _72336_ (_26717_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and _72337_ (_26718_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  or _72338_ (_26719_, _26718_, _26717_);
  or _72339_ (_26720_, _26719_, _26716_);
  and _72340_ (_26721_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  and _72341_ (_26722_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or _72342_ (_26723_, _26722_, _26721_);
  and _72343_ (_26724_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and _72344_ (_26725_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or _72345_ (_26726_, _26725_, _26724_);
  or _72346_ (_26727_, _26726_, _26723_);
  or _72347_ (_26728_, _26727_, _26720_);
  and _72348_ (_26729_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and _72349_ (_26730_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  or _72350_ (_26731_, _26730_, _26729_);
  and _72351_ (_26732_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  and _72352_ (_26733_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or _72353_ (_26734_, _26733_, _26732_);
  or _72354_ (_26735_, _26734_, _26731_);
  and _72355_ (_26736_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and _72356_ (_26737_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  or _72357_ (_26738_, _26737_, _26736_);
  and _72358_ (_26739_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  and _72359_ (_26740_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or _72360_ (_26741_, _26740_, _26739_);
  or _72361_ (_26742_, _26741_, _26738_);
  or _72362_ (_26743_, _26742_, _26735_);
  or _72363_ (_26744_, _26743_, _26728_);
  or _72364_ (_26745_, _26744_, _26713_);
  and _72365_ (_26746_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and _72366_ (_26747_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  or _72367_ (_26748_, _26747_, _26746_);
  and _72368_ (_26749_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  and _72369_ (_26750_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or _72370_ (_26751_, _26750_, _26749_);
  or _72371_ (_26752_, _26751_, _26748_);
  and _72372_ (_26753_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and _72373_ (_26754_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  or _72374_ (_26755_, _26754_, _26753_);
  and _72375_ (_26756_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and _72376_ (_26757_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or _72377_ (_26758_, _26757_, _26756_);
  or _72378_ (_26759_, _26758_, _26755_);
  or _72379_ (_26760_, _26759_, _26752_);
  and _72380_ (_26761_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  and _72381_ (_26762_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or _72382_ (_26763_, _26762_, _26761_);
  and _72383_ (_26764_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and _72384_ (_26765_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  or _72385_ (_26766_, _26765_, _26764_);
  or _72386_ (_26767_, _26766_, _26763_);
  and _72387_ (_26768_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and _72388_ (_26769_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  or _72389_ (_26770_, _26769_, _26768_);
  and _72390_ (_26771_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  and _72391_ (_26772_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or _72392_ (_26773_, _26772_, _26771_);
  or _72393_ (_26774_, _26773_, _26770_);
  or _72394_ (_26775_, _26774_, _26767_);
  or _72395_ (_26776_, _26775_, _26760_);
  and _72396_ (_26777_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  and _72397_ (_26778_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or _72398_ (_26779_, _26778_, _26777_);
  and _72399_ (_26780_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and _72400_ (_26781_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  or _72401_ (_26782_, _26781_, _26780_);
  or _72402_ (_26783_, _26782_, _26779_);
  and _72403_ (_26784_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  and _72404_ (_26785_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or _72405_ (_26786_, _26785_, _26784_);
  and _72406_ (_26787_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  and _72407_ (_26788_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  or _72408_ (_26789_, _26788_, _26787_);
  or _72409_ (_26790_, _26789_, _26786_);
  or _72410_ (_26791_, _26790_, _26783_);
  and _72411_ (_26792_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and _72412_ (_26793_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  or _72413_ (_26794_, _26793_, _26792_);
  and _72414_ (_26795_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  and _72415_ (_26796_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or _72416_ (_26797_, _26796_, _26795_);
  or _72417_ (_26798_, _26797_, _26794_);
  and _72418_ (_26799_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and _72419_ (_26800_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  or _72420_ (_26801_, _26800_, _26799_);
  and _72421_ (_26802_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  and _72422_ (_26803_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or _72423_ (_26804_, _26803_, _26802_);
  or _72424_ (_26805_, _26804_, _26801_);
  or _72425_ (_26806_, _26805_, _26798_);
  or _72426_ (_26807_, _26806_, _26791_);
  or _72427_ (_26808_, _26807_, _26776_);
  or _72428_ (_26809_, _26808_, _26745_);
  or _72429_ (_26810_, _26809_, _26682_);
  and _72430_ (_26811_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and _72431_ (_26812_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  or _72432_ (_26813_, _26812_, _26811_);
  and _72433_ (_26814_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  and _72434_ (_26815_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or _72435_ (_26816_, _26815_, _26814_);
  or _72436_ (_26817_, _26816_, _26813_);
  and _72437_ (_26818_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and _72438_ (_26819_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  or _72439_ (_26820_, _26819_, _26818_);
  and _72440_ (_26821_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and _72441_ (_26822_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or _72442_ (_26823_, _26822_, _26821_);
  or _72443_ (_26824_, _26823_, _26820_);
  or _72444_ (_26825_, _26824_, _26817_);
  and _72445_ (_26826_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  and _72446_ (_26827_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or _72447_ (_26828_, _26827_, _26826_);
  and _72448_ (_26829_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and _72449_ (_26830_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  or _72450_ (_26831_, _26830_, _26829_);
  or _72451_ (_26832_, _26831_, _26828_);
  and _72452_ (_26833_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  and _72453_ (_26834_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or _72454_ (_26835_, _26834_, _26833_);
  and _72455_ (_26836_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and _72456_ (_26837_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  or _72457_ (_26838_, _26837_, _26836_);
  or _72458_ (_26839_, _26838_, _26835_);
  or _72459_ (_26840_, _26839_, _26832_);
  or _72460_ (_26841_, _26840_, _26825_);
  and _72461_ (_26842_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  and _72462_ (_26843_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or _72463_ (_26844_, _26843_, _26842_);
  and _72464_ (_26845_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and _72465_ (_26846_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or _72466_ (_26847_, _26846_, _26845_);
  or _72467_ (_26848_, _26847_, _26844_);
  and _72468_ (_26849_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  and _72469_ (_26850_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or _72470_ (_26851_, _26850_, _26849_);
  and _72471_ (_26852_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  and _72472_ (_26853_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or _72473_ (_26854_, _26853_, _26852_);
  or _72474_ (_26855_, _26854_, _26851_);
  or _72475_ (_26856_, _26855_, _26848_);
  and _72476_ (_26857_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and _72477_ (_26858_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or _72478_ (_26859_, _26858_, _26857_);
  and _72479_ (_26860_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  and _72480_ (_26861_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or _72481_ (_26862_, _26861_, _26860_);
  or _72482_ (_26863_, _26862_, _26859_);
  and _72483_ (_26864_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and _72484_ (_26865_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or _72485_ (_26866_, _26865_, _26864_);
  and _72486_ (_26867_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  and _72487_ (_26868_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or _72488_ (_26869_, _26868_, _26867_);
  or _72489_ (_26870_, _26869_, _26866_);
  or _72490_ (_26871_, _26870_, _26863_);
  or _72491_ (_26872_, _26871_, _26856_);
  or _72492_ (_26873_, _26872_, _26841_);
  and _72493_ (_26874_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  and _72494_ (_26875_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or _72495_ (_26876_, _26875_, _26874_);
  and _72496_ (_26877_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and _72497_ (_26878_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or _72498_ (_26879_, _26878_, _26877_);
  or _72499_ (_26880_, _26879_, _26876_);
  and _72500_ (_26881_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  and _72501_ (_26882_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or _72502_ (_26883_, _26882_, _26881_);
  and _72503_ (_26884_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and _72504_ (_26885_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or _72505_ (_26886_, _26885_, _26884_);
  or _72506_ (_26887_, _26886_, _26883_);
  or _72507_ (_26888_, _26887_, _26880_);
  and _72508_ (_26889_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and _72509_ (_26890_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or _72510_ (_26891_, _26890_, _26889_);
  and _72511_ (_26892_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  and _72512_ (_26893_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or _72513_ (_26894_, _26893_, _26892_);
  or _72514_ (_26895_, _26894_, _26891_);
  and _72515_ (_26896_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and _72516_ (_26897_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  or _72517_ (_26898_, _26897_, _26896_);
  and _72518_ (_26899_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  and _72519_ (_26900_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  or _72520_ (_26901_, _26900_, _26899_);
  or _72521_ (_26902_, _26901_, _26898_);
  or _72522_ (_26903_, _26902_, _26895_);
  or _72523_ (_26904_, _26903_, _26888_);
  and _72524_ (_26905_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and _72525_ (_26906_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  or _72526_ (_26907_, _26906_, _26905_);
  and _72527_ (_26908_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  and _72528_ (_26909_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or _72529_ (_26910_, _26909_, _26908_);
  or _72530_ (_26911_, _26910_, _26907_);
  and _72531_ (_26912_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and _72532_ (_26913_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or _72533_ (_26914_, _26913_, _26912_);
  and _72534_ (_26915_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  and _72535_ (_26916_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or _72536_ (_26917_, _26916_, _26915_);
  or _72537_ (_26918_, _26917_, _26914_);
  or _72538_ (_26919_, _26918_, _26911_);
  and _72539_ (_26920_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  and _72540_ (_26921_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or _72541_ (_26922_, _26921_, _26920_);
  and _72542_ (_26923_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and _72543_ (_26924_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or _72544_ (_26925_, _26924_, _26923_);
  or _72545_ (_26926_, _26925_, _26922_);
  and _72546_ (_26927_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  and _72547_ (_26928_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or _72548_ (_26929_, _26928_, _26927_);
  and _72549_ (_26930_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and _72550_ (_26931_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or _72551_ (_26932_, _26931_, _26930_);
  or _72552_ (_26933_, _26932_, _26929_);
  or _72553_ (_26934_, _26933_, _26926_);
  or _72554_ (_26935_, _26934_, _26919_);
  or _72555_ (_26936_, _26935_, _26904_);
  or _72556_ (_26937_, _26936_, _26873_);
  and _72557_ (_26938_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and _72558_ (_26939_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  or _72559_ (_26940_, _26939_, _26938_);
  and _72560_ (_26941_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  and _72561_ (_26942_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  or _72562_ (_26943_, _26942_, _26941_);
  or _72563_ (_26944_, _26943_, _26940_);
  and _72564_ (_26945_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and _72565_ (_26946_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  or _72566_ (_26947_, _26946_, _26945_);
  and _72567_ (_26948_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  and _72568_ (_26949_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or _72569_ (_26950_, _26949_, _26948_);
  or _72570_ (_26951_, _26950_, _26947_);
  or _72571_ (_26952_, _26951_, _26944_);
  and _72572_ (_26953_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  and _72573_ (_26954_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or _72574_ (_26955_, _26954_, _26953_);
  and _72575_ (_26956_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and _72576_ (_26957_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or _72577_ (_26958_, _26957_, _26956_);
  or _72578_ (_26959_, _26958_, _26955_);
  and _72579_ (_26960_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and _72580_ (_26961_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or _72581_ (_26962_, _26961_, _26960_);
  and _72582_ (_26963_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  and _72583_ (_26964_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or _72584_ (_26965_, _26964_, _26963_);
  or _72585_ (_26966_, _26965_, _26962_);
  or _72586_ (_26967_, _26966_, _26959_);
  or _72587_ (_26968_, _26967_, _26952_);
  and _72588_ (_26969_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  and _72589_ (_26970_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or _72590_ (_26971_, _26970_, _26969_);
  and _72591_ (_26972_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and _72592_ (_26973_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or _72593_ (_26974_, _26973_, _26972_);
  or _72594_ (_26975_, _26974_, _26971_);
  and _72595_ (_26976_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  and _72596_ (_26977_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or _72597_ (_26978_, _26977_, _26976_);
  and _72598_ (_26979_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and _72599_ (_26980_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or _72600_ (_26981_, _26980_, _26979_);
  or _72601_ (_26982_, _26981_, _26978_);
  or _72602_ (_26983_, _26982_, _26975_);
  and _72603_ (_26984_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  and _72604_ (_26985_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or _72605_ (_26986_, _26985_, _26984_);
  and _72606_ (_26987_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and _72607_ (_26988_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  or _72608_ (_26989_, _26988_, _26987_);
  or _72609_ (_26990_, _26989_, _26986_);
  and _72610_ (_26991_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and _72611_ (_26992_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  or _72612_ (_26993_, _26992_, _26991_);
  and _72613_ (_26994_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  and _72614_ (_26995_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or _72615_ (_26996_, _26995_, _26994_);
  or _72616_ (_26997_, _26996_, _26993_);
  or _72617_ (_26998_, _26997_, _26990_);
  or _72618_ (_26999_, _26998_, _26983_);
  or _72619_ (_27000_, _26999_, _26968_);
  and _72620_ (_27001_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  and _72621_ (_27002_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or _72622_ (_27003_, _27002_, _27001_);
  and _72623_ (_27004_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and _72624_ (_27005_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or _72625_ (_27006_, _27005_, _27004_);
  or _72626_ (_27007_, _27006_, _27003_);
  and _72627_ (_27008_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  and _72628_ (_27009_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or _72629_ (_27010_, _27009_, _27008_);
  and _72630_ (_27011_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and _72631_ (_27012_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or _72632_ (_27013_, _27012_, _27011_);
  or _72633_ (_27014_, _27013_, _27010_);
  or _72634_ (_27015_, _27014_, _27007_);
  and _72635_ (_27016_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and _72636_ (_27017_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  or _72637_ (_27018_, _27017_, _27016_);
  and _72638_ (_27019_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and _72639_ (_27020_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or _72640_ (_27021_, _27020_, _27019_);
  or _72641_ (_27022_, _27021_, _27018_);
  and _72642_ (_27023_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and _72643_ (_27024_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  or _72644_ (_27025_, _27024_, _27023_);
  and _72645_ (_27026_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  and _72646_ (_27027_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or _72647_ (_27028_, _27027_, _27026_);
  or _72648_ (_27029_, _27028_, _27025_);
  or _72649_ (_27030_, _27029_, _27022_);
  or _72650_ (_27031_, _27030_, _27015_);
  and _72651_ (_27032_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and _72652_ (_27033_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and _72653_ (_27034_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and _72654_ (_27035_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or _72655_ (_27036_, _27035_, _27034_);
  or _72656_ (_27037_, _27036_, _27033_);
  or _72657_ (_27038_, _27037_, _27032_);
  and _72658_ (_27039_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and _72659_ (_27040_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and _72660_ (_27041_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _72661_ (_27042_, _27041_, _27040_);
  or _72662_ (_27043_, _27042_, _27039_);
  or _72663_ (_27044_, _27043_, _27038_);
  and _72664_ (_27045_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and _72665_ (_27046_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or _72666_ (_27047_, _27046_, _27045_);
  and _72667_ (_27048_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and _72668_ (_27049_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or _72669_ (_27050_, _27049_, _27048_);
  or _72670_ (_27051_, _27050_, _27047_);
  and _72671_ (_27052_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and _72672_ (_27053_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or _72673_ (_27054_, _27053_, _27052_);
  and _72674_ (_27055_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and _72675_ (_27056_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or _72676_ (_27057_, _27056_, _27055_);
  or _72677_ (_27058_, _27057_, _27054_);
  or _72678_ (_27059_, _27058_, _27051_);
  or _72679_ (_27060_, _27059_, _27044_);
  or _72680_ (_27061_, _27060_, _27031_);
  or _72681_ (_27062_, _27061_, _27000_);
  or _72682_ (_27063_, _27062_, _26937_);
  or _72683_ (_27064_, _27063_, _26810_);
  and _72684_ (_27065_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or _72685_ (_27066_, _27065_, _27064_);
  and _72686_ (_27067_, _27066_, _00006_);
  or _72687_ (_27068_, _27067_, _26555_);
  and _72688_ (_00003_[7], _27068_, _38997_);
  and _72689_ (_27069_, _26196_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _72690_ (_27070_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _72691_ (_27071_, _27070_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _72692_ (_27072_, _27071_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _72693_ (_27073_, _27072_, _27069_);
  and _72694_ (_27074_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _72695_ (_27075_, _27074_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _72696_ (_27076_, _27075_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _72697_ (_27077_, _27076_, _27073_);
  and _72698_ (_27078_, _27077_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _72699_ (_27079_, _27078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _72700_ (_27080_, _27079_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _72701_ (_27081_, _27079_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _72702_ (_27082_, _27081_, _27080_);
  and _72703_ (_27083_, _27082_, _21983_);
  nor _72704_ (_27084_, _27078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _72705_ (_27085_, _27084_, _27079_);
  and _72706_ (_27086_, _27085_, _21983_);
  nor _72707_ (_27087_, _27077_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor _72708_ (_27088_, _27087_, _27078_);
  and _72709_ (_27089_, _27088_, _21983_);
  nor _72710_ (_27090_, _27085_, _21983_);
  nor _72711_ (_27091_, _27090_, _27086_);
  and _72712_ (_27092_, _27075_, _27073_);
  nor _72713_ (_27093_, _27092_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _72714_ (_27094_, _27092_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _72715_ (_27095_, _27094_, _27093_);
  and _72716_ (_27096_, _27095_, _21983_);
  nor _72717_ (_27097_, _27095_, _21983_);
  and _72718_ (_27098_, _27073_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _72719_ (_27099_, _27098_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _72720_ (_27100_, _27099_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _72721_ (_27101_, _27100_, _27092_);
  and _72722_ (_27102_, _27101_, _21983_);
  nor _72723_ (_27103_, _27101_, _21983_);
  nor _72724_ (_27104_, _27103_, _27102_);
  not _72725_ (_27105_, _27104_);
  nor _72726_ (_27106_, _27098_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor _72727_ (_27107_, _27106_, _27099_);
  and _72728_ (_27108_, _27107_, _21983_);
  nor _72729_ (_27109_, _27073_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _72730_ (_27110_, _27109_, _27098_);
  and _72731_ (_27111_, _27110_, _21983_);
  nor _72732_ (_27112_, _27107_, _21983_);
  nor _72733_ (_27113_, _27112_, _27108_);
  and _72734_ (_27114_, _27071_, _27069_);
  nor _72735_ (_27115_, _27114_, _16218_);
  and _72736_ (_27116_, _27114_, _16218_);
  nor _72737_ (_27117_, _27116_, _27115_);
  not _72738_ (_27118_, _27117_);
  and _72739_ (_27119_, _27118_, _21983_);
  nor _72740_ (_27120_, _27118_, _21983_);
  and _72741_ (_27121_, _27070_, _27069_);
  nor _72742_ (_27122_, _27121_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _72743_ (_27123_, _27122_, _27114_);
  and _72744_ (_27124_, _27123_, _21690_);
  nor _72745_ (_27125_, _27123_, _21690_);
  nor _72746_ (_27126_, _27125_, _27124_);
  not _72747_ (_27127_, _27126_);
  and _72748_ (_27128_, _27069_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _72749_ (_27129_, _27128_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _72750_ (_27130_, _27129_, _27121_);
  and _72751_ (_27131_, _27130_, _21732_);
  nor _72752_ (_27132_, _27130_, _21732_);
  nor _72753_ (_27133_, _27132_, _27131_);
  not _72754_ (_27134_, _27133_);
  nor _72755_ (_27135_, _27069_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _72756_ (_27136_, _27135_, _27128_);
  and _72757_ (_27137_, _27136_, _21774_);
  nor _72758_ (_27138_, _26196_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _72759_ (_27139_, _27138_, _27069_);
  not _72760_ (_27140_, _27139_);
  and _72761_ (_27141_, _21816_, _27140_);
  nor _72762_ (_27142_, _21816_, _27140_);
  nor _72763_ (_27143_, _27142_, _27141_);
  not _72764_ (_27144_, _27143_);
  nor _72765_ (_27145_, _26210_, _26165_);
  not _72766_ (_27146_, _27145_);
  and _72767_ (_27147_, _27146_, _21857_);
  and _72768_ (_27148_, _21898_, _16194_);
  and _72769_ (_27149_, _21940_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _72770_ (_27150_, _21898_, _16194_);
  nor _72771_ (_27151_, _27150_, _27148_);
  and _72772_ (_27152_, _27151_, _27149_);
  nor _72773_ (_27153_, _27152_, _27148_);
  nor _72774_ (_27154_, _27146_, _21857_);
  nor _72775_ (_27155_, _27154_, _27147_);
  not _72776_ (_27156_, _27155_);
  nor _72777_ (_27157_, _27156_, _27153_);
  nor _72778_ (_27158_, _27157_, _27147_);
  nor _72779_ (_27159_, _27158_, _27144_);
  nor _72780_ (_27160_, _27159_, _27141_);
  nor _72781_ (_27161_, _27136_, _21774_);
  nor _72782_ (_27162_, _27161_, _27137_);
  not _72783_ (_27163_, _27162_);
  nor _72784_ (_27164_, _27163_, _27160_);
  nor _72785_ (_27165_, _27164_, _27137_);
  nor _72786_ (_27166_, _27165_, _27134_);
  nor _72787_ (_27167_, _27166_, _27131_);
  nor _72788_ (_27168_, _27167_, _27127_);
  nor _72789_ (_27169_, _27168_, _27124_);
  nor _72790_ (_27170_, _27169_, _27120_);
  or _72791_ (_27171_, _27170_, _27119_);
  nor _72792_ (_27172_, _27110_, _21983_);
  nor _72793_ (_27173_, _27172_, _27111_);
  and _72794_ (_27174_, _27173_, _27171_);
  and _72795_ (_27175_, _27174_, _27113_);
  or _72796_ (_27176_, _27175_, _27111_);
  nor _72797_ (_27177_, _27176_, _27108_);
  nor _72798_ (_27178_, _27177_, _27105_);
  nor _72799_ (_27179_, _27178_, _27102_);
  nor _72800_ (_27180_, _27179_, _27097_);
  nor _72801_ (_27181_, _27180_, _27096_);
  nor _72802_ (_27182_, _27088_, _21983_);
  nor _72803_ (_27183_, _27182_, _27089_);
  not _72804_ (_27184_, _27183_);
  nor _72805_ (_27185_, _27184_, _27181_);
  and _72806_ (_27186_, _27185_, _27091_);
  or _72807_ (_27187_, _27186_, _27089_);
  nor _72808_ (_27188_, _27187_, _27086_);
  nor _72809_ (_27189_, _27082_, _21983_);
  nor _72810_ (_27190_, _27189_, _27083_);
  not _72811_ (_27191_, _27190_);
  nor _72812_ (_27192_, _27191_, _27188_);
  nor _72813_ (_27193_, _27192_, _27083_);
  nor _72814_ (_27194_, _27080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _72815_ (_27195_, _27080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _72816_ (_27196_, _27195_, _27194_);
  not _72817_ (_27197_, _27196_);
  and _72818_ (_27198_, _27197_, _21983_);
  nor _72819_ (_27199_, _27197_, _21983_);
  nor _72820_ (_27200_, _27199_, _27198_);
  and _72821_ (_27201_, _27200_, _27193_);
  nor _72822_ (_27202_, _27200_, _27193_);
  or _72823_ (_27203_, _27202_, _27201_);
  nor _72824_ (_27204_, _27203_, cy_reg);
  and _72825_ (_27205_, _27196_, cy_reg);
  nor _72826_ (_27206_, _27205_, _27204_);
  nand _72827_ (_27207_, _27206_, _14142_);
  or _72828_ (_27208_, _27206_, _14142_);
  and _72829_ (_27209_, _27208_, _27207_);
  not _72830_ (_27210_, cy_reg);
  nor _72831_ (_27211_, _27185_, _27089_);
  and _72832_ (_27212_, _27211_, _27091_);
  nor _72833_ (_27213_, _27211_, _27091_);
  nor _72834_ (_27214_, _27213_, _27212_);
  and _72835_ (_27215_, _27214_, _27210_);
  nor _72836_ (_27216_, _27085_, _27210_);
  nor _72837_ (_27217_, _27216_, _27215_);
  nand _72838_ (_27218_, _27217_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _72839_ (_27219_, _27217_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _72840_ (_27220_, _27219_, _27218_);
  and _72841_ (_27221_, _27184_, _27181_);
  nor _72842_ (_27222_, _27221_, _27185_);
  nor _72843_ (_27223_, _27222_, cy_reg);
  nor _72844_ (_27224_, _27088_, _27210_);
  nor _72845_ (_27225_, _27224_, _27223_);
  nand _72846_ (_27226_, _27225_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _72847_ (_27227_, _27225_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _72848_ (_27228_, _27227_, _27226_);
  and _72849_ (_27229_, _27177_, _27105_);
  nor _72850_ (_27230_, _27229_, _27178_);
  or _72851_ (_27231_, _27230_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nand _72852_ (_27232_, _27230_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _72853_ (_27233_, _27232_, _27231_);
  nor _72854_ (_27234_, _27097_, _27096_);
  nor _72855_ (_27235_, _27234_, _27179_);
  and _72856_ (_27236_, _27234_, _27179_);
  nor _72857_ (_27237_, _27236_, _27235_);
  or _72858_ (_27238_, _27237_, _14106_);
  nand _72859_ (_27239_, _27237_, _14106_);
  and _72860_ (_27240_, _27239_, _27238_);
  or _72861_ (_27241_, _27240_, _27233_);
  or _72862_ (_27242_, _27241_, cy_reg);
  nor _72863_ (_27243_, _27101_, _14121_);
  and _72864_ (_27244_, _27101_, _14121_);
  or _72865_ (_27245_, _27244_, _27243_);
  nor _72866_ (_27246_, _27095_, _14106_);
  and _72867_ (_27247_, _27095_, _14106_);
  or _72868_ (_27248_, _27247_, _27246_);
  or _72869_ (_27249_, _27248_, _27210_);
  or _72870_ (_27250_, _27249_, _27245_);
  and _72871_ (_27251_, _27250_, _27242_);
  nor _72872_ (_27252_, _27174_, _27111_);
  and _72873_ (_27253_, _27252_, _27113_);
  nor _72874_ (_27254_, _27252_, _27113_);
  nor _72875_ (_27255_, _27254_, _27253_);
  nor _72876_ (_27256_, _27255_, cy_reg);
  and _72877_ (_27257_, _27107_, cy_reg);
  nor _72878_ (_27258_, _27257_, _27256_);
  nor _72879_ (_27259_, _27258_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _72880_ (_27260_, _27258_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _72881_ (_27261_, _27110_, cy_reg);
  nor _72882_ (_27262_, _27173_, _27171_);
  nor _72883_ (_27263_, _27262_, _27174_);
  and _72884_ (_27264_, _27263_, _27210_);
  nor _72885_ (_27265_, _27264_, _27261_);
  and _72886_ (_27266_, _27265_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _72887_ (_27267_, _27265_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _72888_ (_27268_, _27117_, _27210_);
  nor _72889_ (_27269_, _27119_, _27120_);
  nor _72890_ (_27270_, _27269_, _27169_);
  and _72891_ (_27271_, _27269_, _27169_);
  or _72892_ (_27272_, _27271_, _27270_);
  and _72893_ (_27273_, _27272_, _27210_);
  nor _72894_ (_27274_, _27273_, _27268_);
  and _72895_ (_27275_, _27274_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _72896_ (_27276_, _27274_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _72897_ (_27277_, _27123_, cy_reg);
  and _72898_ (_27278_, _27167_, _27127_);
  nor _72899_ (_27279_, _27278_, _27168_);
  and _72900_ (_27280_, _27279_, _27210_);
  nor _72901_ (_27281_, _27280_, _27277_);
  and _72902_ (_27282_, _27281_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _72903_ (_27283_, _27281_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _72904_ (_27284_, _27165_, _27134_);
  nor _72905_ (_27285_, _27284_, _27166_);
  and _72906_ (_27286_, _27285_, _27210_);
  and _72907_ (_27287_, _27130_, cy_reg);
  nor _72908_ (_27288_, _27287_, _27286_);
  and _72909_ (_27289_, _27288_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _72910_ (_27290_, _27288_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _72911_ (_27291_, _27136_, cy_reg);
  and _72912_ (_27292_, _27163_, _27160_);
  nor _72913_ (_27293_, _27292_, _27164_);
  and _72914_ (_27294_, _27293_, _27210_);
  nor _72915_ (_27295_, _27294_, _27291_);
  and _72916_ (_27296_, _27295_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _72917_ (_27297_, _27158_, _27144_);
  nor _72918_ (_27298_, _27297_, _27159_);
  and _72919_ (_27299_, _27298_, _27210_);
  nor _72920_ (_27300_, _27139_, _27210_);
  nor _72921_ (_27301_, _27300_, _27299_);
  and _72922_ (_27302_, _27301_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _72923_ (_27303_, _27301_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _72924_ (_27304_, _27156_, _27153_);
  nor _72925_ (_27305_, _27304_, _27157_);
  and _72926_ (_27306_, _27305_, _27210_);
  nor _72927_ (_27307_, _27145_, _27210_);
  nor _72928_ (_27308_, _27307_, _27306_);
  and _72929_ (_27309_, _27308_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _72930_ (_27310_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _72931_ (_27311_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _72932_ (_27312_, _27311_, _27310_);
  not _72933_ (_27313_, _27312_);
  and _72934_ (_27314_, _21940_, _27210_);
  nand _72935_ (_27315_, _27314_, _27313_);
  or _72936_ (_27316_, _27314_, _27313_);
  and _72937_ (_27317_, _27316_, _27315_);
  and _72938_ (_27318_, cy_reg, _16194_);
  nor _72939_ (_27319_, _27151_, _27149_);
  nor _72940_ (_27320_, _27319_, _27152_);
  and _72941_ (_27321_, _27320_, _27210_);
  nor _72942_ (_27322_, _27321_, _27318_);
  nor _72943_ (_27323_, _27322_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _72944_ (_27324_, _27322_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _72945_ (_27325_, _27324_, _27323_);
  or _72946_ (_27326_, _27325_, _27317_);
  nor _72947_ (_27327_, _27308_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _72948_ (_27328_, _27327_, _27326_);
  or _72949_ (_27329_, _27328_, _27309_);
  or _72950_ (_27330_, _27329_, _27303_);
  or _72951_ (_27331_, _27330_, _27302_);
  nor _72952_ (_27332_, _27295_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or _72953_ (_27333_, _27332_, _27331_);
  or _72954_ (_27334_, _27333_, _27296_);
  or _72955_ (_27335_, _27334_, _27290_);
  or _72956_ (_27336_, _27335_, _27289_);
  or _72957_ (_27337_, _27336_, _27283_);
  or _72958_ (_27338_, _27337_, _27282_);
  or _72959_ (_27339_, _27338_, _27276_);
  or _72960_ (_27340_, _27339_, _27275_);
  or _72961_ (_27341_, _27340_, _27267_);
  or _72962_ (_27342_, _27341_, _27266_);
  or _72963_ (_27343_, _27342_, _27260_);
  or _72964_ (_27344_, _27343_, _27259_);
  or _72965_ (_27345_, _27344_, _27251_);
  or _72966_ (_27346_, _27345_, _27228_);
  or _72967_ (_27347_, _27346_, _27220_);
  and _72968_ (_27348_, _27191_, _27188_);
  nor _72969_ (_27349_, _27348_, _27192_);
  nor _72970_ (_27350_, _27349_, cy_reg);
  nor _72971_ (_27351_, _27082_, _27210_);
  nor _72972_ (_27352_, _27351_, _27350_);
  and _72973_ (_27353_, _27352_, _14137_);
  nor _72974_ (_27354_, _27352_, _14137_);
  or _72975_ (_27355_, _27354_, _27353_);
  or _72976_ (_27356_, _27355_, _27347_);
  or _72977_ (_27357_, _27356_, _27209_);
  and _72978_ (_27358_, _26323_, _26190_);
  nor _72979_ (_27359_, _27358_, _26236_);
  and _72980_ (_27360_, _26366_, _26190_);
  nor _72981_ (_27361_, _27360_, _26280_);
  and _72982_ (_27362_, _27361_, _27359_);
  not _72983_ (_27363_, _26545_);
  and _72984_ (_27364_, _27363_, _26502_);
  and _72985_ (_27365_, _27364_, _27362_);
  not _72986_ (_27366_, _26457_);
  and _72987_ (_27367_, _27366_, _26413_);
  or _72988_ (_27368_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _72989_ (_27369_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _72990_ (_27370_, \oc8051_symbolic_cxrom1.regvalid [1], _27369_);
  and _72991_ (_27371_, _27370_, _15852_);
  and _72992_ (_27372_, _27371_, _27368_);
  or _72993_ (_27373_, \oc8051_symbolic_cxrom1.regvalid [13], _27369_);
  or _72994_ (_27374_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _72995_ (_27375_, _27374_, _27373_);
  not _72996_ (_27376_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _72997_ (_27377_, _27376_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _72998_ (_27378_, _27377_, _27375_);
  or _72999_ (_27379_, _27378_, _27372_);
  not _73000_ (_27380_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _73001_ (_27381_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _73002_ (_27382_, _27381_, _27376_);
  nor _73003_ (_27383_, _27382_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _73004_ (_27384_, _27382_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _73005_ (_27385_, _27384_, _27383_);
  and _73006_ (_27386_, _27385_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _73007_ (_27387_, _27381_, _27376_);
  nor _73008_ (_27388_, _27387_, _27382_);
  nand _73009_ (_27389_, \oc8051_symbolic_cxrom1.regvalid [7], _27369_);
  nand _73010_ (_27390_, _27389_, _27388_);
  or _73011_ (_27391_, _27390_, _27386_);
  and _73012_ (_27392_, _27391_, _27380_);
  nor _73013_ (_27393_, _27385_, _18609_);
  and _73014_ (_27394_, _27385_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _73015_ (_27395_, _27394_, _27393_);
  or _73016_ (_27396_, _27388_, _27395_);
  and _73017_ (_27397_, _27396_, _27392_);
  or _73018_ (_27398_, _27397_, _27379_);
  and _73019_ (_27399_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _73020_ (_27400_, \oc8051_symbolic_cxrom1.regvalid [0], _27369_);
  or _73021_ (_27401_, _27400_, _27399_);
  and _73022_ (_27402_, _27401_, _27376_);
  and _73023_ (_27403_, \oc8051_symbolic_cxrom1.regvalid [4], _27369_);
  and _73024_ (_27404_, \oc8051_symbolic_cxrom1.regvalid [12], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _73025_ (_27405_, _27404_, _27403_);
  and _73026_ (_27406_, _27405_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _73027_ (_27407_, _27406_, _27402_);
  and _73028_ (_27408_, _27407_, _27380_);
  and _73029_ (_27409_, _15852_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _73030_ (_27410_, _27409_, _27369_);
  and _73031_ (_27411_, _27409_, _27369_);
  nor _73032_ (_27412_, _27411_, _27410_);
  nand _73033_ (_27413_, _27412_, _18508_);
  and _73034_ (_27414_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _73035_ (_27415_, _27414_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _73036_ (_27416_, _27415_, _27409_);
  and _73037_ (_27417_, _27416_, _27373_);
  and _73038_ (_27418_, _27417_, _27413_);
  or _73039_ (_27419_, _27412_, \oc8051_symbolic_cxrom1.regvalid [9]);
  not _73040_ (_27420_, _27416_);
  nand _73041_ (_27421_, _27412_, _18635_);
  and _73042_ (_27422_, _27421_, _27420_);
  and _73043_ (_27423_, _27422_, _27419_);
  or _73044_ (_27424_, _27423_, _27418_);
  and _73045_ (_27425_, _27424_, _27408_);
  not _73046_ (_27426_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand _73047_ (_27427_, _27412_, _27426_);
  or _73048_ (_27428_, \oc8051_symbolic_cxrom1.regvalid [15], _27369_);
  and _73049_ (_27429_, _27428_, _27416_);
  and _73050_ (_27430_, _27429_, _27427_);
  or _73051_ (_27431_, _27412_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nand _73052_ (_27432_, _27412_, _18609_);
  and _73053_ (_27433_, _27432_, _27420_);
  and _73054_ (_27434_, _27433_, _27431_);
  or _73055_ (_27435_, _27434_, _27430_);
  and _73056_ (_27436_, \oc8051_symbolic_cxrom1.regvalid [14], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _73057_ (_27437_, \oc8051_symbolic_cxrom1.regvalid [6], _27369_);
  or _73058_ (_27438_, _27437_, _27376_);
  or _73059_ (_27439_, _27438_, _27436_);
  or _73060_ (_27440_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _73061_ (_27441_, \oc8051_symbolic_cxrom1.regvalid [10], _27369_);
  and _73062_ (_27442_, _27441_, _27440_);
  or _73063_ (_27443_, _27442_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _73064_ (_27444_, _27443_, _27439_);
  and _73065_ (_27445_, _27444_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _73066_ (_27446_, _27405_, _27377_);
  or _73067_ (_27447_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _73068_ (_27448_, \oc8051_symbolic_cxrom1.regvalid [0], _27369_);
  and _73069_ (_27449_, _27448_, _15852_);
  and _73070_ (_27450_, _27449_, _27447_);
  or _73071_ (_27451_, _27450_, _27446_);
  and _73072_ (_27452_, _27451_, _27445_);
  and _73073_ (_27453_, _27452_, _27435_);
  or _73074_ (_27454_, _27453_, _27425_);
  not _73075_ (_27455_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _73076_ (_27456_, _27451_, _27444_);
  and _73077_ (_27457_, _27456_, _27455_);
  and _73078_ (_27458_, _27457_, _27454_);
  and _73079_ (_27459_, _27458_, _27398_);
  or _73080_ (_27460_, \oc8051_symbolic_cxrom1.regvalid [2], _27380_);
  or _73081_ (_27461_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _73082_ (_27462_, _27461_, _27460_);
  or _73083_ (_27463_, _27462_, _27385_);
  or _73084_ (_27464_, \oc8051_symbolic_cxrom1.regvalid [10], _27380_);
  or _73085_ (_27465_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand _73086_ (_27466_, _27465_, _27464_);
  and _73087_ (_27467_, _27466_, _27385_);
  nor _73088_ (_27468_, _27467_, _27388_);
  and _73089_ (_27469_, _27468_, _27463_);
  and _73090_ (_27470_, _27385_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _73091_ (_27471_, _27403_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _73092_ (_27472_, _27471_, _27470_);
  and _73093_ (_27473_, _27385_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or _73094_ (_27474_, _27437_, _27380_);
  or _73095_ (_27475_, _27474_, _27473_);
  and _73096_ (_27476_, _27475_, _27388_);
  and _73097_ (_27477_, _27476_, _27472_);
  or _73098_ (_27478_, _27477_, _27469_);
  nand _73099_ (_27479_, _27412_, _18543_);
  or _73100_ (_27480_, \oc8051_symbolic_cxrom1.regvalid [14], _27369_);
  and _73101_ (_27481_, _27480_, _27479_);
  or _73102_ (_27482_, _27481_, _27420_);
  or _73103_ (_27483_, _27412_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand _73104_ (_27484_, _27412_, _18644_);
  and _73105_ (_27485_, _27484_, _27483_);
  or _73106_ (_27486_, _27485_, _27416_);
  and _73107_ (_27487_, _27486_, _27482_);
  or _73108_ (_27488_, _27487_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _73109_ (_27489_, _27412_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nand _73110_ (_27490_, _27412_, _18657_);
  and _73111_ (_27491_, _27490_, _27420_);
  and _73112_ (_27492_, _27491_, _27489_);
  nand _73113_ (_27493_, _27412_, _18532_);
  or _73114_ (_27494_, \oc8051_symbolic_cxrom1.regvalid [12], _27369_);
  and _73115_ (_27495_, _27494_, _27416_);
  and _73116_ (_27496_, _27495_, _27493_);
  or _73117_ (_27497_, _27496_, _27380_);
  or _73118_ (_27498_, _27497_, _27492_);
  or _73119_ (_27499_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _73120_ (_27500_, _27499_, _27428_);
  or _73121_ (_27501_, _27500_, _27376_);
  or _73122_ (_27502_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _73123_ (_27503_, \oc8051_symbolic_cxrom1.regvalid [11], _27369_);
  and _73124_ (_27504_, _27503_, _27502_);
  or _73125_ (_27505_, _27504_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _73126_ (_27506_, _27505_, _27501_);
  and _73127_ (_27507_, _27506_, _27414_);
  and _73128_ (_27508_, _27380_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _73129_ (_27509_, _27375_, _27376_);
  or _73130_ (_27510_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _73131_ (_27511_, \oc8051_symbolic_cxrom1.regvalid [9], _27369_);
  and _73132_ (_27512_, _27511_, _27510_);
  or _73133_ (_27513_, _27512_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _73134_ (_27514_, _27513_, _27509_);
  and _73135_ (_27515_, _27514_, _27508_);
  or _73136_ (_27516_, _27515_, _27507_);
  and _73137_ (_27517_, _27506_, _27380_);
  or _73138_ (_27518_, _27517_, _27379_);
  and _73139_ (_27519_, _27518_, _27516_);
  and _73140_ (_27520_, _27519_, _27498_);
  and _73141_ (_27521_, _27520_, _27488_);
  and _73142_ (_27522_, _27521_, _27478_);
  or _73143_ (_27523_, _27522_, _27459_);
  nor _73144_ (_27524_, _26178_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _73145_ (_27525_, _26210_, _26185_);
  nor _73146_ (_27526_, _27525_, _27524_);
  nor _73147_ (_27527_, _27526_, _16190_);
  not _73148_ (_27528_, _27527_);
  and _73149_ (_27529_, _26156_, _16194_);
  and _73150_ (_27530_, _26210_, _26164_);
  nor _73151_ (_27531_, _27530_, _27529_);
  nor _73152_ (_27532_, _27531_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _73153_ (_27533_, _21603_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _73154_ (_27534_, _18657_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _73155_ (_27535_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _73156_ (_27536_, _27535_, _27534_);
  and _73157_ (_27537_, _27536_, _27533_);
  and _73158_ (_27538_, _18635_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _73159_ (_27539_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _73160_ (_27540_, _27539_, _27538_);
  and _73161_ (_27541_, _27540_, _21596_);
  nor _73162_ (_27542_, _27541_, _27537_);
  not _73163_ (_27543_, _27542_);
  nor _73164_ (_27544_, _27543_, _27532_);
  and _73165_ (_27545_, _27544_, _27528_);
  not _73166_ (_27546_, _27545_);
  and _73167_ (_27547_, _27546_, _26190_);
  nor _73168_ (_27548_, _21608_, _16198_);
  and _73169_ (_27549_, _27548_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _73170_ (_27550_, _27548_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _73171_ (_27551_, _27550_, _27549_);
  nand _73172_ (_27552_, _27551_, _18622_);
  and _73173_ (_27553_, _21608_, _16198_);
  nor _73174_ (_27554_, _27553_, _27548_);
  not _73175_ (_27555_, _27554_);
  nor _73176_ (_27556_, _27555_, _21670_);
  and _73177_ (_27557_, _27556_, _27552_);
  and _73178_ (_27558_, _27551_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _73179_ (_27559_, _27551_, _18609_);
  or _73180_ (_27560_, _27559_, _27558_);
  and _73181_ (_27561_, _27560_, _27555_);
  or _73182_ (_27562_, _27561_, _27557_);
  and _73183_ (_27563_, _27562_, _21608_);
  nand _73184_ (_27564_, _27551_, _18630_);
  nor _73185_ (_27565_, _27555_, _21679_);
  and _73186_ (_27566_, _27565_, _27564_);
  and _73187_ (_27567_, _27551_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _73188_ (_27568_, _27551_, _18635_);
  or _73189_ (_27569_, _27568_, _27567_);
  and _73190_ (_27570_, _27569_, _27555_);
  or _73191_ (_27571_, _27570_, _27566_);
  and _73192_ (_27572_, _27571_, _21603_);
  or _73193_ (_27573_, _27572_, _27563_);
  nand _73194_ (_27574_, _27551_, _18646_);
  or _73195_ (_27575_, _27551_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _73196_ (_27576_, _27575_, _27555_);
  and _73197_ (_27577_, _27576_, _27574_);
  or _73198_ (_27578_, _27551_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _73199_ (_27579_, _27555_, _26149_);
  and _73200_ (_27580_, _27579_, _27578_);
  or _73201_ (_27581_, _27580_, _27577_);
  and _73202_ (_27582_, _27581_, _21595_);
  nand _73203_ (_27583_, _27551_, _18663_);
  nor _73204_ (_27584_, _27555_, _21675_);
  and _73205_ (_27585_, _27584_, _27583_);
  and _73206_ (_27586_, _27551_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _73207_ (_27587_, _27551_, _18657_);
  or _73208_ (_27588_, _27587_, _27586_);
  and _73209_ (_27589_, _27588_, _27555_);
  or _73210_ (_27590_, _27589_, _27585_);
  and _73211_ (_27591_, _27590_, _21605_);
  or _73212_ (_27592_, _27591_, _27582_);
  or _73213_ (_27593_, _27592_, _27573_);
  and _73214_ (_27594_, _27593_, _21689_);
  and _73215_ (_27595_, _27594_, _27547_);
  and _73216_ (_27596_, _27595_, _27523_);
  and _73217_ (_27597_, _15585_, _26138_);
  and _73218_ (_27598_, _27597_, _27596_);
  and _73219_ (_27599_, _27598_, _27367_);
  and _73220_ (_27600_, _27599_, _27365_);
  and _73221_ (property_invalid_jnc, _27600_, _27357_);
  and _73222_ (_27601_, _27196_, _27210_);
  nor _73223_ (_27602_, _27203_, _27210_);
  nor _73224_ (_27603_, _27602_, _27601_);
  and _73225_ (_27604_, _27603_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _73226_ (_27605_, _27603_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or _73227_ (_27606_, _27088_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand _73228_ (_27607_, _27088_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _73229_ (_27608_, _27607_, _27606_);
  and _73230_ (_27609_, _27085_, _14132_);
  nor _73231_ (_27610_, _27085_, _14132_);
  or _73232_ (_27611_, _27610_, _27609_);
  or _73233_ (_27612_, _27611_, _27608_);
  or _73234_ (_27613_, _27612_, cy_reg);
  or _73235_ (_27614_, _27214_, _14132_);
  nand _73236_ (_27615_, _27214_, _14132_);
  and _73237_ (_27616_, _27615_, _27614_);
  or _73238_ (_27617_, _27222_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand _73239_ (_27618_, _27222_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _73240_ (_27619_, _27618_, _27617_);
  or _73241_ (_27620_, _27619_, _27210_);
  or _73242_ (_27621_, _27620_, _27616_);
  and _73243_ (_27622_, _27621_, _27613_);
  and _73244_ (_27623_, _27095_, _27210_);
  nor _73245_ (_27624_, _27237_, _27210_);
  nor _73246_ (_27625_, _27624_, _27623_);
  and _73247_ (_27626_, _27625_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _73248_ (_27627_, _27625_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _73249_ (_27628_, _27107_, _27210_);
  nor _73250_ (_27629_, _27255_, _27210_);
  nor _73251_ (_27630_, _27629_, _27628_);
  and _73252_ (_27631_, _27630_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _73253_ (_27632_, _27630_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _73254_ (_27633_, _27117_, cy_reg);
  and _73255_ (_27634_, _27272_, cy_reg);
  nor _73256_ (_27635_, _27634_, _27633_);
  and _73257_ (_27636_, _27635_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _73258_ (_27637_, _27635_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _73259_ (_27638_, _27123_, _27210_);
  and _73260_ (_27639_, _27279_, cy_reg);
  nor _73261_ (_27640_, _27639_, _27638_);
  and _73262_ (_27641_, _27640_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _73263_ (_27642_, _27640_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _73264_ (_27643_, _27285_, cy_reg);
  and _73265_ (_27644_, _27130_, _27210_);
  nor _73266_ (_27645_, _27644_, _27643_);
  and _73267_ (_27646_, _27645_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _73268_ (_27647_, _27645_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _73269_ (_27648_, _27136_, _27210_);
  and _73270_ (_27649_, _27293_, cy_reg);
  nor _73271_ (_27650_, _27649_, _27648_);
  and _73272_ (_27651_, _27650_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _73273_ (_27652_, _27139_, cy_reg);
  and _73274_ (_27653_, _27298_, cy_reg);
  nor _73275_ (_27654_, _27653_, _27652_);
  and _73276_ (_27655_, _27654_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _73277_ (_27656_, _27654_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _73278_ (_27657_, _27305_, cy_reg);
  nor _73279_ (_27658_, _27145_, cy_reg);
  nor _73280_ (_27659_, _27658_, _27657_);
  and _73281_ (_27660_, _27659_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _73282_ (_27661_, cy_reg, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _73283_ (_27662_, _27320_, cy_reg);
  nor _73284_ (_27663_, _27662_, _27661_);
  and _73285_ (_27664_, _27663_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _73286_ (_27665_, _27312_, _21940_);
  nor _73287_ (_27666_, _27312_, _21940_);
  or _73288_ (_27667_, _27666_, _27665_);
  or _73289_ (_27668_, _27667_, _27210_);
  nand _73290_ (_27669_, _27312_, _27210_);
  and _73291_ (_27670_, _27669_, _27668_);
  nor _73292_ (_27671_, _27663_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _73293_ (_27672_, _27671_, _27670_);
  or _73294_ (_27673_, _27672_, _27664_);
  nor _73295_ (_27674_, _27659_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _73296_ (_27675_, _27674_, _27673_);
  or _73297_ (_27676_, _27675_, _27660_);
  or _73298_ (_27677_, _27676_, _27656_);
  or _73299_ (_27678_, _27677_, _27655_);
  nor _73300_ (_27679_, _27650_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or _73301_ (_27680_, _27679_, _27678_);
  or _73302_ (_27681_, _27680_, _27651_);
  or _73303_ (_27682_, _27681_, _27647_);
  or _73304_ (_27683_, _27682_, _27646_);
  or _73305_ (_27684_, _27683_, _27642_);
  or _73306_ (_27685_, _27684_, _27641_);
  or _73307_ (_27686_, _27685_, _27637_);
  or _73308_ (_27687_, _27686_, _27636_);
  and _73309_ (_27688_, _27110_, _27210_);
  and _73310_ (_27689_, _27263_, cy_reg);
  nor _73311_ (_27690_, _27689_, _27688_);
  nor _73312_ (_27691_, _27690_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _73313_ (_27692_, _27690_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _73314_ (_27693_, _27692_, _27691_);
  or _73315_ (_27694_, _27693_, _27687_);
  or _73316_ (_27695_, _27694_, _27632_);
  or _73317_ (_27696_, _27695_, _27631_);
  and _73318_ (_27697_, _27101_, _27210_);
  and _73319_ (_27698_, _27230_, cy_reg);
  nor _73320_ (_27699_, _27698_, _27697_);
  and _73321_ (_27700_, _27699_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _73322_ (_27701_, _27699_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _73323_ (_27702_, _27701_, _27700_);
  or _73324_ (_27703_, _27702_, _27696_);
  or _73325_ (_27704_, _27703_, _27627_);
  or _73326_ (_27705_, _27704_, _27626_);
  or _73327_ (_27706_, _27705_, _27622_);
  nor _73328_ (_27707_, _27082_, cy_reg);
  nor _73329_ (_27708_, _27349_, _27210_);
  nor _73330_ (_27709_, _27708_, _27707_);
  and _73331_ (_27710_, _27709_, _14137_);
  nor _73332_ (_27711_, _27709_, _14137_);
  or _73333_ (_27712_, _27711_, _27710_);
  or _73334_ (_27713_, _27712_, _27706_);
  or _73335_ (_27714_, _27713_, _27605_);
  or _73336_ (_27715_, _27714_, _27604_);
  and _73337_ (_27716_, _27362_, _26547_);
  and _73338_ (_27717_, _27716_, _27599_);
  and _73339_ (property_invalid_jc, _27717_, _27715_);
  or _73340_ (_27718_, _21898_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand _73341_ (_27719_, _21898_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _73342_ (_27720_, _27719_, _27718_);
  and _73343_ (_27721_, _21940_, _27455_);
  nor _73344_ (_27722_, _21940_, _27455_);
  or _73345_ (_27723_, _27722_, _27721_);
  or _73346_ (_27724_, _27723_, _27720_);
  or _73347_ (_27725_, _21816_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand _73348_ (_27726_, _21816_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _73349_ (_27727_, _27726_, _27725_);
  and _73350_ (_27728_, _21857_, _27376_);
  nor _73351_ (_27729_, _21857_, _27376_);
  or _73352_ (_27730_, _27729_, _27728_);
  or _73353_ (_27731_, _27730_, _27727_);
  or _73354_ (_27732_, _27731_, _27724_);
  or _73355_ (_27733_, _21732_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand _73356_ (_27734_, _21732_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _73357_ (_27735_, _27734_, _27733_);
  not _73358_ (_27736_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _73359_ (_27737_, _21774_, _27736_);
  and _73360_ (_27738_, _21774_, _27736_);
  or _73361_ (_27739_, _27738_, _27737_);
  or _73362_ (_27740_, _27739_, _27735_);
  not _73363_ (_27741_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _73364_ (_27742_, _21983_, _27741_);
  nor _73365_ (_27743_, _21983_, _27741_);
  or _73366_ (_27744_, _27743_, _27742_);
  not _73367_ (_27745_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _73368_ (_27746_, _21690_, _27745_);
  nor _73369_ (_27747_, _21690_, _27745_);
  or _73370_ (_27748_, _27747_, _27746_);
  or _73371_ (_27749_, _27748_, _27744_);
  or _73372_ (_27750_, _27749_, _27740_);
  or _73373_ (_27751_, _27750_, _27732_);
  nor _73374_ (_27752_, _27196_, _14142_);
  and _73375_ (_27753_, _27196_, _14142_);
  or _73376_ (_27754_, _27753_, _27752_);
  nor _73377_ (_27755_, _27082_, _14137_);
  and _73378_ (_27756_, _27082_, _14137_);
  or _73379_ (_27757_, _27756_, _27755_);
  or _73380_ (_27758_, _27757_, _27612_);
  or _73381_ (_27759_, _27758_, _27754_);
  nor _73382_ (_27760_, _26546_, _14110_);
  and _73383_ (_27761_, _26546_, _14110_);
  or _73384_ (_27762_, _27761_, _27760_);
  nor _73385_ (_27763_, _26413_, _14116_);
  and _73386_ (_27764_, _26413_, _14116_);
  or _73387_ (_27765_, _27764_, _27763_);
  or _73388_ (_27766_, _27765_, _27762_);
  and _73389_ (_27767_, _26457_, _14121_);
  nor _73390_ (_27768_, _26457_, _14121_);
  or _73391_ (_27769_, _27768_, _27767_);
  or _73392_ (_27770_, _27769_, _27248_);
  or _73393_ (_27771_, _27770_, _27766_);
  or _73394_ (_27772_, _27771_, _27759_);
  or _73395_ (_27773_, _27772_, _27751_);
  nor _73396_ (_27774_, _26323_, _26550_);
  and _73397_ (_27775_, _27361_, _27774_);
  and _73398_ (_27776_, _27775_, _27598_);
  and _73399_ (property_invalid_ajmp, _27776_, _27773_);
  and _73400_ (_27777_, _26210_, _26193_);
  and _73401_ (_27778_, _26199_, _26165_);
  and _73402_ (_27779_, _26203_, _26196_);
  or _73403_ (_27780_, _27779_, _27778_);
  or _73404_ (_27781_, _27780_, _27777_);
  and _73405_ (_27782_, _26209_, _26158_);
  or _73406_ (_27783_, _27782_, _27140_);
  or _73407_ (_27784_, _27783_, _27781_);
  and _73408_ (_27785_, _26216_, _26210_);
  or _73409_ (_27786_, _27785_, _27139_);
  and _73410_ (_27787_, _26225_, _26196_);
  and _73411_ (_27788_, _26231_, _26158_);
  and _73412_ (_27789_, _26221_, _26165_);
  or _73413_ (_27790_, _27789_, _27788_);
  or _73414_ (_27791_, _27790_, _27787_);
  or _73415_ (_27792_, _27791_, _27786_);
  nand _73416_ (_27793_, _27792_, _27784_);
  nor _73417_ (_27794_, _27793_, _27545_);
  nand _73418_ (_27795_, _27794_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _73419_ (_27796_, _27794_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _73420_ (_27797_, _27796_, _27795_);
  and _73421_ (_27798_, _26461_, _26210_);
  and _73422_ (_27799_, _26466_, _26165_);
  and _73423_ (_27800_, _26470_, _26196_);
  or _73424_ (_27801_, _27800_, _27799_);
  or _73425_ (_27802_, _27801_, _27798_);
  and _73426_ (_27803_, _26476_, _26158_);
  or _73427_ (_27804_, _27803_, _27140_);
  or _73428_ (_27805_, _27804_, _27802_);
  and _73429_ (_27806_, _26482_, _26210_);
  or _73430_ (_27807_, _27806_, _27139_);
  and _73431_ (_27808_, _26491_, _26196_);
  and _73432_ (_27809_, _26497_, _26158_);
  and _73433_ (_27810_, _26487_, _26165_);
  or _73434_ (_27811_, _27810_, _27809_);
  or _73435_ (_27812_, _27811_, _27808_);
  or _73436_ (_27813_, _27812_, _27807_);
  nand _73437_ (_27814_, _27813_, _27805_);
  nor _73438_ (_27815_, _27814_, _27545_);
  nand _73439_ (_27816_, _27815_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or _73440_ (_27817_, _27815_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _73441_ (_27818_, _27817_, _27816_);
  or _73442_ (_27819_, _27818_, _27797_);
  and _73443_ (_27820_, _26326_, _26210_);
  and _73444_ (_27821_, _26331_, _26165_);
  and _73445_ (_27822_, _26335_, _26196_);
  or _73446_ (_27823_, _27822_, _27821_);
  or _73447_ (_27824_, _27823_, _27820_);
  and _73448_ (_27825_, _26341_, _26158_);
  or _73449_ (_27826_, _27825_, _27140_);
  or _73450_ (_27827_, _27826_, _27824_);
  and _73451_ (_27828_, _26352_, _26165_);
  or _73452_ (_27829_, _27828_, _27139_);
  and _73453_ (_27830_, _26356_, _26196_);
  and _73454_ (_27831_, _26362_, _26158_);
  and _73455_ (_27832_, _26347_, _26210_);
  or _73456_ (_27833_, _27832_, _27831_);
  or _73457_ (_27834_, _27833_, _27830_);
  or _73458_ (_27835_, _27834_, _27829_);
  nand _73459_ (_27836_, _27835_, _27827_);
  nor _73460_ (_27837_, _27836_, _27545_);
  nand _73461_ (_27838_, _27837_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _73462_ (_27839_, _27837_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _73463_ (_27840_, _27839_, _27838_);
  and _73464_ (_27841_, _26510_, _26165_);
  and _73465_ (_27842_, _26505_, _26210_);
  and _73466_ (_27843_, _26514_, _26196_);
  or _73467_ (_27844_, _27843_, _27842_);
  or _73468_ (_27845_, _27844_, _27841_);
  and _73469_ (_27846_, _26520_, _26158_);
  or _73470_ (_27847_, _27846_, _27140_);
  or _73471_ (_27848_, _27847_, _27845_);
  and _73472_ (_27849_, _26526_, _26210_);
  or _73473_ (_27850_, _27849_, _27139_);
  and _73474_ (_27851_, _26535_, _26196_);
  and _73475_ (_27852_, _26541_, _26158_);
  and _73476_ (_27853_, _26531_, _26165_);
  or _73477_ (_27854_, _27853_, _27852_);
  or _73478_ (_27855_, _27854_, _27851_);
  or _73479_ (_27856_, _27855_, _27850_);
  nand _73480_ (_27857_, _27856_, _27848_);
  nor _73481_ (_27858_, _27857_, _27545_);
  nand _73482_ (_27859_, _27858_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or _73483_ (_27860_, _27858_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _73484_ (_27861_, _27860_, _27859_);
  or _73485_ (_27862_, _27861_, _27840_);
  or _73486_ (_27863_, _27862_, _27819_);
  and _73487_ (_27864_, _26288_, _26165_);
  and _73488_ (_27865_, _26283_, _26210_);
  and _73489_ (_27866_, _26292_, _26196_);
  or _73490_ (_27867_, _27866_, _27865_);
  or _73491_ (_27868_, _27867_, _27864_);
  and _73492_ (_27869_, _26298_, _26158_);
  or _73493_ (_27870_, _27869_, _27140_);
  or _73494_ (_27871_, _27870_, _27868_);
  and _73495_ (_27872_, _26304_, _26210_);
  or _73496_ (_27873_, _27872_, _27139_);
  and _73497_ (_27874_, _26313_, _26196_);
  and _73498_ (_27875_, _26319_, _26158_);
  and _73499_ (_27876_, _26309_, _26165_);
  or _73500_ (_27877_, _27876_, _27875_);
  or _73501_ (_27878_, _27877_, _27874_);
  or _73502_ (_27879_, _27878_, _27873_);
  nand _73503_ (_27880_, _27879_, _27871_);
  nor _73504_ (_27881_, _27880_, _27545_);
  nor _73505_ (_27882_, _27881_, _27380_);
  and _73506_ (_27883_, _27881_, _27380_);
  or _73507_ (_27884_, _27883_, _27882_);
  and _73508_ (_27885_, _26372_, _26210_);
  and _73509_ (_27886_, _26377_, _26165_);
  and _73510_ (_27887_, _26381_, _26196_);
  or _73511_ (_27888_, _27887_, _27886_);
  or _73512_ (_27889_, _27888_, _27885_);
  and _73513_ (_27890_, _26387_, _26158_);
  or _73514_ (_27891_, _27890_, _27140_);
  or _73515_ (_27892_, _27891_, _27889_);
  and _73516_ (_27893_, _26393_, _26210_);
  or _73517_ (_27894_, _27893_, _27139_);
  and _73518_ (_27895_, _26402_, _26196_);
  and _73519_ (_27896_, _26408_, _26158_);
  and _73520_ (_27897_, _26398_, _26165_);
  or _73521_ (_27898_, _27897_, _27896_);
  or _73522_ (_27899_, _27898_, _27895_);
  or _73523_ (_27900_, _27899_, _27894_);
  nand _73524_ (_27901_, _27900_, _27892_);
  nor _73525_ (_27902_, _27901_, _27545_);
  and _73526_ (_27903_, _27902_, _27745_);
  nor _73527_ (_27904_, _27902_, _27745_);
  or _73528_ (_27905_, _27904_, _27903_);
  or _73529_ (_27906_, _27905_, _27884_);
  and _73530_ (_27907_, _26260_, _26210_);
  and _73531_ (_27908_, _26269_, _26196_);
  nor _73532_ (_27909_, _27908_, _27907_);
  and _73533_ (_27910_, _26275_, _26158_);
  and _73534_ (_27911_, _26265_, _26165_);
  nor _73535_ (_27912_, _27911_, _27910_);
  and _73536_ (_27913_, _27912_, _27909_);
  nor _73537_ (_27914_, _27913_, _27139_);
  and _73538_ (_27915_, _26239_, _26210_);
  and _73539_ (_27916_, _26248_, _26196_);
  nor _73540_ (_27917_, _27916_, _27915_);
  and _73541_ (_27918_, _26254_, _26158_);
  and _73542_ (_27919_, _26244_, _26165_);
  nor _73543_ (_27920_, _27919_, _27918_);
  and _73544_ (_27921_, _27920_, _27917_);
  nor _73545_ (_27922_, _27921_, _27140_);
  nor _73546_ (_27923_, _27922_, _27914_);
  nor _73547_ (_27924_, _27923_, _27545_);
  nor _73548_ (_27925_, _27924_, _27376_);
  and _73549_ (_27926_, _27924_, _27376_);
  or _73550_ (_27927_, _27926_, _27925_);
  and _73551_ (_27928_, _26416_, _26210_);
  and _73552_ (_27929_, _26421_, _26165_);
  and _73553_ (_27930_, _26425_, _26196_);
  or _73554_ (_27931_, _27930_, _27929_);
  or _73555_ (_27932_, _27931_, _27928_);
  and _73556_ (_27933_, _26431_, _26158_);
  or _73557_ (_27934_, _27933_, _27140_);
  or _73558_ (_27935_, _27934_, _27932_);
  and _73559_ (_27936_, _26437_, _26210_);
  or _73560_ (_27937_, _27936_, _27139_);
  and _73561_ (_27938_, _26446_, _26196_);
  and _73562_ (_27939_, _26452_, _26158_);
  and _73563_ (_27940_, _26442_, _26165_);
  or _73564_ (_27941_, _27940_, _27939_);
  or _73565_ (_27942_, _27941_, _27938_);
  or _73566_ (_27943_, _27942_, _27937_);
  nand _73567_ (_27944_, _27943_, _27935_);
  nor _73568_ (_27945_, _27944_, _27545_);
  nor _73569_ (_27946_, _27945_, _27741_);
  and _73570_ (_27947_, _27945_, _27741_);
  or _73571_ (_27948_, _27947_, _27946_);
  or _73572_ (_27949_, _27948_, _27927_);
  or _73573_ (_27950_, _27949_, _27906_);
  or _73574_ (_27951_, _27950_, _27863_);
  or _73575_ (_27952_, _21898_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand _73576_ (_27953_, _21898_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _73577_ (_27954_, _27953_, _27952_);
  nor _73578_ (_27955_, _21940_, _14110_);
  and _73579_ (_27956_, _21940_, _14110_);
  or _73580_ (_27957_, _27956_, _27955_);
  or _73581_ (_27958_, _27957_, _27954_);
  or _73582_ (_27959_, _21816_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand _73583_ (_27960_, _21816_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _73584_ (_27961_, _27960_, _27959_);
  and _73585_ (_27962_, _21857_, _14121_);
  nor _73586_ (_27963_, _21857_, _14121_);
  or _73587_ (_27964_, _27963_, _27962_);
  or _73588_ (_27965_, _27964_, _27961_);
  or _73589_ (_27966_, _27965_, _27958_);
  or _73590_ (_27967_, _21732_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _73591_ (_27968_, _21732_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _73592_ (_27969_, _27968_, _27967_);
  and _73593_ (_27970_, _21774_, _14127_);
  nor _73594_ (_27971_, _21774_, _14127_);
  or _73595_ (_27972_, _27971_, _27970_);
  or _73596_ (_27973_, _27972_, _27969_);
  and _73597_ (_27974_, _21983_, _14142_);
  nor _73598_ (_27975_, _21983_, _14142_);
  or _73599_ (_27976_, _27975_, _27974_);
  nor _73600_ (_27977_, _21690_, _14137_);
  and _73601_ (_27978_, _21690_, _14137_);
  or _73602_ (_27979_, _27978_, _27977_);
  or _73603_ (_27980_, _27979_, _27976_);
  or _73604_ (_27981_, _27980_, _27973_);
  or _73605_ (_27982_, _27981_, _27966_);
  or _73606_ (_27983_, _27982_, _27951_);
  not _73607_ (_27984_, _26546_);
  and _73608_ (_27985_, _27984_, _26458_);
  and _73609_ (_27986_, _27361_, _26550_);
  and _73610_ (_27987_, _27986_, _27358_);
  and _73611_ (_27988_, _27987_, _27985_);
  and _73612_ (_27989_, _27988_, _27598_);
  and _73613_ (property_invalid_ljmp, _27989_, _27983_);
  and _73614_ (_27990_, _27203_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _73615_ (_27991_, _27203_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _73616_ (_27992_, _27255_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _73617_ (_27993_, _27255_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _73618_ (_27994_, _27263_, _14110_);
  nor _73619_ (_27995_, _27263_, _14110_);
  and _73620_ (_27996_, _27272_, _27741_);
  nor _73621_ (_27997_, _27272_, _27741_);
  and _73622_ (_27998_, _27279_, _27745_);
  nor _73623_ (_27999_, _27279_, _27745_);
  not _73624_ (_28000_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _73625_ (_28001_, _27285_, _28000_);
  nor _73626_ (_28002_, _27285_, _28000_);
  and _73627_ (_28003_, _27293_, _27736_);
  and _73628_ (_28004_, _27298_, _27369_);
  nor _73629_ (_28005_, _27298_, _27369_);
  and _73630_ (_28006_, _27305_, _27376_);
  or _73631_ (_28007_, _27320_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand _73632_ (_28008_, _27320_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _73633_ (_28009_, _28008_, _28007_);
  or _73634_ (_28010_, _28009_, _27667_);
  nor _73635_ (_28011_, _27305_, _27376_);
  or _73636_ (_28012_, _28011_, _28010_);
  or _73637_ (_28013_, _28012_, _28006_);
  or _73638_ (_28014_, _28013_, _28005_);
  or _73639_ (_28015_, _28014_, _28004_);
  nor _73640_ (_28016_, _27293_, _27736_);
  or _73641_ (_28017_, _28016_, _28015_);
  or _73642_ (_28018_, _28017_, _28003_);
  or _73643_ (_28019_, _28018_, _28002_);
  or _73644_ (_28020_, _28019_, _28001_);
  or _73645_ (_28021_, _28020_, _27999_);
  or _73646_ (_28022_, _28021_, _27998_);
  or _73647_ (_28023_, _28022_, _27997_);
  or _73648_ (_28024_, _28023_, _27996_);
  or _73649_ (_28025_, _28024_, _27995_);
  or _73650_ (_28026_, _28025_, _27994_);
  or _73651_ (_28027_, _28026_, _27993_);
  or _73652_ (_28028_, _28027_, _27992_);
  or _73653_ (_28029_, _28028_, _27241_);
  or _73654_ (_28030_, _28029_, _27619_);
  or _73655_ (_28031_, _28030_, _27616_);
  nor _73656_ (_28032_, _27349_, _14137_);
  and _73657_ (_28033_, _27349_, _14137_);
  or _73658_ (_28034_, _28033_, _28032_);
  or _73659_ (_28035_, _28034_, _28031_);
  or _73660_ (_28036_, _28035_, _27991_);
  or _73661_ (_28037_, _28036_, _27990_);
  not _73662_ (_28038_, _26413_);
  and _73663_ (_28039_, _26457_, _28038_);
  and _73664_ (_28040_, _28039_, _26547_);
  and _73665_ (_28041_, _28040_, _27362_);
  and _73666_ (_28042_, _28041_, _27598_);
  and _73667_ (property_invalid_sjmp, _28042_, _28037_);
  and _73668_ (_28043_, _27549_, _27072_);
  and _73669_ (_28044_, _28043_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _73670_ (_28045_, _28044_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _73671_ (_28046_, _28045_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _73672_ (_28047_, _28046_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _73673_ (_28048_, _28047_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _73674_ (_28049_, _28048_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _73675_ (_28050_, _28049_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _73676_ (_28051_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _73677_ (_28052_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _73678_ (_28053_, _28052_, _28051_);
  nor _73679_ (_28054_, _28049_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _73680_ (_28055_, _28054_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _73681_ (_28056_, _28055_, _28053_);
  nor _73682_ (_28057_, _28056_, _28050_);
  or _73683_ (_28058_, _28054_, _28050_);
  and _73684_ (_28059_, _28058_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _73685_ (_28060_, _28043_, _27075_);
  nor _73686_ (_28061_, _28045_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _73687_ (_28062_, _28061_, _28060_);
  and _73688_ (_28063_, _28062_, _14121_);
  and _73689_ (_28064_, _27549_, _27071_);
  nor _73690_ (_28065_, _28064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _73691_ (_28066_, _28065_, _28043_);
  and _73692_ (_28067_, _28066_, _27741_);
  nor _73693_ (_28068_, _28066_, _27741_);
  or _73694_ (_28069_, _28068_, _28067_);
  or _73695_ (_28070_, _28069_, _28063_);
  and _73696_ (_28071_, _27549_, _27070_);
  and _73697_ (_28072_, _27549_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _73698_ (_28073_, _28072_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _73699_ (_28074_, _28073_, _28071_);
  nor _73700_ (_28075_, _28074_, _28000_);
  or _73701_ (_28076_, _27551_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand _73702_ (_28077_, _27551_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _73703_ (_28078_, _28077_, _28076_);
  and _73704_ (_28079_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _73705_ (_28080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _73706_ (_28081_, _28080_, _28079_);
  nand _73707_ (_28082_, _28081_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _73708_ (_28083_, _28081_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _73709_ (_28084_, _28083_, _28082_);
  nand _73710_ (_28085_, _28084_, _27313_);
  or _73711_ (_28086_, _27554_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand _73712_ (_28087_, _27554_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _73713_ (_28088_, _28087_, _28086_);
  or _73714_ (_28089_, _28088_, _28085_);
  or _73715_ (_28090_, _28089_, _28078_);
  or _73716_ (_28091_, _28090_, _28075_);
  nor _73717_ (_28092_, _28043_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor _73718_ (_28093_, _28092_, _28044_);
  nor _73719_ (_28094_, _28093_, _14110_);
  and _73720_ (_28095_, _28093_, _14110_);
  or _73721_ (_28096_, _28095_, _28094_);
  or _73722_ (_28097_, _28096_, _28091_);
  nor _73723_ (_28098_, _28071_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _73724_ (_28099_, _28098_, _28064_);
  nor _73725_ (_28100_, _28099_, _27745_);
  and _73726_ (_28101_, _28099_, _27745_);
  or _73727_ (_28102_, _28101_, _28100_);
  or _73728_ (_28103_, _28102_, _28097_);
  nor _73729_ (_28104_, _28062_, _14121_);
  nor _73730_ (_28105_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _73731_ (_28106_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _73732_ (_28107_, _28106_, _28105_);
  or _73733_ (_28108_, _28107_, _28044_);
  nand _73734_ (_28109_, _28107_, _28044_);
  and _73735_ (_28110_, _28109_, _28108_);
  nor _73736_ (_28111_, _27549_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _73737_ (_28112_, _28111_, _28072_);
  nand _73738_ (_28113_, _28112_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or _73739_ (_28114_, _28112_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _73740_ (_28115_, _28114_, _28113_);
  and _73741_ (_28116_, _28074_, _28000_);
  or _73742_ (_28117_, _28116_, _28115_);
  or _73743_ (_28118_, _28117_, _28110_);
  or _73744_ (_28119_, _28118_, _28104_);
  or _73745_ (_28120_, _28119_, _28103_);
  or _73746_ (_28121_, _28120_, _28070_);
  and _73747_ (_28122_, _28060_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _73748_ (_28123_, _28122_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor _73749_ (_28124_, _28123_, _28048_);
  and _73750_ (_28125_, _28124_, _14127_);
  nor _73751_ (_28126_, _28124_, _14127_);
  or _73752_ (_28127_, _28126_, _28125_);
  or _73753_ (_28128_, _28127_, _28121_);
  not _73754_ (_28129_, _28053_);
  and _73755_ (_28130_, _28129_, _28050_);
  nor _73756_ (_28131_, _28046_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _73757_ (_28132_, _28131_, _28047_);
  nor _73758_ (_28133_, _28132_, _14106_);
  and _73759_ (_28134_, _28132_, _14106_);
  or _73760_ (_28135_, _28134_, _28133_);
  nor _73761_ (_28136_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _73762_ (_28137_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _73763_ (_28138_, _28137_, _28136_);
  not _73764_ (_28139_, _28138_);
  and _73765_ (_28140_, _28139_, _28048_);
  nor _73766_ (_28141_, _28139_, _28048_);
  or _73767_ (_28142_, _28141_, _28140_);
  or _73768_ (_28143_, _28142_, _28135_);
  or _73769_ (_28144_, _28143_, _28130_);
  or _73770_ (_28145_, _28144_, _28128_);
  or _73771_ (_28146_, _28145_, _28059_);
  or _73772_ (_28147_, _28146_, _28057_);
  not _73773_ (_28148_, _26502_);
  and _73774_ (_28149_, _28148_, _26369_);
  and _73775_ (_28150_, _28149_, _27984_);
  or _73776_ (_28151_, _28150_, _27365_);
  and _73777_ (_28152_, _28151_, _28039_);
  and _73778_ (_28153_, _26545_, _26413_);
  and _73779_ (_28154_, _28153_, _26369_);
  and _73780_ (_28155_, _26502_, _27366_);
  and _73781_ (_28156_, _28155_, _28154_);
  and _73782_ (_28157_, _26545_, _26502_);
  and _73783_ (_28158_, _27358_, _26236_);
  and _73784_ (_28159_, _28158_, _27361_);
  nand _73785_ (_28160_, _28159_, _27367_);
  nor _73786_ (_28161_, _28160_, _28157_);
  or _73787_ (_28162_, _28161_, _28156_);
  or _73788_ (_28163_, _28162_, _28152_);
  and _73789_ (_28164_, _28163_, _27598_);
  and _73790_ (property_invalid_pcp3, _28164_, _28147_);
  and _73791_ (_28165_, _28148_, _27360_);
  and _73792_ (_28166_, _27364_, _26368_);
  or _73793_ (_28167_, _28166_, _28165_);
  and _73794_ (_28168_, _28167_, _28038_);
  or _73795_ (_28169_, _26413_, _27358_);
  and _73796_ (_28170_, _28169_, _27984_);
  and _73797_ (_28171_, _28170_, _27986_);
  or _73798_ (_28172_, _28154_, _27366_);
  or _73799_ (_28173_, _28172_, _28171_);
  or _73800_ (_28174_, _28173_, _28168_);
  and _73801_ (_28175_, _27984_, _26369_);
  and _73802_ (_28176_, _28153_, _27360_);
  and _73803_ (_28177_, _28176_, _26502_);
  or _73804_ (_28178_, _28177_, _26457_);
  or _73805_ (_28179_, _28178_, _28175_);
  and _73806_ (_28180_, _28179_, _28174_);
  or _73807_ (_28181_, _27987_, _26551_);
  and _73808_ (_28182_, _28181_, _27366_);
  or _73809_ (_28183_, _28182_, _28149_);
  and _73810_ (_28184_, _28183_, _26413_);
  and _73811_ (_28185_, _27358_, _26280_);
  and _73812_ (_28186_, _28185_, _28148_);
  and _73813_ (_28187_, _27986_, _26545_);
  or _73814_ (_28188_, _28187_, _28186_);
  and _73815_ (_28189_, _28188_, _28039_);
  and _73816_ (_28190_, _28157_, _27367_);
  and _73817_ (_28191_, _28190_, _28185_);
  and _73818_ (_28192_, _26546_, _26368_);
  and _73819_ (_28193_, _28192_, _26458_);
  or _73820_ (_28194_, _28193_, _28191_);
  or _73821_ (_28195_, _28194_, _28189_);
  or _73822_ (_28196_, _28195_, _28184_);
  or _73823_ (_28197_, _28196_, _28180_);
  nor _73824_ (_28198_, _27123_, _27745_);
  nor _73825_ (_28199_, _27110_, _14110_);
  or _73826_ (_28200_, _28199_, _28198_);
  and _73827_ (_28201_, _27123_, _27745_);
  and _73828_ (_28202_, _27110_, _14110_);
  or _73829_ (_28203_, _28202_, _28201_);
  or _73830_ (_28204_, _28203_, _28200_);
  and _73831_ (_28205_, _27117_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _73832_ (_28206_, _27130_, _28000_);
  or _73833_ (_28207_, _28206_, _28205_);
  and _73834_ (_28208_, _27130_, _28000_);
  not _73835_ (_28209_, _27098_);
  nor _73836_ (_28210_, _28107_, _28209_);
  or _73837_ (_28211_, _28210_, _28208_);
  or _73838_ (_28212_, _28211_, _28207_);
  and _73839_ (_28213_, _27139_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _73840_ (_28214_, _27139_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _73841_ (_28215_, _28214_, _28213_);
  and _73842_ (_28216_, _27145_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand _73843_ (_28217_, _28081_, _27312_);
  nor _73844_ (_28218_, _27145_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _73845_ (_28219_, _28218_, _28217_);
  or _73846_ (_28220_, _28219_, _28216_);
  or _73847_ (_28221_, _28220_, _28215_);
  nor _73848_ (_28222_, _27136_, _27736_);
  and _73849_ (_28223_, _27136_, _27736_);
  or _73850_ (_28224_, _28223_, _28222_);
  or _73851_ (_28225_, _28224_, _28221_);
  and _73852_ (_28226_, _28107_, _28209_);
  nor _73853_ (_28227_, _27117_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or _73854_ (_28228_, _28227_, _28226_);
  or _73855_ (_28229_, _28228_, _28225_);
  or _73856_ (_28230_, _28229_, _28212_);
  or _73857_ (_28231_, _28230_, _28204_);
  or _73858_ (_28232_, _28231_, _27248_);
  or _73859_ (_28233_, _28232_, _27245_);
  or _73860_ (_28234_, _28233_, _27759_);
  and _73861_ (_28235_, _28234_, _27598_);
  and _73862_ (property_invalid_pcp2, _28235_, _28197_);
  not _73863_ (_28236_, _26235_);
  and _73864_ (_28237_, _26280_, _28236_);
  or _73865_ (_28238_, _28237_, _28158_);
  nor _73866_ (_28239_, _27366_, _26366_);
  and _73867_ (_28240_, _28239_, _28238_);
  and _73868_ (_28241_, _26545_, _28236_);
  and _73869_ (_28242_, _28241_, _26457_);
  or _73870_ (_28243_, _28165_, _28038_);
  or _73871_ (_28244_, _28243_, _28242_);
  or _73872_ (_28245_, _28244_, _28186_);
  or _73873_ (_28246_, _28245_, _28240_);
  and _73874_ (_28247_, _26551_, _26547_);
  and _73875_ (_28248_, _27363_, _27360_);
  and _73876_ (_28249_, _28248_, _26502_);
  or _73877_ (_28250_, _28159_, _26413_);
  or _73878_ (_28251_, _28250_, _28249_);
  or _73879_ (_28252_, _28251_, _28247_);
  and _73880_ (_28253_, _28252_, _28246_);
  and _73881_ (_28254_, _28176_, _26457_);
  and _73882_ (_28255_, _27359_, _26548_);
  nor _73883_ (_28256_, _27363_, _26502_);
  and _73884_ (_28257_, _28256_, _26368_);
  and _73885_ (_28258_, _28257_, _28039_);
  or _73886_ (_28259_, _28258_, _28255_);
  or _73887_ (_28260_, _28259_, _28254_);
  or _73888_ (_28261_, _28185_, _27360_);
  nand _73889_ (_28262_, _27984_, _26501_);
  nor _73890_ (_28263_, _28262_, _27360_);
  or _73891_ (_28264_, _28263_, _26458_);
  and _73892_ (_28265_, _28264_, _28261_);
  and _73893_ (_28266_, _28248_, _27366_);
  and _73894_ (_28267_, _28237_, _27985_);
  or _73895_ (_28268_, _28267_, _28266_);
  or _73896_ (_28269_, _28268_, _28265_);
  or _73897_ (_28270_, _28269_, _28260_);
  or _73898_ (_28271_, _28270_, _28253_);
  nor _73899_ (_28272_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _73900_ (_28273_, _27072_, _21597_);
  and _73901_ (_28274_, _28273_, _27075_);
  or _73902_ (_28275_, _28274_, _28272_);
  nor _73903_ (_28276_, _28275_, _27100_);
  nor _73904_ (_28277_, _28276_, _14121_);
  and _73905_ (_28278_, _28273_, _27076_);
  and _73906_ (_28279_, _28278_, _16238_);
  nor _73907_ (_28280_, _28278_, _16238_);
  or _73908_ (_28281_, _28280_, _28279_);
  nand _73909_ (_28282_, _28281_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _73910_ (_28283_, _28281_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _73911_ (_28284_, _28283_, _28282_);
  or _73912_ (_28285_, _28284_, _28277_);
  and _73913_ (_28286_, _27078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nand _73914_ (_28287_, _28286_, _28138_);
  or _73915_ (_28288_, _28286_, _28138_);
  and _73916_ (_28289_, _28288_, _28287_);
  and _73917_ (_28290_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5], _16190_);
  and _73918_ (_28291_, _27130_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _73919_ (_28292_, _28291_, _28290_);
  or _73920_ (_28293_, _28292_, _28000_);
  nand _73921_ (_28294_, _28292_, _28000_);
  and _73922_ (_28295_, _28294_, _28293_);
  or _73923_ (_28296_, _28295_, _28289_);
  or _73924_ (_28297_, _28296_, _28285_);
  and _73925_ (_28298_, _27114_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _73926_ (_28299_, _27070_, _21597_);
  nor _73927_ (_28300_, _28299_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _73928_ (_28301_, _28300_, _28298_);
  and _73929_ (_28302_, _28301_, _27745_);
  nor _73930_ (_28303_, _28301_, _27745_);
  and _73931_ (_28304_, _21602_, _27376_);
  nor _73932_ (_28305_, _21602_, _27376_);
  or _73933_ (_28306_, _28305_, _28084_);
  or _73934_ (_28307_, _28306_, _28304_);
  or _73935_ (_28308_, _28307_, _28303_);
  or _73936_ (_28309_, _28308_, _28302_);
  nor _73937_ (_28310_, _28298_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _73938_ (_28311_, _28310_, _28273_);
  nor _73939_ (_28312_, _28311_, _27741_);
  and _73940_ (_28313_, _21599_, _27369_);
  nor _73941_ (_28314_, _21599_, _27369_);
  nor _73942_ (_28315_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _73943_ (_28316_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _73944_ (_28317_, _28316_, _28315_);
  not _73945_ (_28318_, _28317_);
  nor _73946_ (_28319_, _28318_, _21597_);
  and _73947_ (_28320_, _28318_, _21597_);
  or _73948_ (_28321_, _28320_, _27312_);
  or _73949_ (_28322_, _28321_, _28319_);
  or _73950_ (_28323_, _28322_, _28314_);
  or _73951_ (_28324_, _28323_, _28313_);
  or _73952_ (_28325_, _28324_, _28312_);
  nor _73953_ (_28326_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _73954_ (_28327_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _73955_ (_28328_, _28327_, _28326_);
  or _73956_ (_28329_, _28328_, _28274_);
  nand _73957_ (_28330_, _28328_, _28274_);
  and _73958_ (_28331_, _28330_, _28329_);
  and _73959_ (_28332_, _28311_, _27741_);
  or _73960_ (_28333_, _28332_, _28331_);
  or _73961_ (_28334_, _28333_, _28325_);
  or _73962_ (_28335_, _28334_, _28309_);
  and _73963_ (_28336_, _28276_, _14121_);
  nand _73964_ (_28337_, _28273_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _73965_ (_28338_, _28337_, _28107_);
  and _73966_ (_28339_, _28210_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _73967_ (_28340_, _28339_, _28338_);
  or _73968_ (_28341_, _28273_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _73969_ (_28342_, _28341_, _28337_);
  and _73970_ (_28343_, _28342_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _73971_ (_28344_, _28342_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _73972_ (_28345_, _28344_, _28343_);
  or _73973_ (_28346_, _28345_, _28340_);
  or _73974_ (_28347_, _28346_, _28336_);
  or _73975_ (_28348_, _28347_, _28335_);
  or _73976_ (_28349_, _28348_, _28297_);
  and _73977_ (_28350_, _27080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _73978_ (_28351_, _28350_, _28053_);
  nand _73979_ (_28352_, _28350_, _28053_);
  and _73980_ (_28353_, _28352_, _28351_);
  nand _73981_ (_28354_, _27079_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _73982_ (_28355_, _28354_, _16246_);
  nor _73983_ (_28356_, _28355_, _28350_);
  and _73984_ (_28357_, _28356_, _14137_);
  nor _73985_ (_28358_, _28356_, _14137_);
  or _73986_ (_28359_, _28358_, _28357_);
  or _73987_ (_28360_, _28359_, _28353_);
  or _73988_ (_28361_, _28360_, _28349_);
  and _73989_ (_28362_, _28361_, _27598_);
  and _73990_ (property_invalid_pcp1, _28362_, _28271_);
  and _73991_ (_28363_, _26138_, pc_change_r);
  and _73992_ (_28364_, _28363_, _27596_);
  and _73993_ (_28365_, acc_reg[0], acc_reg[1]);
  and _73994_ (_28366_, _28365_, acc_reg[2]);
  and _73995_ (_28367_, _28366_, acc_reg[3]);
  and _73996_ (_28368_, _28367_, acc_reg[4]);
  and _73997_ (_28369_, _28368_, acc_reg[5]);
  and _73998_ (_28370_, _28369_, acc_reg[6]);
  nor _73999_ (_28371_, acc_reg[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _74000_ (_28372_, acc_reg[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _74001_ (_28373_, _28372_, _28371_);
  nor _74002_ (_28374_, _28369_, acc_reg[6]);
  nor _74003_ (_28375_, _28374_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _74004_ (_28376_, _28375_, _28373_);
  nor _74005_ (_28377_, _28376_, _28370_);
  not _74006_ (_28378_, _28373_);
  and _74007_ (_28379_, _28378_, _28370_);
  nor _74008_ (_28380_, _28368_, acc_reg[5]);
  nor _74009_ (_28381_, _28380_, _28369_);
  nor _74010_ (_28382_, _28381_, _33948_);
  and _74011_ (_28383_, _28381_, _33948_);
  or _74012_ (_28384_, _28383_, _28382_);
  or _74013_ (_28385_, _28384_, _28379_);
  or _74014_ (_28386_, _28374_, _28370_);
  and _74015_ (_28387_, _28386_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _74016_ (_28388_, _28366_, acc_reg[3]);
  nor _74017_ (_28389_, _28388_, _28367_);
  and _74018_ (_28390_, _28389_, _34032_);
  nor _74019_ (_28391_, _28389_, _34032_);
  or _74020_ (_28392_, _28391_, _28390_);
  and _74021_ (_28393_, acc_reg[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _74022_ (_28394_, acc_reg[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _74023_ (_28395_, _28394_, _28393_);
  not _74024_ (_28396_, acc_reg[0]);
  and _74025_ (_28397_, _28396_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nand _74026_ (_28398_, _28397_, _28395_);
  or _74027_ (_28399_, _28396_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _74028_ (_28400_, _28399_, _28395_);
  and _74029_ (_28401_, _28400_, _28398_);
  nor _74030_ (_28402_, _28365_, acc_reg[2]);
  nor _74031_ (_28403_, _28402_, _28366_);
  nor _74032_ (_28404_, _28403_, _34059_);
  and _74033_ (_28405_, _28403_, _34059_);
  or _74034_ (_28406_, _28405_, _28404_);
  or _74035_ (_28407_, _28406_, _28401_);
  or _74036_ (_28408_, _28407_, _28392_);
  nor _74037_ (_28409_, _28367_, acc_reg[4]);
  nor _74038_ (_28410_, _28409_, _28368_);
  nor _74039_ (_28411_, _28410_, _33984_);
  and _74040_ (_28412_, _28410_, _33984_);
  or _74041_ (_28413_, _28412_, _28411_);
  or _74042_ (_28414_, _28413_, _28408_);
  or _74043_ (_28415_, _28414_, _28387_);
  or _74044_ (_28416_, _28415_, _28385_);
  or _74045_ (_28417_, _28416_, _28377_);
  and _74046_ (_28418_, _28417_, pc_inc_acc_r);
  and _74047_ (property_invalid_inc_acc, _28418_, _28364_);
  not _74048_ (_28419_, op1_out_r[0]);
  and _74049_ (_28420_, _28419_, op1_out_r[1]);
  and _74050_ (_28421_, op1_out_r[2], op1_out_r[3]);
  and _74051_ (_28422_, _28421_, _28420_);
  not _74052_ (_28423_, op1_out_r[5]);
  and _74053_ (_28424_, op1_out_r[4], _28423_);
  and _74054_ (_28425_, op1_out_r[7], op1_out_r[6]);
  and _74055_ (_28426_, _28425_, _28424_);
  and _74056_ (_28427_, _28426_, _28422_);
  nor _74057_ (_28428_, _28419_, op1_out_r[1]);
  not _74058_ (_28429_, op1_out_r[3]);
  and _74059_ (_28430_, op1_out_r[2], _28429_);
  and _74060_ (_28431_, _28430_, _28428_);
  and _74061_ (_28432_, _28431_, _28426_);
  nor _74062_ (_28433_, _28432_, _28427_);
  and _74063_ (_28434_, _28428_, _28421_);
  and _74064_ (_28435_, _28434_, _28426_);
  nor _74065_ (_28436_, op1_out_r[2], op1_out_r[3]);
  and _74066_ (_28437_, _28436_, _28428_);
  nor _74067_ (_28438_, op1_out_r[4], op1_out_r[5]);
  not _74068_ (_28439_, op1_out_r[7]);
  and _74069_ (_28440_, _28439_, op1_out_r[6]);
  and _74070_ (_28441_, _28440_, _28438_);
  and _74071_ (_28442_, _28441_, _28437_);
  nor _74072_ (_28443_, _28442_, _28435_);
  and _74073_ (_28444_, _28443_, _28433_);
  and _74074_ (_28445_, op1_out_r[0], op1_out_r[1]);
  and _74075_ (_28446_, _28445_, _28421_);
  and _74076_ (_28447_, _28438_, _28425_);
  and _74077_ (_28448_, _28447_, _28446_);
  and _74078_ (_28449_, _28436_, _28420_);
  and _74079_ (_28450_, _28449_, _28426_);
  nor _74080_ (_28451_, _28450_, _28448_);
  and _74081_ (_28452_, _28440_, _28424_);
  and _74082_ (_28453_, _28452_, _28446_);
  nor _74083_ (_28454_, op1_out_r[4], _28423_);
  and _74084_ (_28455_, _28454_, _28440_);
  and _74085_ (_28456_, _28455_, _28449_);
  nor _74086_ (_28457_, _28456_, _28453_);
  and _74087_ (_28458_, _28457_, _28451_);
  and _74088_ (_28459_, _28458_, _28444_);
  nor _74089_ (_28460_, _28439_, op1_out_r[6]);
  and _74090_ (_28461_, _28460_, _28454_);
  and _74091_ (_28462_, _28461_, _28431_);
  and _74092_ (_28463_, _28430_, _28420_);
  and _74093_ (_28464_, _28463_, _28461_);
  nor _74094_ (_28465_, _28464_, _28462_);
  and _74095_ (_28466_, op1_out_r[4], op1_out_r[5]);
  and _74096_ (_28467_, _28466_, _28460_);
  and _74097_ (_28468_, _28467_, _28434_);
  nor _74098_ (_28469_, op1_out_r[2], _28429_);
  and _74099_ (_28470_, _28469_, _28445_);
  and _74100_ (_28471_, _28470_, _28467_);
  nor _74101_ (_28472_, _28471_, _28468_);
  and _74102_ (_28473_, _28472_, _28465_);
  and _74103_ (_28474_, _28467_, _28463_);
  nor _74104_ (_28475_, op1_out_r[0], op1_out_r[1]);
  and _74105_ (_28476_, _28475_, _28469_);
  and _74106_ (_28477_, _28476_, _28467_);
  nor _74107_ (_28478_, _28477_, _28474_);
  and _74108_ (_28479_, _28445_, _28436_);
  and _74109_ (_28480_, _28479_, _28426_);
  and _74110_ (_28481_, _28463_, _28426_);
  nor _74111_ (_28482_, _28481_, _28480_);
  and _74112_ (_28483_, _28482_, _28478_);
  and _74113_ (_28484_, _28483_, _28473_);
  and _74114_ (_28485_, _28484_, _28459_);
  and _74115_ (_28486_, _28467_, _28437_);
  and _74116_ (_28487_, _28445_, _28430_);
  and _74117_ (_28488_, _28487_, _28467_);
  nor _74118_ (_28489_, _28488_, _28486_);
  and _74119_ (_28490_, _28475_, _28436_);
  and _74120_ (_28491_, _28490_, _28467_);
  and _74121_ (_28492_, _28469_, _28420_);
  and _74122_ (_28493_, _28492_, _28467_);
  nor _74123_ (_28494_, _28493_, _28491_);
  and _74124_ (_28495_, _28494_, _28489_);
  and _74125_ (_28496_, _28467_, _28449_);
  and _74126_ (_28497_, _28461_, _28446_);
  nor _74127_ (_28498_, _28497_, _28496_);
  and _74128_ (_28499_, _28454_, _28425_);
  and _74129_ (_28500_, _28499_, _28479_);
  and _74130_ (_28501_, _28446_, _28426_);
  nor _74131_ (_28502_, _28501_, _28500_);
  and _74132_ (_28503_, _28502_, _28498_);
  and _74133_ (_28504_, _28503_, _28495_);
  and _74134_ (_28505_, _28466_, _28440_);
  and _74135_ (_28506_, _28505_, _28463_);
  and _74136_ (_28507_, _28505_, _28431_);
  nor _74137_ (_28508_, _28507_, _28506_);
  and _74138_ (_28509_, _28475_, _28430_);
  and _74139_ (_28510_, _28509_, _28467_);
  and _74140_ (_28511_, _28509_, _28505_);
  nor _74141_ (_28512_, _28511_, _28510_);
  and _74142_ (_28513_, _28512_, _28508_);
  and _74143_ (_28514_, _28475_, _28421_);
  and _74144_ (_28515_, _28514_, _28426_);
  and _74145_ (_28516_, _28470_, _28426_);
  nor _74146_ (_28517_, _28516_, _28515_);
  and _74147_ (_28518_, _28467_, _28431_);
  and _74148_ (_28519_, _28467_, _28422_);
  nor _74149_ (_28520_, _28519_, _28518_);
  and _74150_ (_28521_, _28520_, _28517_);
  and _74151_ (_28522_, _28521_, _28513_);
  and _74152_ (_28523_, _28522_, _28504_);
  and _74153_ (_28524_, _28523_, _28485_);
  and _74154_ (_28525_, _28460_, _28438_);
  and _74155_ (_28526_, _28525_, _28437_);
  nor _74156_ (_28527_, op1_out_r[7], op1_out_r[6]);
  and _74157_ (_28528_, _28527_, _28454_);
  and _74158_ (_28529_, _28528_, _28431_);
  nor _74159_ (_28530_, _28529_, _28526_);
  and _74160_ (_28531_, _28525_, _28470_);
  and _74161_ (_28532_, _28525_, _28490_);
  nor _74162_ (_28533_, _28532_, _28531_);
  and _74163_ (_28534_, _28533_, _28530_);
  and _74164_ (_28535_, _28455_, _28431_);
  and _74165_ (_28536_, _28509_, _28455_);
  nor _74166_ (_28537_, _28536_, _28535_);
  and _74167_ (_28538_, _28527_, _28438_);
  and _74168_ (_28539_, _28538_, _28431_);
  and _74169_ (_28540_, _28538_, _28509_);
  nor _74170_ (_28541_, _28540_, _28539_);
  and _74171_ (_28542_, _28541_, _28537_);
  and _74172_ (_28543_, _28542_, _28534_);
  and _74173_ (_28544_, _28466_, _28425_);
  and _74174_ (_28545_, _28544_, _28509_);
  and _74175_ (_28546_, _28544_, _28479_);
  nor _74176_ (_28547_, _28546_, _28545_);
  and _74177_ (_28548_, _28525_, _28422_);
  and _74178_ (_28549_, _28460_, _28424_);
  and _74179_ (_28550_, _28549_, _28490_);
  nor _74180_ (_28551_, _28550_, _28548_);
  and _74181_ (_28552_, _28551_, _28547_);
  and _74182_ (_28553_, _28525_, _28514_);
  and _74183_ (_28554_, _28469_, _28428_);
  and _74184_ (_28555_, _28554_, _28528_);
  nor _74185_ (_28556_, _28555_, _28553_);
  and _74186_ (_28557_, _28549_, _28437_);
  and _74187_ (_28558_, _28525_, _28449_);
  nor _74188_ (_28559_, _28558_, _28557_);
  and _74189_ (_28560_, _28559_, _28556_);
  and _74190_ (_28561_, _28560_, _28552_);
  and _74191_ (_28562_, _28561_, _28543_);
  and _74192_ (_28563_, _28499_, _28434_);
  and _74193_ (_28564_, _28499_, _28422_);
  nor _74194_ (_28565_, _28564_, _28563_);
  and _74195_ (_28566_, _28514_, _28499_);
  and _74196_ (_28567_, _28525_, _28463_);
  nor _74197_ (_28568_, _28567_, _28566_);
  and _74198_ (_28569_, _28568_, _28565_);
  and _74199_ (_28570_, _28479_, _28461_);
  and _74200_ (_28571_, _28525_, _28509_);
  nor _74201_ (_28572_, _28571_, _28570_);
  and _74202_ (_28573_, _28554_, _28549_);
  and _74203_ (_28574_, _28505_, _28446_);
  nor _74204_ (_28575_, _28574_, _28573_);
  and _74205_ (_28576_, _28575_, _28572_);
  and _74206_ (_28577_, _28576_, _28569_);
  and _74207_ (_28578_, _28490_, _28461_);
  and _74208_ (_28579_, _28527_, _28424_);
  and _74209_ (_28580_, _28579_, _28446_);
  nor _74210_ (_28581_, _28580_, _28578_);
  and _74211_ (_28582_, _28538_, _28463_);
  and _74212_ (_28583_, _28479_, _28455_);
  nor _74213_ (_28584_, _28583_, _28582_);
  and _74214_ (_28585_, _28584_, _28581_);
  and _74215_ (_28586_, _28525_, _28479_);
  and _74216_ (_28587_, _28525_, _28431_);
  nor _74217_ (_28588_, _28587_, _28586_);
  and _74218_ (_28589_, _28461_, _28437_);
  and _74219_ (_28590_, _28487_, _28461_);
  nor _74220_ (_28591_, _28590_, _28589_);
  and _74221_ (_28592_, _28591_, _28588_);
  and _74222_ (_28593_, _28592_, _28585_);
  and _74223_ (_28594_, _28593_, _28577_);
  and _74224_ (_28595_, _28594_, _28562_);
  and _74225_ (_28596_, _28595_, _28524_);
  and _74226_ (_28597_, _28528_, _28487_);
  and _74227_ (_28598_, _28527_, _28466_);
  and _74228_ (_28599_, _28598_, _28554_);
  nor _74229_ (_28600_, _28599_, _28597_);
  and _74230_ (_28601_, _28505_, _28476_);
  and _74231_ (_28602_, _28505_, _28422_);
  nor _74232_ (_28603_, _28602_, _28601_);
  and _74233_ (_28604_, _28603_, _28600_);
  and _74234_ (_28605_, _28598_, _28476_);
  and _74235_ (_28606_, _28598_, _28422_);
  nor _74236_ (_28607_, _28606_, _28605_);
  and _74237_ (_28608_, _28528_, _28492_);
  and _74238_ (_28609_, _28528_, _28476_);
  nor _74239_ (_28610_, _28609_, _28608_);
  and _74240_ (_28611_, _28610_, _28607_);
  and _74241_ (_28612_, _28611_, _28604_);
  and _74242_ (_28613_, _28554_, _28467_);
  and _74243_ (_28614_, _28455_, _28422_);
  nor _74244_ (_28615_, _28614_, _28613_);
  and _74245_ (_28616_, _28499_, _28431_);
  and _74246_ (_28617_, _28455_, _28434_);
  nor _74247_ (_28618_, _28617_, _28616_);
  and _74248_ (_28619_, _28618_, _28615_);
  and _74249_ (_28620_, _28505_, _28492_);
  and _74250_ (_28621_, _28598_, _28492_);
  nor _74251_ (_28622_, _28621_, _28620_);
  and _74252_ (_28623_, _28505_, _28487_);
  and _74253_ (_28624_, _28598_, _28487_);
  nor _74254_ (_28625_, _28624_, _28623_);
  and _74255_ (_28626_, _28625_, _28622_);
  and _74256_ (_28627_, _28626_, _28619_);
  and _74257_ (_28628_, _28627_, _28612_);
  and _74258_ (_28629_, _28549_, _28422_);
  and _74259_ (_28630_, _28549_, _28434_);
  nor _74260_ (_28631_, _28630_, _28629_);
  and _74261_ (_28632_, _28549_, _28470_);
  and _74262_ (_28633_, _28549_, _28514_);
  nor _74263_ (_28634_, _28633_, _28632_);
  and _74264_ (_28635_, _28634_, _28631_);
  and _74265_ (_28636_, _28461_, _28422_);
  and _74266_ (_28637_, _28461_, _28434_);
  nor _74267_ (_28638_, _28637_, _28636_);
  and _74268_ (_28639_, _28470_, _28461_);
  and _74269_ (_28640_, _28514_, _28461_);
  nor _74270_ (_28641_, _28640_, _28639_);
  and _74271_ (_28642_, _28641_, _28638_);
  and _74272_ (_28643_, _28642_, _28635_);
  and _74273_ (_28644_, _28544_, _28487_);
  and _74274_ (_28645_, _28544_, _28476_);
  nor _74275_ (_28646_, _28645_, _28644_);
  and _74276_ (_28647_, _28452_, _28431_);
  and _74277_ (_28648_, _28479_, _28452_);
  nor _74278_ (_28649_, _28648_, _28647_);
  and _74279_ (_28650_, _28649_, _28646_);
  and _74280_ (_28651_, _28549_, _28487_);
  and _74281_ (_28652_, _28549_, _28476_);
  nor _74282_ (_28653_, _28652_, _28651_);
  and _74283_ (_28654_, _28487_, _28441_);
  and _74284_ (_28655_, _28549_, _28492_);
  nor _74285_ (_28656_, _28655_, _28654_);
  and _74286_ (_28657_, _28656_, _28653_);
  and _74287_ (_28658_, _28657_, _28650_);
  and _74288_ (_28659_, _28658_, _28643_);
  and _74289_ (_28660_, _28659_, _28628_);
  and _74290_ (_28661_, _28452_, _28449_);
  and _74291_ (_28662_, _28505_, _28449_);
  nor _74292_ (_28663_, _28662_, _28661_);
  and _74293_ (_28664_, _28441_, _28422_);
  and _74294_ (_28665_, _28455_, _28446_);
  nor _74295_ (_28666_, _28665_, _28664_);
  and _74296_ (_28667_, _28666_, _28663_);
  and _74297_ (_28668_, _28452_, _28437_);
  and _74298_ (_28669_, _28505_, _28479_);
  nor _74299_ (_28670_, _28669_, _28668_);
  and _74300_ (_28671_, _28509_, _28452_);
  and _74301_ (_28672_, _28490_, _28452_);
  nor _74302_ (_28673_, _28672_, _28671_);
  and _74303_ (_28674_, _28673_, _28670_);
  and _74304_ (_28675_, _28674_, _28667_);
  and _74305_ (_28676_, _28598_, _28437_);
  and _74306_ (_28677_, _28554_, _28447_);
  nor _74307_ (_28678_, _28677_, _28676_);
  and _74308_ (_28679_, _28554_, _28499_);
  and _74309_ (_28680_, _28447_, _28434_);
  nor _74310_ (_28681_, _28680_, _28679_);
  and _74311_ (_28682_, _28681_, _28678_);
  and _74312_ (_28683_, _28490_, _28455_);
  and _74313_ (_28684_, _28455_, _28437_);
  nor _74314_ (_28685_, _28684_, _28683_);
  and _74315_ (_28686_, _28598_, _28449_);
  and _74316_ (_28687_, _28598_, _28490_);
  nor _74317_ (_28688_, _28687_, _28686_);
  and _74318_ (_28689_, _28688_, _28685_);
  and _74319_ (_28690_, _28689_, _28682_);
  and _74320_ (_28691_, _28690_, _28675_);
  and _74321_ (_28692_, _28499_, _28449_);
  and _74322_ (_28693_, _28499_, _28437_);
  nor _74323_ (_28694_, _28693_, _28692_);
  and _74324_ (_28695_, _28449_, _28447_);
  and _74325_ (_28696_, _28509_, _28447_);
  nor _74326_ (_28697_, _28696_, _28695_);
  and _74327_ (_28698_, _28697_, _28694_);
  and _74328_ (_28699_, _28499_, _28490_);
  and _74329_ (_28700_, _28499_, _28492_);
  nor _74330_ (_28701_, _28700_, _28699_);
  and _74331_ (_28702_, _28463_, _28447_);
  and _74332_ (_28703_, _28499_, _28476_);
  nor _74333_ (_28704_, _28703_, _28702_);
  and _74334_ (_28705_, _28704_, _28701_);
  and _74335_ (_28706_, _28705_, _28698_);
  and _74336_ (_28707_, _28579_, _28449_);
  and _74337_ (_28708_, _28492_, _28447_);
  nor _74338_ (_28709_, _28708_, _28707_);
  and _74339_ (_28710_, _28579_, _28463_);
  and _74340_ (_28711_, _28579_, _28509_);
  nor _74341_ (_28712_, _28711_, _28710_);
  and _74342_ (_28713_, _28712_, _28709_);
  and _74343_ (_28714_, _28487_, _28447_);
  and _74344_ (_28715_, _28470_, _28447_);
  nor _74345_ (_28716_, _28715_, _28714_);
  and _74346_ (_28717_, _28447_, _28437_);
  and _74347_ (_28718_, _28476_, _28447_);
  nor _74348_ (_28719_, _28718_, _28717_);
  and _74349_ (_28720_, _28719_, _28716_);
  and _74350_ (_28721_, _28720_, _28713_);
  and _74351_ (_28722_, _28721_, _28706_);
  and _74352_ (_28723_, _28722_, _28691_);
  and _74353_ (_28724_, _28723_, _28660_);
  and _74354_ (_28725_, _28724_, _28596_);
  and _74355_ (_28726_, _28538_, _28476_);
  and _74356_ (_28727_, _28538_, _28492_);
  nor _74357_ (_28728_, _28727_, _28726_);
  and _74358_ (_28729_, _28579_, _28554_);
  and _74359_ (_28730_, _28538_, _28487_);
  nor _74360_ (_28731_, _28730_, _28729_);
  and _74361_ (_28732_, _28731_, _28728_);
  and _74362_ (_28733_, _28598_, _28446_);
  and _74363_ (_28734_, _28509_, _28441_);
  nor _74364_ (_28735_, _28734_, _28733_);
  and _74365_ (_28736_, _28449_, _28441_);
  and _74366_ (_28737_, _28490_, _28441_);
  nor _74367_ (_28738_, _28737_, _28736_);
  and _74368_ (_28739_, _28738_, _28735_);
  and _74369_ (_28740_, _28739_, _28732_);
  and _74370_ (_28741_, _28528_, _28446_);
  and _74371_ (_28742_, _28528_, _28437_);
  nor _74372_ (_28743_, _28742_, _28741_);
  and _74373_ (_28744_, _28598_, _28431_);
  and _74374_ (_28745_, _28598_, _28479_);
  nor _74375_ (_28746_, _28745_, _28744_);
  and _74376_ (_28747_, _28746_, _28743_);
  and _74377_ (_28748_, _28487_, _28452_);
  and _74378_ (_28749_, _28441_, _28431_);
  nor _74379_ (_28750_, _28749_, _28748_);
  and _74380_ (_28751_, _28479_, _28441_);
  and _74381_ (_28752_, _28463_, _28441_);
  nor _74382_ (_28753_, _28752_, _28751_);
  and _74383_ (_28754_, _28753_, _28750_);
  and _74384_ (_28755_, _28754_, _28747_);
  and _74385_ (_28756_, _28755_, _28740_);
  and _74386_ (_28757_, _28470_, _28452_);
  and _74387_ (_28758_, _28514_, _28452_);
  nor _74388_ (_28759_, _28758_, _28757_);
  and _74389_ (_28760_, _28549_, _28509_);
  and _74390_ (_28761_, _28554_, _28538_);
  nor _74391_ (_28762_, _28761_, _28760_);
  and _74392_ (_28763_, _28762_, _28759_);
  and _74393_ (_28764_, _28525_, _28434_);
  and _74394_ (_28765_, _28549_, _28463_);
  nor _74395_ (_28766_, _28765_, _28764_);
  and _74396_ (_28767_, _28549_, _28479_);
  and _74397_ (_28768_, _28549_, _28431_);
  nor _74398_ (_28769_, _28768_, _28767_);
  and _74399_ (_28770_, _28769_, _28766_);
  and _74400_ (_28771_, _28770_, _28763_);
  and _74401_ (_28772_, _28538_, _28422_);
  and _74402_ (_28773_, _28476_, _28452_);
  nor _74403_ (_28774_, _28773_, _28772_);
  and _74404_ (_28775_, _28538_, _28434_);
  and _74405_ (_28776_, _28538_, _28470_);
  nor _74406_ (_28777_, _28776_, _28775_);
  and _74407_ (_28778_, _28777_, _28774_);
  and _74408_ (_28779_, _28554_, _28452_);
  and _74409_ (_28780_, _28492_, _28452_);
  nor _74410_ (_28781_, _28780_, _28779_);
  and _74411_ (_28782_, _28452_, _28422_);
  and _74412_ (_28783_, _28452_, _28434_);
  nor _74413_ (_28784_, _28783_, _28782_);
  and _74414_ (_28785_, _28784_, _28781_);
  and _74415_ (_28786_, _28785_, _28778_);
  and _74416_ (_28787_, _28786_, _28771_);
  and _74417_ (_28788_, _28787_, _28756_);
  and _74418_ (_28789_, _28492_, _28455_);
  and _74419_ (_28790_, _28598_, _28470_);
  nor _74420_ (_28791_, _28790_, _28789_);
  and _74421_ (_28792_, _28554_, _28505_);
  and _74422_ (_28793_, _28487_, _28455_);
  nor _74423_ (_28794_, _28793_, _28792_);
  and _74424_ (_28795_, _28794_, _28791_);
  and _74425_ (_28796_, _28554_, _28426_);
  and _74426_ (_28797_, _28514_, _28467_);
  nor _74427_ (_28798_, _28797_, _28796_);
  and _74428_ (_28799_, _28479_, _28467_);
  and _74429_ (_28800_, _28476_, _28455_);
  nor _74430_ (_28801_, _28800_, _28799_);
  and _74431_ (_28802_, _28801_, _28798_);
  and _74432_ (_28803_, _28437_, _28426_);
  and _74433_ (_28804_, _28490_, _28426_);
  nor _74434_ (_28805_, _28804_, _28803_);
  and _74435_ (_28806_, _28492_, _28426_);
  and _74436_ (_28807_, _28476_, _28426_);
  nor _74437_ (_28808_, _28807_, _28806_);
  and _74438_ (_28809_, _28808_, _28805_);
  and _74439_ (_28810_, _28809_, _28802_);
  and _74440_ (_28811_, _28810_, _28795_);
  and _74441_ (_28812_, _28505_, _28437_);
  and _74442_ (_28813_, _28505_, _28490_);
  nor _74443_ (_28814_, _28813_, _28812_);
  and _74444_ (_28815_, _28441_, _28434_);
  and _74445_ (_28816_, _28538_, _28436_);
  nor _74446_ (_28817_, _28816_, _28815_);
  and _74447_ (_28818_, _28817_, _28814_);
  and _74448_ (_28819_, _28598_, _28509_);
  and _74449_ (_28820_, _28528_, _28449_);
  nor _74450_ (_28821_, _28820_, _28819_);
  and _74451_ (_28822_, _28579_, _28479_);
  and _74452_ (_28823_, _28463_, _28455_);
  nor _74453_ (_28824_, _28823_, _28822_);
  and _74454_ (_28825_, _28824_, _28821_);
  and _74455_ (_28826_, _28825_, _28818_);
  and _74456_ (_28827_, _28598_, _28463_);
  and _74457_ (_28828_, _28528_, _28490_);
  nor _74458_ (_28829_, _28828_, _28827_);
  and _74459_ (_28830_, _28487_, _28426_);
  and _74460_ (_28831_, _28509_, _28426_);
  nor _74461_ (_28832_, _28831_, _28830_);
  and _74462_ (_28833_, _28832_, _28829_);
  and _74463_ (_28834_, _28579_, _28437_);
  and _74464_ (_28835_, _28579_, _28490_);
  nor _74465_ (_28836_, _28835_, _28834_);
  and _74466_ (_28837_, _28538_, _28446_);
  and _74467_ (_28838_, _28579_, _28431_);
  nor _74468_ (_28839_, _28838_, _28837_);
  and _74469_ (_28840_, _28839_, _28836_);
  and _74470_ (_28841_, _28840_, _28833_);
  and _74471_ (_28842_, _28841_, _28826_);
  and _74472_ (_28843_, _28842_, _28811_);
  and _74473_ (_28844_, _28843_, _28788_);
  and _74474_ (_28845_, _28544_, _28422_);
  and _74475_ (_28846_, _28544_, _28449_);
  nor _74476_ (_28847_, _28846_, _28845_);
  and _74477_ (_28848_, _28544_, _28434_);
  and _74478_ (_28849_, _28528_, _28422_);
  nor _74479_ (_28850_, _28849_, _28848_);
  and _74480_ (_28851_, _28850_, _28847_);
  and _74481_ (_28852_, _28544_, _28514_);
  and _74482_ (_28853_, _28499_, _28446_);
  nor _74483_ (_28854_, _28853_, _28852_);
  and _74484_ (_28855_, _28544_, _28470_);
  and _74485_ (_28856_, _28544_, _28490_);
  nor _74486_ (_28857_, _28856_, _28855_);
  and _74487_ (_28858_, _28857_, _28854_);
  and _74488_ (_28859_, _28858_, _28851_);
  and _74489_ (_28860_, _28492_, _28461_);
  and _74490_ (_28861_, _28554_, _28461_);
  nor _74491_ (_28862_, _28861_, _28860_);
  and _74492_ (_28863_, _28598_, _28434_);
  and _74493_ (_28864_, _28598_, _28514_);
  nor _74494_ (_28865_, _28864_, _28863_);
  and _74495_ (_28866_, _28865_, _28862_);
  and _74496_ (_28867_, _28528_, _28434_);
  and _74497_ (_28868_, _28528_, _28470_);
  nor _74498_ (_28869_, _28868_, _28867_);
  and _74499_ (_28870_, _28528_, _28514_);
  and _74500_ (_28871_, _28554_, _28455_);
  nor _74501_ (_28872_, _28871_, _28870_);
  and _74502_ (_28873_, _28872_, _28869_);
  and _74503_ (_28874_, _28873_, _28866_);
  and _74504_ (_28875_, _28874_, _28859_);
  and _74505_ (_28876_, _28514_, _28447_);
  and _74506_ (_28877_, _28514_, _28455_);
  nor _74507_ (_28878_, _28877_, _28876_);
  and _74508_ (_28879_, _28479_, _28447_);
  and _74509_ (_28880_, _28447_, _28422_);
  nor _74510_ (_28881_, _28880_, _28879_);
  and _74511_ (_28882_, _28881_, _28878_);
  and _74512_ (_28883_, _28514_, _28505_);
  and _74513_ (_28884_, _28470_, _28455_);
  nor _74514_ (_28885_, _28884_, _28883_);
  and _74515_ (_28886_, _28505_, _28434_);
  and _74516_ (_28887_, _28505_, _28470_);
  nor _74517_ (_28888_, _28887_, _28886_);
  and _74518_ (_28889_, _28888_, _28885_);
  and _74519_ (_28890_, _28889_, _28882_);
  and _74520_ (_28891_, _28499_, _28463_);
  and _74521_ (_28892_, _28499_, _28470_);
  nor _74522_ (_28893_, _28892_, _28891_);
  and _74523_ (_28894_, _28544_, _28437_);
  and _74524_ (_28895_, _28499_, _28487_);
  nor _74525_ (_28896_, _28895_, _28894_);
  and _74526_ (_28897_, _28896_, _28893_);
  and _74527_ (_28898_, _28467_, _28446_);
  and _74528_ (_28899_, _28447_, _28431_);
  nor _74529_ (_28900_, _28899_, _28898_);
  and _74530_ (_28901_, _28509_, _28499_);
  and _74531_ (_28902_, _28490_, _28447_);
  nor _74532_ (_28903_, _28902_, _28901_);
  and _74533_ (_28904_, _28903_, _28900_);
  and _74534_ (_28905_, _28904_, _28897_);
  and _74535_ (_28906_, _28905_, _28890_);
  and _74536_ (_28907_, _28906_, _28875_);
  and _74537_ (_28908_, _28525_, _28487_);
  and _74538_ (_28909_, _28525_, _28476_);
  nor _74539_ (_28910_, _28909_, _28908_);
  and _74540_ (_28911_, _28525_, _28492_);
  and _74541_ (_28912_, _28554_, _28525_);
  nor _74542_ (_28913_, _28912_, _28911_);
  and _74543_ (_28914_, _28913_, _28910_);
  and _74544_ (_28915_, _28544_, _28463_);
  and _74545_ (_28916_, _28544_, _28431_);
  nor _74546_ (_28917_, _28916_, _28915_);
  and _74547_ (_28918_, _28525_, _28446_);
  and _74548_ (_28919_, _28549_, _28449_);
  nor _74549_ (_28920_, _28919_, _28918_);
  and _74550_ (_28921_, _28920_, _28917_);
  and _74551_ (_28922_, _28921_, _28914_);
  and _74552_ (_28923_, _28579_, _28422_);
  and _74553_ (_28924_, _28579_, _28434_);
  nor _74554_ (_28925_, _28924_, _28923_);
  and _74555_ (_28926_, _28538_, _28514_);
  and _74556_ (_28927_, _28579_, _28470_);
  nor _74557_ (_28928_, _28927_, _28926_);
  and _74558_ (_28929_, _28928_, _28925_);
  and _74559_ (_28930_, _28579_, _28487_);
  and _74560_ (_28931_, _28579_, _28492_);
  nor _74561_ (_28932_, _28931_, _28930_);
  and _74562_ (_28933_, _28579_, _28476_);
  and _74563_ (_28934_, _28579_, _28514_);
  nor _74564_ (_28935_, _28934_, _28933_);
  and _74565_ (_28936_, _28935_, _28932_);
  and _74566_ (_28937_, _28936_, _28929_);
  and _74567_ (_28938_, _28937_, _28922_);
  and _74568_ (_28939_, _28528_, _28479_);
  and _74569_ (_28940_, _28528_, _28509_);
  nor _74570_ (_28941_, _28940_, _28939_);
  and _74571_ (_28942_, _28476_, _28441_);
  and _74572_ (_28943_, _28528_, _28463_);
  nor _74573_ (_28944_, _28943_, _28942_);
  and _74574_ (_28945_, _28944_, _28941_);
  and _74575_ (_28946_, _28461_, _28449_);
  and _74576_ (_28947_, _28476_, _28461_);
  nor _74577_ (_28948_, _28947_, _28946_);
  and _74578_ (_28949_, _28549_, _28446_);
  and _74579_ (_28950_, _28509_, _28461_);
  nor _74580_ (_28951_, _28950_, _28949_);
  and _74581_ (_28952_, _28951_, _28948_);
  and _74582_ (_28953_, _28952_, _28945_);
  and _74583_ (_28954_, _28544_, _28492_);
  and _74584_ (_28955_, _28470_, _28441_);
  nor _74585_ (_28956_, _28955_, _28954_);
  and _74586_ (_28957_, _28554_, _28544_);
  and _74587_ (_28958_, _28446_, _28441_);
  nor _74588_ (_28959_, _28958_, _28957_);
  and _74589_ (_28960_, _28959_, _28956_);
  and _74590_ (_28961_, _28463_, _28452_);
  and _74591_ (_28962_, _28492_, _28441_);
  nor _74592_ (_28963_, _28962_, _28961_);
  and _74593_ (_28964_, _28514_, _28441_);
  and _74594_ (_28965_, _28554_, _28441_);
  nor _74595_ (_28966_, _28965_, _28964_);
  and _74596_ (_28967_, _28966_, _28963_);
  and _74597_ (_28968_, _28967_, _28960_);
  and _74598_ (_28969_, _28968_, _28953_);
  and _74599_ (_28970_, _28969_, _28938_);
  and _74600_ (_28971_, _28970_, _28907_);
  and _74601_ (_28972_, _28971_, _28844_);
  and _74602_ (_28973_, _28972_, _28725_);
  and _74603_ (_28974_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  not _74604_ (_28975_, _28974_);
  and _74605_ (_28976_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and _74606_ (_28977_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  nor _74607_ (_28978_, _28977_, _28976_);
  and _74608_ (_28979_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  and _74609_ (_28980_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  nor _74610_ (_28981_, _28980_, _28979_);
  and _74611_ (_28982_, _28981_, _28978_);
  and _74612_ (_28983_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and _74613_ (_28984_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  nor _74614_ (_28985_, _28984_, _28983_);
  and _74615_ (_28986_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  and _74616_ (_28987_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  nor _74617_ (_28988_, _28987_, _28986_);
  and _74618_ (_28989_, _28988_, _28985_);
  and _74619_ (_28990_, _28989_, _28982_);
  and _74620_ (_28991_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  and _74621_ (_28992_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  nor _74622_ (_28993_, _28992_, _28991_);
  and _74623_ (_28994_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and _74624_ (_28995_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  nor _74625_ (_28996_, _28995_, _28994_);
  and _74626_ (_28997_, _28996_, _28993_);
  and _74627_ (_28998_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  and _74628_ (_28999_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  nor _74629_ (_29000_, _28999_, _28998_);
  and _74630_ (_29001_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and _74631_ (_29002_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  nor _74632_ (_29003_, _29002_, _29001_);
  and _74633_ (_29004_, _29003_, _29000_);
  and _74634_ (_29005_, _29004_, _28997_);
  and _74635_ (_29006_, _29005_, _28990_);
  and _74636_ (_29007_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and _74637_ (_29008_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  nor _74638_ (_29009_, _29008_, _29007_);
  and _74639_ (_29010_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  and _74640_ (_29011_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  nor _74641_ (_29012_, _29011_, _29010_);
  and _74642_ (_29013_, _29012_, _29009_);
  and _74643_ (_29014_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  and _74644_ (_29015_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  nor _74645_ (_29016_, _29015_, _29014_);
  and _74646_ (_29017_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and _74647_ (_29018_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  nor _74648_ (_29019_, _29018_, _29017_);
  and _74649_ (_29020_, _29019_, _29016_);
  and _74650_ (_29021_, _29020_, _29013_);
  and _74651_ (_29022_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and _74652_ (_29023_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  nor _74653_ (_29024_, _29023_, _29022_);
  and _74654_ (_29025_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  and _74655_ (_29026_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  nor _74656_ (_29027_, _29026_, _29025_);
  and _74657_ (_29028_, _29027_, _29024_);
  and _74658_ (_29029_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and _74659_ (_29030_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  nor _74660_ (_29031_, _29030_, _29029_);
  and _74661_ (_29032_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  and _74662_ (_29033_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  nor _74663_ (_29034_, _29033_, _29032_);
  and _74664_ (_29035_, _29034_, _29031_);
  and _74665_ (_29036_, _29035_, _29028_);
  and _74666_ (_29037_, _29036_, _29021_);
  and _74667_ (_29038_, _29037_, _29006_);
  and _74668_ (_29039_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and _74669_ (_29040_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  nor _74670_ (_29041_, _29040_, _29039_);
  and _74671_ (_29042_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  and _74672_ (_29043_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  nor _74673_ (_29044_, _29043_, _29042_);
  and _74674_ (_29045_, _29044_, _29041_);
  and _74675_ (_29046_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and _74676_ (_29047_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  nor _74677_ (_29048_, _29047_, _29046_);
  and _74678_ (_29049_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  and _74679_ (_29050_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  nor _74680_ (_29051_, _29050_, _29049_);
  and _74681_ (_29052_, _29051_, _29048_);
  and _74682_ (_29053_, _29052_, _29045_);
  and _74683_ (_29054_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  and _74684_ (_29055_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  nor _74685_ (_29056_, _29055_, _29054_);
  and _74686_ (_29057_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and _74687_ (_29058_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  nor _74688_ (_29059_, _29058_, _29057_);
  and _74689_ (_29060_, _29059_, _29056_);
  and _74690_ (_29061_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  and _74691_ (_29062_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  nor _74692_ (_29063_, _29062_, _29061_);
  and _74693_ (_29064_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and _74694_ (_29065_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  nor _74695_ (_29066_, _29065_, _29064_);
  and _74696_ (_29067_, _29066_, _29063_);
  and _74697_ (_29068_, _29067_, _29060_);
  and _74698_ (_29069_, _29068_, _29053_);
  and _74699_ (_29070_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  and _74700_ (_29071_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  nor _74701_ (_29072_, _29071_, _29070_);
  and _74702_ (_29073_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  and _74703_ (_29074_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  nor _74704_ (_29075_, _29074_, _29073_);
  and _74705_ (_29076_, _29075_, _29072_);
  and _74706_ (_29077_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  and _74707_ (_29078_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  nor _74708_ (_29079_, _29078_, _29077_);
  and _74709_ (_29080_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and _74710_ (_29081_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  nor _74711_ (_29082_, _29081_, _29080_);
  and _74712_ (_29083_, _29082_, _29079_);
  and _74713_ (_29084_, _29083_, _29076_);
  and _74714_ (_29085_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and _74715_ (_29086_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  nor _74716_ (_29087_, _29086_, _29085_);
  and _74717_ (_29088_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  and _74718_ (_29089_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  nor _74719_ (_29090_, _29089_, _29088_);
  and _74720_ (_29091_, _29090_, _29087_);
  and _74721_ (_29092_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and _74722_ (_29093_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  nor _74723_ (_29094_, _29093_, _29092_);
  and _74724_ (_29095_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  and _74725_ (_29096_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  nor _74726_ (_29097_, _29096_, _29095_);
  and _74727_ (_29098_, _29097_, _29094_);
  and _74728_ (_29099_, _29098_, _29091_);
  and _74729_ (_29100_, _29099_, _29084_);
  and _74730_ (_29101_, _29100_, _29069_);
  and _74731_ (_29102_, _29101_, _29038_);
  and _74732_ (_29103_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  and _74733_ (_29104_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  nor _74734_ (_29105_, _29104_, _29103_);
  and _74735_ (_29106_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and _74736_ (_29107_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  nor _74737_ (_29108_, _29107_, _29106_);
  and _74738_ (_29109_, _29108_, _29105_);
  and _74739_ (_29110_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  and _74740_ (_29111_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  nor _74741_ (_29112_, _29111_, _29110_);
  and _74742_ (_29113_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and _74743_ (_29114_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  nor _74744_ (_29115_, _29114_, _29113_);
  and _74745_ (_29116_, _29115_, _29112_);
  and _74746_ (_29117_, _29116_, _29109_);
  and _74747_ (_29118_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and _74748_ (_29119_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  nor _74749_ (_29120_, _29119_, _29118_);
  and _74750_ (_29121_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  and _74751_ (_29122_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  nor _74752_ (_29123_, _29122_, _29121_);
  and _74753_ (_29124_, _29123_, _29120_);
  and _74754_ (_29125_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and _74755_ (_29126_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  nor _74756_ (_29127_, _29126_, _29125_);
  and _74757_ (_29128_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  and _74758_ (_29129_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  nor _74759_ (_29130_, _29129_, _29128_);
  and _74760_ (_29131_, _29130_, _29127_);
  and _74761_ (_29132_, _29131_, _29124_);
  and _74762_ (_29133_, _29132_, _29117_);
  and _74763_ (_29134_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  and _74764_ (_29135_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  nor _74765_ (_29136_, _29135_, _29134_);
  and _74766_ (_29137_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and _74767_ (_29138_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  nor _74768_ (_29139_, _29138_, _29137_);
  and _74769_ (_29140_, _29139_, _29136_);
  and _74770_ (_29141_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  and _74771_ (_29142_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  nor _74772_ (_29143_, _29142_, _29141_);
  and _74773_ (_29144_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  and _74774_ (_29145_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  nor _74775_ (_29146_, _29145_, _29144_);
  and _74776_ (_29147_, _29146_, _29143_);
  and _74777_ (_29148_, _29147_, _29140_);
  and _74778_ (_29149_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  and _74779_ (_29150_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  nor _74780_ (_29151_, _29150_, _29149_);
  and _74781_ (_29152_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and _74782_ (_29153_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  nor _74783_ (_29154_, _29153_, _29152_);
  and _74784_ (_29155_, _29154_, _29151_);
  and _74785_ (_29156_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and _74786_ (_29157_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  nor _74787_ (_29158_, _29157_, _29156_);
  and _74788_ (_29159_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  and _74789_ (_29160_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  nor _74790_ (_29161_, _29160_, _29159_);
  and _74791_ (_29162_, _29161_, _29158_);
  and _74792_ (_29163_, _29162_, _29155_);
  and _74793_ (_29164_, _29163_, _29148_);
  and _74794_ (_29165_, _29164_, _29133_);
  and _74795_ (_29166_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and _74796_ (_29167_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  nor _74797_ (_29168_, _29167_, _29166_);
  and _74798_ (_29169_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  and _74799_ (_29170_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  nor _74800_ (_29171_, _29170_, _29169_);
  and _74801_ (_29172_, _29171_, _29168_);
  and _74802_ (_29173_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and _74803_ (_29174_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  nor _74804_ (_29175_, _29174_, _29173_);
  and _74805_ (_29176_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  and _74806_ (_29177_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  nor _74807_ (_29178_, _29177_, _29176_);
  and _74808_ (_29179_, _29178_, _29175_);
  and _74809_ (_29180_, _29179_, _29172_);
  and _74810_ (_29181_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  and _74811_ (_29182_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  nor _74812_ (_29183_, _29182_, _29181_);
  and _74813_ (_29184_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  and _74814_ (_29185_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  nor _74815_ (_29186_, _29185_, _29184_);
  and _74816_ (_29187_, _29186_, _29183_);
  and _74817_ (_29188_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  and _74818_ (_29189_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  nor _74819_ (_29190_, _29189_, _29188_);
  and _74820_ (_29191_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and _74821_ (_29192_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  nor _74822_ (_29193_, _29192_, _29191_);
  and _74823_ (_29194_, _29193_, _29190_);
  and _74824_ (_29195_, _29194_, _29187_);
  and _74825_ (_29196_, _29195_, _29180_);
  and _74826_ (_29197_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and _74827_ (_29198_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  nor _74828_ (_29199_, _29198_, _29197_);
  and _74829_ (_29200_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  and _74830_ (_29201_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  nor _74831_ (_29202_, _29201_, _29200_);
  and _74832_ (_29203_, _29202_, _29199_);
  and _74833_ (_29204_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and _74834_ (_29205_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  nor _74835_ (_29206_, _29205_, _29204_);
  and _74836_ (_29207_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and _74837_ (_29208_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  nor _74838_ (_29209_, _29208_, _29207_);
  and _74839_ (_29210_, _29209_, _29206_);
  and _74840_ (_29211_, _29210_, _29203_);
  and _74841_ (_29212_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  and _74842_ (_29213_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  nor _74843_ (_29214_, _29213_, _29212_);
  and _74844_ (_29215_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and _74845_ (_29216_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  nor _74846_ (_29217_, _29216_, _29215_);
  and _74847_ (_29218_, _29217_, _29214_);
  and _74848_ (_29219_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  and _74849_ (_29220_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  nor _74850_ (_29221_, _29220_, _29219_);
  and _74851_ (_29222_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and _74852_ (_29223_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  nor _74853_ (_29224_, _29223_, _29222_);
  and _74854_ (_29225_, _29224_, _29221_);
  and _74855_ (_29226_, _29225_, _29218_);
  and _74856_ (_29227_, _29226_, _29211_);
  and _74857_ (_29228_, _29227_, _29196_);
  and _74858_ (_29229_, _29228_, _29165_);
  and _74859_ (_29230_, _29229_, _29102_);
  and _74860_ (_29231_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  and _74861_ (_29232_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  nor _74862_ (_29233_, _29232_, _29231_);
  and _74863_ (_29234_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and _74864_ (_29235_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  nor _74865_ (_29236_, _29235_, _29234_);
  and _74866_ (_29237_, _29236_, _29233_);
  and _74867_ (_29238_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  and _74868_ (_29239_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  nor _74869_ (_29240_, _29239_, _29238_);
  and _74870_ (_29241_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and _74871_ (_29242_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  nor _74872_ (_29243_, _29242_, _29241_);
  and _74873_ (_29244_, _29243_, _29240_);
  and _74874_ (_29245_, _29244_, _29237_);
  and _74875_ (_29246_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and _74876_ (_29247_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  nor _74877_ (_29248_, _29247_, _29246_);
  and _74878_ (_29249_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  and _74879_ (_29250_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  nor _74880_ (_29251_, _29250_, _29249_);
  and _74881_ (_29252_, _29251_, _29248_);
  and _74882_ (_29253_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and _74883_ (_29254_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  nor _74884_ (_29255_, _29254_, _29253_);
  and _74885_ (_29256_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  and _74886_ (_29257_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  nor _74887_ (_29258_, _29257_, _29256_);
  and _74888_ (_29259_, _29258_, _29255_);
  and _74889_ (_29260_, _29259_, _29252_);
  and _74890_ (_29261_, _29260_, _29245_);
  and _74891_ (_29262_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and _74892_ (_29263_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  nor _74893_ (_29264_, _29263_, _29262_);
  and _74894_ (_29265_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  and _74895_ (_29266_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  nor _74896_ (_29267_, _29266_, _29265_);
  and _74897_ (_29268_, _29267_, _29264_);
  and _74898_ (_29269_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and _74899_ (_29270_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  nor _74900_ (_29271_, _29270_, _29269_);
  and _74901_ (_29272_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  and _74902_ (_29273_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  nor _74903_ (_29274_, _29273_, _29272_);
  and _74904_ (_29275_, _29274_, _29271_);
  and _74905_ (_29276_, _29275_, _29268_);
  and _74906_ (_29277_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  and _74907_ (_29278_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  nor _74908_ (_29279_, _29278_, _29277_);
  and _74909_ (_29280_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and _74910_ (_29281_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  nor _74911_ (_29282_, _29281_, _29280_);
  and _74912_ (_29283_, _29282_, _29279_);
  and _74913_ (_29284_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and _74914_ (_29285_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  nor _74915_ (_29286_, _29285_, _29284_);
  and _74916_ (_29287_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  and _74917_ (_29288_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  nor _74918_ (_29289_, _29288_, _29287_);
  and _74919_ (_29290_, _29289_, _29286_);
  and _74920_ (_29291_, _29290_, _29283_);
  and _74921_ (_29292_, _29291_, _29276_);
  and _74922_ (_29293_, _29292_, _29261_);
  and _74923_ (_29294_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  and _74924_ (_29295_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  nor _74925_ (_29296_, _29295_, _29294_);
  and _74926_ (_29297_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and _74927_ (_29298_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  nor _74928_ (_29299_, _29298_, _29297_);
  and _74929_ (_29300_, _29299_, _29296_);
  and _74930_ (_29301_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  and _74931_ (_29302_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  nor _74932_ (_29303_, _29302_, _29301_);
  and _74933_ (_29304_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and _74934_ (_29305_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  nor _74935_ (_29306_, _29305_, _29304_);
  and _74936_ (_29307_, _29306_, _29303_);
  and _74937_ (_29308_, _29307_, _29300_);
  and _74938_ (_29309_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  and _74939_ (_29310_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  nor _74940_ (_29311_, _29310_, _29309_);
  and _74941_ (_29312_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and _74942_ (_29313_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  nor _74943_ (_29314_, _29313_, _29312_);
  and _74944_ (_29315_, _29314_, _29311_);
  and _74945_ (_29316_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and _74946_ (_29317_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  nor _74947_ (_29318_, _29317_, _29316_);
  and _74948_ (_29319_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  and _74949_ (_29320_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  nor _74950_ (_29321_, _29320_, _29319_);
  and _74951_ (_29322_, _29321_, _29318_);
  and _74952_ (_29323_, _29322_, _29315_);
  and _74953_ (_29324_, _29323_, _29308_);
  and _74954_ (_29325_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and _74955_ (_29326_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  nor _74956_ (_29327_, _29326_, _29325_);
  and _74957_ (_29328_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  and _74958_ (_29329_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  nor _74959_ (_29330_, _29329_, _29328_);
  and _74960_ (_29331_, _29330_, _29327_);
  and _74961_ (_29332_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and _74962_ (_29333_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  nor _74963_ (_29334_, _29333_, _29332_);
  and _74964_ (_29335_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and _74965_ (_29336_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  nor _74966_ (_29337_, _29336_, _29335_);
  and _74967_ (_29338_, _29337_, _29334_);
  and _74968_ (_29339_, _29338_, _29331_);
  and _74969_ (_29340_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  and _74970_ (_29341_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  nor _74971_ (_29342_, _29341_, _29340_);
  and _74972_ (_29343_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and _74973_ (_29344_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  nor _74974_ (_29345_, _29344_, _29343_);
  and _74975_ (_29346_, _29345_, _29342_);
  and _74976_ (_29347_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  and _74977_ (_29348_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  nor _74978_ (_29349_, _29348_, _29347_);
  and _74979_ (_29350_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  and _74980_ (_29351_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  nor _74981_ (_29352_, _29351_, _29350_);
  and _74982_ (_29353_, _29352_, _29349_);
  and _74983_ (_29354_, _29353_, _29346_);
  and _74984_ (_29355_, _29354_, _29339_);
  and _74985_ (_29356_, _29355_, _29324_);
  and _74986_ (_29357_, _29356_, _29293_);
  and _74987_ (_29358_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  and _74988_ (_29359_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  nor _74989_ (_29360_, _29359_, _29358_);
  and _74990_ (_29361_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and _74991_ (_29362_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  nor _74992_ (_29363_, _29362_, _29361_);
  and _74993_ (_29364_, _29363_, _29360_);
  and _74994_ (_29365_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  and _74995_ (_29366_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  nor _74996_ (_29367_, _29366_, _29365_);
  and _74997_ (_29368_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and _74998_ (_29369_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  nor _74999_ (_29370_, _29369_, _29368_);
  and _75000_ (_29371_, _29370_, _29367_);
  and _75001_ (_29372_, _29371_, _29364_);
  and _75002_ (_29373_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and _75003_ (_29374_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  nor _75004_ (_29375_, _29374_, _29373_);
  and _75005_ (_29376_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and _75006_ (_29377_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  nor _75007_ (_29378_, _29377_, _29376_);
  and _75008_ (_29379_, _29378_, _29375_);
  and _75009_ (_29380_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and _75010_ (_29381_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  nor _75011_ (_29382_, _29381_, _29380_);
  and _75012_ (_29383_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  and _75013_ (_29384_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  nor _75014_ (_29385_, _29384_, _29383_);
  and _75015_ (_29386_, _29385_, _29382_);
  and _75016_ (_29387_, _29386_, _29379_);
  and _75017_ (_29388_, _29387_, _29372_);
  and _75018_ (_29389_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and _75019_ (_29390_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  nor _75020_ (_29391_, _29390_, _29389_);
  and _75021_ (_29392_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  and _75022_ (_29393_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  nor _75023_ (_29394_, _29393_, _29392_);
  and _75024_ (_29395_, _29394_, _29391_);
  and _75025_ (_29396_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and _75026_ (_29397_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  nor _75027_ (_29398_, _29397_, _29396_);
  and _75028_ (_29399_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  and _75029_ (_29400_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  nor _75030_ (_29401_, _29400_, _29399_);
  and _75031_ (_29402_, _29401_, _29398_);
  and _75032_ (_29403_, _29402_, _29395_);
  and _75033_ (_29404_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  and _75034_ (_29405_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  nor _75035_ (_29406_, _29405_, _29404_);
  and _75036_ (_29407_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  and _75037_ (_29408_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  nor _75038_ (_29409_, _29408_, _29407_);
  and _75039_ (_29410_, _29409_, _29406_);
  and _75040_ (_29411_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  and _75041_ (_29412_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  nor _75042_ (_29413_, _29412_, _29411_);
  and _75043_ (_29414_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and _75044_ (_29415_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  nor _75045_ (_29416_, _29415_, _29414_);
  and _75046_ (_29417_, _29416_, _29413_);
  and _75047_ (_29418_, _29417_, _29410_);
  and _75048_ (_29419_, _29418_, _29403_);
  and _75049_ (_29420_, _29419_, _29388_);
  and _75050_ (_29421_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  and _75051_ (_29422_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  nor _75052_ (_29423_, _29422_, _29421_);
  and _75053_ (_29424_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and _75054_ (_29425_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  nor _75055_ (_29426_, _29425_, _29424_);
  and _75056_ (_29427_, _29426_, _29423_);
  and _75057_ (_29428_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  and _75058_ (_29429_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  nor _75059_ (_29430_, _29429_, _29428_);
  and _75060_ (_29431_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and _75061_ (_29432_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  nor _75062_ (_29433_, _29432_, _29431_);
  and _75063_ (_29434_, _29433_, _29430_);
  and _75064_ (_29435_, _29434_, _29427_);
  and _75065_ (_29436_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and _75066_ (_29437_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  nor _75067_ (_29438_, _29437_, _29436_);
  and _75068_ (_29439_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  and _75069_ (_29440_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  nor _75070_ (_29441_, _29440_, _29439_);
  and _75071_ (_29442_, _29441_, _29438_);
  and _75072_ (_29443_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and _75073_ (_29444_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  nor _75074_ (_29445_, _29444_, _29443_);
  and _75075_ (_29446_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and _75076_ (_29447_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  nor _75077_ (_29448_, _29447_, _29446_);
  and _75078_ (_29449_, _29448_, _29445_);
  and _75079_ (_29450_, _29449_, _29442_);
  and _75080_ (_29451_, _29450_, _29435_);
  and _75081_ (_29452_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and _75082_ (_29453_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor _75083_ (_29454_, _29453_, _29452_);
  and _75084_ (_29455_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and _75085_ (_29456_, _28538_, _28479_);
  and _75086_ (_29457_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor _75087_ (_29458_, _29457_, _29455_);
  and _75088_ (_29459_, _29458_, _29454_);
  and _75089_ (_29460_, _28538_, _28490_);
  and _75090_ (_29461_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and _75091_ (_29462_, _28538_, _28449_);
  and _75092_ (_29463_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and _75093_ (_29464_, _28538_, _28437_);
  and _75094_ (_29465_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or _75095_ (_29466_, _29465_, _29463_);
  nor _75096_ (_29467_, _29466_, _29461_);
  and _75097_ (_29468_, _29467_, _29459_);
  and _75098_ (_29469_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and _75099_ (_29470_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor _75100_ (_29471_, _29470_, _29469_);
  and _75101_ (_29472_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and _75102_ (_29473_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor _75103_ (_29474_, _29473_, _29472_);
  and _75104_ (_29475_, _29474_, _29471_);
  and _75105_ (_29476_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and _75106_ (_29477_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor _75107_ (_29478_, _29477_, _29476_);
  and _75108_ (_29479_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and _75109_ (_29480_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor _75110_ (_29481_, _29480_, _29479_);
  and _75111_ (_29482_, _29481_, _29478_);
  and _75112_ (_29483_, _29482_, _29475_);
  and _75113_ (_29484_, _29483_, _29468_);
  and _75114_ (_29485_, _29484_, _29451_);
  and _75115_ (_29486_, _29485_, _29420_);
  and _75116_ (_29487_, _29486_, _29357_);
  and _75117_ (_29488_, _29487_, _29230_);
  and _75118_ (_29489_, _29488_, _28975_);
  and _75119_ (_29490_, iram_op1_reg[0], iram_op1_reg[1]);
  and _75120_ (_29491_, _29490_, iram_op1_reg[2]);
  nor _75121_ (_29492_, _29490_, iram_op1_reg[2]);
  nor _75122_ (_29493_, _29492_, _29491_);
  nor _75123_ (_29494_, _29493_, _29489_);
  and _75124_ (_29495_, _29493_, _29489_);
  or _75125_ (_29496_, _29495_, _29494_);
  and _75126_ (_29497_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  not _75127_ (_29498_, _29497_);
  and _75128_ (_29499_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  and _75129_ (_29500_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  nor _75130_ (_29501_, _29500_, _29499_);
  and _75131_ (_29502_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and _75132_ (_29503_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  nor _75133_ (_29504_, _29503_, _29502_);
  and _75134_ (_29505_, _29504_, _29501_);
  and _75135_ (_29506_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and _75136_ (_29507_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  nor _75137_ (_29508_, _29507_, _29506_);
  and _75138_ (_29509_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and _75139_ (_29510_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  nor _75140_ (_29511_, _29510_, _29509_);
  and _75141_ (_29512_, _29511_, _29508_);
  and _75142_ (_29513_, _29512_, _29505_);
  and _75143_ (_29514_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and _75144_ (_29515_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  nor _75145_ (_29516_, _29515_, _29514_);
  and _75146_ (_29517_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  and _75147_ (_29518_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  nor _75148_ (_29519_, _29518_, _29517_);
  and _75149_ (_29520_, _29519_, _29516_);
  and _75150_ (_29521_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  and _75151_ (_29522_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  nor _75152_ (_29523_, _29522_, _29521_);
  and _75153_ (_29524_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and _75154_ (_29525_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  nor _75155_ (_29526_, _29525_, _29524_);
  and _75156_ (_29527_, _29526_, _29523_);
  and _75157_ (_29528_, _29527_, _29520_);
  and _75158_ (_29529_, _29528_, _29513_);
  and _75159_ (_29530_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and _75160_ (_29531_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  nor _75161_ (_29532_, _29531_, _29530_);
  and _75162_ (_29533_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  and _75163_ (_29534_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  nor _75164_ (_29535_, _29534_, _29533_);
  and _75165_ (_29536_, _29535_, _29532_);
  and _75166_ (_29537_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and _75167_ (_29538_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  nor _75168_ (_29539_, _29538_, _29537_);
  and _75169_ (_29540_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  and _75170_ (_29541_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  nor _75171_ (_29542_, _29541_, _29540_);
  and _75172_ (_29543_, _29542_, _29539_);
  and _75173_ (_29544_, _29543_, _29536_);
  and _75174_ (_29545_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  and _75175_ (_29546_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  nor _75176_ (_29547_, _29546_, _29545_);
  and _75177_ (_29548_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  and _75178_ (_29549_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  nor _75179_ (_29550_, _29549_, _29548_);
  and _75180_ (_29551_, _29550_, _29547_);
  and _75181_ (_29552_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  and _75182_ (_29553_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  nor _75183_ (_29554_, _29553_, _29552_);
  and _75184_ (_29555_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and _75185_ (_29556_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  nor _75186_ (_29557_, _29556_, _29555_);
  and _75187_ (_29558_, _29557_, _29554_);
  and _75188_ (_29559_, _29558_, _29551_);
  and _75189_ (_29560_, _29559_, _29544_);
  and _75190_ (_29561_, _29560_, _29529_);
  and _75191_ (_29562_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and _75192_ (_29563_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  nor _75193_ (_29564_, _29563_, _29562_);
  and _75194_ (_29565_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  and _75195_ (_29566_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  nor _75196_ (_29567_, _29566_, _29565_);
  and _75197_ (_29568_, _29567_, _29564_);
  and _75198_ (_29569_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and _75199_ (_29570_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  nor _75200_ (_29571_, _29570_, _29569_);
  and _75201_ (_29572_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and _75202_ (_29573_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  nor _75203_ (_29574_, _29573_, _29572_);
  and _75204_ (_29575_, _29574_, _29571_);
  and _75205_ (_29576_, _29575_, _29568_);
  and _75206_ (_29577_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  and _75207_ (_29578_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  nor _75208_ (_29579_, _29578_, _29577_);
  and _75209_ (_29580_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and _75210_ (_29581_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  nor _75211_ (_29582_, _29581_, _29580_);
  and _75212_ (_29583_, _29582_, _29579_);
  and _75213_ (_29584_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  and _75214_ (_29585_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  nor _75215_ (_29586_, _29585_, _29584_);
  and _75216_ (_29587_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and _75217_ (_29588_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  nor _75218_ (_29589_, _29588_, _29587_);
  and _75219_ (_29590_, _29589_, _29586_);
  and _75220_ (_29591_, _29590_, _29583_);
  and _75221_ (_29592_, _29591_, _29576_);
  and _75222_ (_29593_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  and _75223_ (_29594_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  nor _75224_ (_29595_, _29594_, _29593_);
  and _75225_ (_29596_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and _75226_ (_29597_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  nor _75227_ (_29598_, _29597_, _29596_);
  and _75228_ (_29599_, _29598_, _29595_);
  and _75229_ (_29600_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  and _75230_ (_29601_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  nor _75231_ (_29602_, _29601_, _29600_);
  and _75232_ (_29603_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  and _75233_ (_29604_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  nor _75234_ (_29605_, _29604_, _29603_);
  and _75235_ (_29606_, _29605_, _29602_);
  and _75236_ (_29607_, _29606_, _29599_);
  and _75237_ (_29608_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and _75238_ (_29609_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  nor _75239_ (_29610_, _29609_, _29608_);
  and _75240_ (_29611_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  and _75241_ (_29612_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  nor _75242_ (_29613_, _29612_, _29611_);
  and _75243_ (_29614_, _29613_, _29610_);
  and _75244_ (_29615_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and _75245_ (_29616_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  nor _75246_ (_29617_, _29616_, _29615_);
  and _75247_ (_29618_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  and _75248_ (_29619_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  nor _75249_ (_29620_, _29619_, _29618_);
  and _75250_ (_29621_, _29620_, _29617_);
  and _75251_ (_29622_, _29621_, _29614_);
  and _75252_ (_29623_, _29622_, _29607_);
  and _75253_ (_29624_, _29623_, _29592_);
  and _75254_ (_29625_, _29624_, _29561_);
  and _75255_ (_29626_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  and _75256_ (_29627_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  nor _75257_ (_29628_, _29627_, _29626_);
  and _75258_ (_29629_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and _75259_ (_29630_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  nor _75260_ (_29631_, _29630_, _29629_);
  and _75261_ (_29632_, _29631_, _29628_);
  and _75262_ (_29633_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  and _75263_ (_29634_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  nor _75264_ (_29635_, _29634_, _29633_);
  and _75265_ (_29636_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  and _75266_ (_29637_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  nor _75267_ (_29638_, _29637_, _29636_);
  and _75268_ (_29639_, _29638_, _29635_);
  and _75269_ (_29640_, _29639_, _29632_);
  and _75270_ (_29641_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and _75271_ (_29642_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  nor _75272_ (_29643_, _29642_, _29641_);
  and _75273_ (_29644_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  and _75274_ (_29645_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  nor _75275_ (_29646_, _29645_, _29644_);
  and _75276_ (_29647_, _29646_, _29643_);
  and _75277_ (_29648_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and _75278_ (_29649_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  nor _75279_ (_29650_, _29649_, _29648_);
  and _75280_ (_29651_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  and _75281_ (_29652_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  nor _75282_ (_29653_, _29652_, _29651_);
  and _75283_ (_29654_, _29653_, _29650_);
  and _75284_ (_29655_, _29654_, _29647_);
  and _75285_ (_29656_, _29655_, _29640_);
  and _75286_ (_29657_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  and _75287_ (_29658_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  nor _75288_ (_29659_, _29658_, _29657_);
  and _75289_ (_29660_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and _75290_ (_29661_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  nor _75291_ (_29662_, _29661_, _29660_);
  and _75292_ (_29663_, _29662_, _29659_);
  and _75293_ (_29664_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and _75294_ (_29665_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  nor _75295_ (_29666_, _29665_, _29664_);
  and _75296_ (_29667_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and _75297_ (_29668_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  nor _75298_ (_29669_, _29668_, _29667_);
  and _75299_ (_29670_, _29669_, _29666_);
  and _75300_ (_29671_, _29670_, _29663_);
  and _75301_ (_29672_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  and _75302_ (_29673_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  nor _75303_ (_29674_, _29673_, _29672_);
  and _75304_ (_29675_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and _75305_ (_29676_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  nor _75306_ (_29677_, _29676_, _29675_);
  and _75307_ (_29678_, _29677_, _29674_);
  and _75308_ (_29679_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and _75309_ (_29680_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  nor _75310_ (_29681_, _29680_, _29679_);
  and _75311_ (_29682_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  and _75312_ (_29683_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  nor _75313_ (_29684_, _29683_, _29682_);
  and _75314_ (_29685_, _29684_, _29681_);
  and _75315_ (_29686_, _29685_, _29678_);
  and _75316_ (_29687_, _29686_, _29671_);
  and _75317_ (_29688_, _29687_, _29656_);
  and _75318_ (_29689_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and _75319_ (_29690_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  nor _75320_ (_29691_, _29690_, _29689_);
  and _75321_ (_29692_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  and _75322_ (_29693_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  nor _75323_ (_29694_, _29693_, _29692_);
  and _75324_ (_29695_, _29694_, _29691_);
  and _75325_ (_29696_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and _75326_ (_29697_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  nor _75327_ (_29698_, _29697_, _29696_);
  and _75328_ (_29699_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  and _75329_ (_29700_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  nor _75330_ (_29701_, _29700_, _29699_);
  and _75331_ (_29702_, _29701_, _29698_);
  and _75332_ (_29703_, _29702_, _29695_);
  and _75333_ (_29704_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  and _75334_ (_29705_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  nor _75335_ (_29706_, _29705_, _29704_);
  and _75336_ (_29707_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and _75337_ (_29708_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  nor _75338_ (_29709_, _29708_, _29707_);
  and _75339_ (_29710_, _29709_, _29706_);
  and _75340_ (_29711_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  and _75341_ (_29712_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  nor _75342_ (_29713_, _29712_, _29711_);
  and _75343_ (_29714_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and _75344_ (_29715_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  nor _75345_ (_29716_, _29715_, _29714_);
  and _75346_ (_29717_, _29716_, _29713_);
  and _75347_ (_29718_, _29717_, _29710_);
  and _75348_ (_29719_, _29718_, _29703_);
  and _75349_ (_29720_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  and _75350_ (_29721_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  nor _75351_ (_29722_, _29721_, _29720_);
  and _75352_ (_29723_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and _75353_ (_29724_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  nor _75354_ (_29725_, _29724_, _29723_);
  and _75355_ (_29726_, _29725_, _29722_);
  and _75356_ (_29727_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and _75357_ (_29728_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  nor _75358_ (_29729_, _29728_, _29727_);
  and _75359_ (_29730_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  and _75360_ (_29731_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  nor _75361_ (_29732_, _29731_, _29730_);
  and _75362_ (_29733_, _29732_, _29729_);
  and _75363_ (_29734_, _29733_, _29726_);
  and _75364_ (_29735_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  and _75365_ (_29736_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  nor _75366_ (_29737_, _29736_, _29735_);
  and _75367_ (_29738_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  and _75368_ (_29739_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  nor _75369_ (_29740_, _29739_, _29738_);
  and _75370_ (_29741_, _29740_, _29737_);
  and _75371_ (_29742_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  and _75372_ (_29743_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  nor _75373_ (_29744_, _29743_, _29742_);
  and _75374_ (_29745_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and _75375_ (_29746_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  nor _75376_ (_29747_, _29746_, _29745_);
  and _75377_ (_29748_, _29747_, _29744_);
  and _75378_ (_29749_, _29748_, _29741_);
  and _75379_ (_29750_, _29749_, _29734_);
  and _75380_ (_29751_, _29750_, _29719_);
  and _75381_ (_29752_, _29751_, _29688_);
  and _75382_ (_29753_, _29752_, _29625_);
  and _75383_ (_29754_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  and _75384_ (_29755_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  nor _75385_ (_29756_, _29755_, _29754_);
  and _75386_ (_29757_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and _75387_ (_29758_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  nor _75388_ (_29759_, _29758_, _29757_);
  and _75389_ (_29760_, _29759_, _29756_);
  and _75390_ (_29761_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  and _75391_ (_29762_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  nor _75392_ (_29763_, _29762_, _29761_);
  and _75393_ (_29764_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and _75394_ (_29765_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  nor _75395_ (_29766_, _29765_, _29764_);
  and _75396_ (_29767_, _29766_, _29763_);
  and _75397_ (_29768_, _29767_, _29760_);
  and _75398_ (_29769_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and _75399_ (_29770_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  nor _75400_ (_29771_, _29770_, _29769_);
  and _75401_ (_29772_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  and _75402_ (_29773_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  nor _75403_ (_29774_, _29773_, _29772_);
  and _75404_ (_29775_, _29774_, _29771_);
  and _75405_ (_29776_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and _75406_ (_29777_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  nor _75407_ (_29778_, _29777_, _29776_);
  and _75408_ (_29779_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  and _75409_ (_29780_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  nor _75410_ (_29781_, _29780_, _29779_);
  and _75411_ (_29782_, _29781_, _29778_);
  and _75412_ (_29783_, _29782_, _29775_);
  and _75413_ (_29784_, _29783_, _29768_);
  and _75414_ (_29785_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  and _75415_ (_29786_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  nor _75416_ (_29787_, _29786_, _29785_);
  and _75417_ (_29788_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and _75418_ (_29789_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  nor _75419_ (_29790_, _29789_, _29788_);
  and _75420_ (_29791_, _29790_, _29787_);
  and _75421_ (_29792_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and _75422_ (_29793_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  nor _75423_ (_29794_, _29793_, _29792_);
  and _75424_ (_29795_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and _75425_ (_29796_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  nor _75426_ (_29797_, _29796_, _29795_);
  and _75427_ (_29798_, _29797_, _29794_);
  and _75428_ (_29799_, _29798_, _29791_);
  and _75429_ (_29800_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  and _75430_ (_29801_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  nor _75431_ (_29802_, _29801_, _29800_);
  and _75432_ (_29803_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and _75433_ (_29804_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  nor _75434_ (_29805_, _29804_, _29803_);
  and _75435_ (_29806_, _29805_, _29802_);
  and _75436_ (_29807_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  and _75437_ (_29808_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  nor _75438_ (_29809_, _29808_, _29807_);
  and _75439_ (_29810_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and _75440_ (_29811_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  nor _75441_ (_29812_, _29811_, _29810_);
  and _75442_ (_29813_, _29812_, _29809_);
  and _75443_ (_29814_, _29813_, _29806_);
  and _75444_ (_29815_, _29814_, _29799_);
  and _75445_ (_29816_, _29815_, _29784_);
  and _75446_ (_29817_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and _75447_ (_29818_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  nor _75448_ (_29819_, _29818_, _29817_);
  and _75449_ (_29820_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  and _75450_ (_29821_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  nor _75451_ (_29822_, _29821_, _29820_);
  and _75452_ (_29823_, _29822_, _29819_);
  and _75453_ (_29824_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and _75454_ (_29825_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  nor _75455_ (_29826_, _29825_, _29824_);
  and _75456_ (_29827_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and _75457_ (_29828_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  nor _75458_ (_29829_, _29828_, _29827_);
  and _75459_ (_29830_, _29829_, _29826_);
  and _75460_ (_29831_, _29830_, _29823_);
  and _75461_ (_29832_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  and _75462_ (_29833_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  nor _75463_ (_29834_, _29833_, _29832_);
  and _75464_ (_29835_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and _75465_ (_29836_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  nor _75466_ (_29837_, _29836_, _29835_);
  and _75467_ (_29838_, _29837_, _29834_);
  and _75468_ (_29839_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  and _75469_ (_29840_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  nor _75470_ (_29841_, _29840_, _29839_);
  and _75471_ (_29842_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and _75472_ (_29843_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  nor _75473_ (_29844_, _29843_, _29842_);
  and _75474_ (_29845_, _29844_, _29841_);
  and _75475_ (_29846_, _29845_, _29838_);
  and _75476_ (_29847_, _29846_, _29831_);
  and _75477_ (_29848_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  and _75478_ (_29849_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  nor _75479_ (_29850_, _29849_, _29848_);
  and _75480_ (_29851_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and _75481_ (_29852_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  nor _75482_ (_29853_, _29852_, _29851_);
  and _75483_ (_29854_, _29853_, _29850_);
  and _75484_ (_29855_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  and _75485_ (_29856_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  nor _75486_ (_29857_, _29856_, _29855_);
  and _75487_ (_29858_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  and _75488_ (_29859_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  nor _75489_ (_29860_, _29859_, _29858_);
  and _75490_ (_29861_, _29860_, _29857_);
  and _75491_ (_29862_, _29861_, _29854_);
  and _75492_ (_29863_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and _75493_ (_29864_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  nor _75494_ (_29865_, _29864_, _29863_);
  and _75495_ (_29866_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  and _75496_ (_29867_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  nor _75497_ (_29868_, _29867_, _29866_);
  and _75498_ (_29869_, _29868_, _29865_);
  and _75499_ (_29870_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and _75500_ (_29871_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  nor _75501_ (_29872_, _29871_, _29870_);
  and _75502_ (_29873_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  and _75503_ (_29874_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  nor _75504_ (_29875_, _29874_, _29873_);
  and _75505_ (_29876_, _29875_, _29872_);
  and _75506_ (_29877_, _29876_, _29869_);
  and _75507_ (_29878_, _29877_, _29862_);
  and _75508_ (_29879_, _29878_, _29847_);
  and _75509_ (_29880_, _29879_, _29816_);
  and _75510_ (_29881_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and _75511_ (_29882_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  nor _75512_ (_29883_, _29882_, _29881_);
  and _75513_ (_29884_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  and _75514_ (_29885_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  nor _75515_ (_29886_, _29885_, _29884_);
  and _75516_ (_29887_, _29886_, _29883_);
  and _75517_ (_29888_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and _75518_ (_29889_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  nor _75519_ (_29890_, _29889_, _29888_);
  and _75520_ (_29891_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  and _75521_ (_29892_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  nor _75522_ (_29893_, _29892_, _29891_);
  and _75523_ (_29894_, _29893_, _29890_);
  and _75524_ (_29895_, _29894_, _29887_);
  and _75525_ (_29896_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  and _75526_ (_29897_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  nor _75527_ (_29898_, _29897_, _29896_);
  and _75528_ (_29899_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and _75529_ (_29900_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  nor _75530_ (_29901_, _29900_, _29899_);
  and _75531_ (_29902_, _29901_, _29898_);
  and _75532_ (_29903_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  and _75533_ (_29904_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  nor _75534_ (_29905_, _29904_, _29903_);
  and _75535_ (_29906_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and _75536_ (_29907_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  nor _75537_ (_29908_, _29907_, _29906_);
  and _75538_ (_29909_, _29908_, _29905_);
  and _75539_ (_29910_, _29909_, _29902_);
  and _75540_ (_29911_, _29910_, _29895_);
  and _75541_ (_29912_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and _75542_ (_29913_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  nor _75543_ (_29914_, _29913_, _29912_);
  and _75544_ (_29915_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  and _75545_ (_29916_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  nor _75546_ (_29917_, _29916_, _29915_);
  and _75547_ (_29918_, _29917_, _29914_);
  and _75548_ (_29919_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and _75549_ (_29920_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  nor _75550_ (_29921_, _29920_, _29919_);
  and _75551_ (_29922_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  and _75552_ (_29923_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  nor _75553_ (_29924_, _29923_, _29922_);
  and _75554_ (_29925_, _29924_, _29921_);
  and _75555_ (_29926_, _29925_, _29918_);
  and _75556_ (_29927_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  and _75557_ (_29928_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  nor _75558_ (_29929_, _29928_, _29927_);
  and _75559_ (_29930_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  and _75560_ (_29931_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  nor _75561_ (_29932_, _29931_, _29930_);
  and _75562_ (_29933_, _29932_, _29929_);
  and _75563_ (_29934_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  and _75564_ (_29935_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  nor _75565_ (_29936_, _29935_, _29934_);
  and _75566_ (_29937_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and _75567_ (_29938_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  nor _75568_ (_29939_, _29938_, _29937_);
  and _75569_ (_29940_, _29939_, _29936_);
  and _75570_ (_29941_, _29940_, _29933_);
  and _75571_ (_29942_, _29941_, _29926_);
  and _75572_ (_29943_, _29942_, _29911_);
  and _75573_ (_29944_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and _75574_ (_29945_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  nor _75575_ (_29946_, _29945_, _29944_);
  and _75576_ (_29947_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  and _75577_ (_29948_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  nor _75578_ (_29949_, _29948_, _29947_);
  and _75579_ (_29950_, _29949_, _29946_);
  and _75580_ (_29951_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and _75581_ (_29952_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  nor _75582_ (_29953_, _29952_, _29951_);
  and _75583_ (_29954_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  and _75584_ (_29955_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  nor _75585_ (_29956_, _29955_, _29954_);
  and _75586_ (_29957_, _29956_, _29953_);
  and _75587_ (_29958_, _29957_, _29950_);
  and _75588_ (_29959_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  and _75589_ (_29960_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  nor _75590_ (_29961_, _29960_, _29959_);
  and _75591_ (_29962_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and _75592_ (_29963_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  nor _75593_ (_29964_, _29963_, _29962_);
  and _75594_ (_29965_, _29964_, _29961_);
  and _75595_ (_29966_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  and _75596_ (_29967_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  nor _75597_ (_29968_, _29967_, _29966_);
  and _75598_ (_29969_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and _75599_ (_29970_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  nor _75600_ (_29971_, _29970_, _29969_);
  and _75601_ (_29972_, _29971_, _29968_);
  and _75602_ (_29973_, _29972_, _29965_);
  and _75603_ (_29974_, _29973_, _29958_);
  and _75604_ (_29975_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and _75605_ (_29976_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor _75606_ (_29977_, _29976_, _29975_);
  and _75607_ (_29978_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and _75608_ (_29979_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor _75609_ (_29980_, _29979_, _29978_);
  and _75610_ (_29981_, _29980_, _29977_);
  and _75611_ (_29982_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and _75612_ (_29983_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and _75613_ (_29984_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or _75614_ (_29985_, _29984_, _29983_);
  nor _75615_ (_29986_, _29985_, _29982_);
  and _75616_ (_29987_, _29986_, _29981_);
  and _75617_ (_29988_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and _75618_ (_29989_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor _75619_ (_29990_, _29989_, _29988_);
  and _75620_ (_29991_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and _75621_ (_29992_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor _75622_ (_29993_, _29992_, _29991_);
  and _75623_ (_29994_, _29993_, _29990_);
  and _75624_ (_29995_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and _75625_ (_29996_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor _75626_ (_29997_, _29996_, _29995_);
  and _75627_ (_29998_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and _75628_ (_29999_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor _75629_ (_30000_, _29999_, _29998_);
  and _75630_ (_30001_, _30000_, _29997_);
  and _75631_ (_30002_, _30001_, _29994_);
  and _75632_ (_30003_, _30002_, _29987_);
  and _75633_ (_30004_, _30003_, _29974_);
  and _75634_ (_30005_, _30004_, _29943_);
  and _75635_ (_30006_, _30005_, _29880_);
  and _75636_ (_30007_, _30006_, _29753_);
  and _75637_ (_30008_, _30007_, _29498_);
  and _75638_ (_30009_, _29491_, iram_op1_reg[3]);
  and _75639_ (_30010_, _30009_, iram_op1_reg[4]);
  nor _75640_ (_30011_, _30009_, iram_op1_reg[4]);
  nor _75641_ (_30012_, _30011_, _30010_);
  and _75642_ (_30013_, _30012_, _30008_);
  nor _75643_ (_30014_, _30012_, _30008_);
  or _75644_ (_30015_, _30014_, _30013_);
  and _75645_ (_30016_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  not _75646_ (_30017_, _30016_);
  and _75647_ (_30018_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and _75648_ (_30019_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  nor _75649_ (_30020_, _30019_, _30018_);
  and _75650_ (_30021_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  and _75651_ (_30022_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  nor _75652_ (_30023_, _30022_, _30021_);
  and _75653_ (_30024_, _30023_, _30020_);
  and _75654_ (_30025_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and _75655_ (_30026_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  nor _75656_ (_30027_, _30026_, _30025_);
  and _75657_ (_30028_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  and _75658_ (_30029_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  nor _75659_ (_30030_, _30029_, _30028_);
  and _75660_ (_30031_, _30030_, _30027_);
  and _75661_ (_30032_, _30031_, _30024_);
  and _75662_ (_30033_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  and _75663_ (_30034_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  nor _75664_ (_30035_, _30034_, _30033_);
  and _75665_ (_30036_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and _75666_ (_30037_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  nor _75667_ (_30038_, _30037_, _30036_);
  and _75668_ (_30039_, _30038_, _30035_);
  and _75669_ (_30040_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  and _75670_ (_30041_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  nor _75671_ (_30042_, _30041_, _30040_);
  and _75672_ (_30043_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and _75673_ (_30044_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  nor _75674_ (_30045_, _30044_, _30043_);
  and _75675_ (_30046_, _30045_, _30042_);
  and _75676_ (_30047_, _30046_, _30039_);
  and _75677_ (_30048_, _30047_, _30032_);
  and _75678_ (_30049_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and _75679_ (_30050_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  nor _75680_ (_30051_, _30050_, _30049_);
  and _75681_ (_30052_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  and _75682_ (_30053_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  nor _75683_ (_30054_, _30053_, _30052_);
  and _75684_ (_30055_, _30054_, _30051_);
  and _75685_ (_30056_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and _75686_ (_30057_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  nor _75687_ (_30058_, _30057_, _30056_);
  and _75688_ (_30059_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  and _75689_ (_30060_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  nor _75690_ (_30061_, _30060_, _30059_);
  and _75691_ (_30062_, _30061_, _30058_);
  and _75692_ (_30063_, _30062_, _30055_);
  and _75693_ (_30064_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  and _75694_ (_30065_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  nor _75695_ (_30066_, _30065_, _30064_);
  and _75696_ (_30067_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  and _75697_ (_30068_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  nor _75698_ (_30069_, _30068_, _30067_);
  and _75699_ (_30070_, _30069_, _30066_);
  and _75700_ (_30071_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  and _75701_ (_30072_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  nor _75702_ (_30073_, _30072_, _30071_);
  and _75703_ (_30074_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and _75704_ (_30075_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  nor _75705_ (_30076_, _30075_, _30074_);
  and _75706_ (_30077_, _30076_, _30073_);
  and _75707_ (_30078_, _30077_, _30070_);
  and _75708_ (_30079_, _30078_, _30063_);
  and _75709_ (_30080_, _30079_, _30048_);
  and _75710_ (_30081_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and _75711_ (_30082_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  nor _75712_ (_30083_, _30082_, _30081_);
  and _75713_ (_30084_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  and _75714_ (_30085_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  nor _75715_ (_30086_, _30085_, _30084_);
  and _75716_ (_30087_, _30086_, _30083_);
  and _75717_ (_30088_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and _75718_ (_30089_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  nor _75719_ (_30090_, _30089_, _30088_);
  and _75720_ (_30091_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and _75721_ (_30092_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  nor _75722_ (_30093_, _30092_, _30091_);
  and _75723_ (_30094_, _30093_, _30090_);
  and _75724_ (_30095_, _30094_, _30087_);
  and _75725_ (_30096_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  and _75726_ (_30097_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  nor _75727_ (_30098_, _30097_, _30096_);
  and _75728_ (_30099_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and _75729_ (_30100_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  nor _75730_ (_30101_, _30100_, _30099_);
  and _75731_ (_30102_, _30101_, _30098_);
  and _75732_ (_30103_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  and _75733_ (_30104_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  nor _75734_ (_30105_, _30104_, _30103_);
  and _75735_ (_30106_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and _75736_ (_30107_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  nor _75737_ (_30108_, _30107_, _30106_);
  and _75738_ (_30109_, _30108_, _30105_);
  and _75739_ (_30110_, _30109_, _30102_);
  and _75740_ (_30111_, _30110_, _30095_);
  and _75741_ (_30112_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and _75742_ (_30113_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  nor _75743_ (_30114_, _30113_, _30112_);
  and _75744_ (_30115_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  and _75745_ (_30116_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  nor _75746_ (_30117_, _30116_, _30115_);
  and _75747_ (_30118_, _30117_, _30114_);
  and _75748_ (_30119_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and _75749_ (_30120_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  nor _75750_ (_30121_, _30120_, _30119_);
  and _75751_ (_30122_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  and _75752_ (_30123_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  nor _75753_ (_30124_, _30123_, _30122_);
  and _75754_ (_30125_, _30124_, _30121_);
  and _75755_ (_30126_, _30125_, _30118_);
  and _75756_ (_30127_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  and _75757_ (_30128_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  nor _75758_ (_30129_, _30128_, _30127_);
  and _75759_ (_30130_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and _75760_ (_30131_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  nor _75761_ (_30132_, _30131_, _30130_);
  and _75762_ (_30133_, _30132_, _30129_);
  and _75763_ (_30134_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  and _75764_ (_30135_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  nor _75765_ (_30136_, _30135_, _30134_);
  and _75766_ (_30137_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  and _75767_ (_30138_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  nor _75768_ (_30139_, _30138_, _30137_);
  and _75769_ (_30140_, _30139_, _30136_);
  and _75770_ (_30141_, _30140_, _30133_);
  and _75771_ (_30142_, _30141_, _30126_);
  and _75772_ (_30143_, _30142_, _30111_);
  and _75773_ (_30144_, _30143_, _30080_);
  and _75774_ (_30145_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  and _75775_ (_30146_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  nor _75776_ (_30147_, _30146_, _30145_);
  and _75777_ (_30148_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and _75778_ (_30149_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  nor _75779_ (_30150_, _30149_, _30148_);
  and _75780_ (_30151_, _30150_, _30147_);
  and _75781_ (_30152_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and _75782_ (_30153_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  nor _75783_ (_30154_, _30153_, _30152_);
  and _75784_ (_30155_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and _75785_ (_30156_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  nor _75786_ (_30157_, _30156_, _30155_);
  and _75787_ (_30158_, _30157_, _30154_);
  and _75788_ (_30159_, _30158_, _30151_);
  and _75789_ (_30160_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  and _75790_ (_30161_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  nor _75791_ (_30162_, _30161_, _30160_);
  and _75792_ (_30163_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and _75793_ (_30164_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  nor _75794_ (_30165_, _30164_, _30163_);
  and _75795_ (_30166_, _30165_, _30162_);
  and _75796_ (_30167_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  and _75797_ (_30168_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  nor _75798_ (_30169_, _30168_, _30167_);
  and _75799_ (_30170_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and _75800_ (_30171_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  nor _75801_ (_30172_, _30171_, _30170_);
  and _75802_ (_30173_, _30172_, _30169_);
  and _75803_ (_30174_, _30173_, _30166_);
  and _75804_ (_30175_, _30174_, _30159_);
  and _75805_ (_30176_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and _75806_ (_30177_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  nor _75807_ (_30178_, _30177_, _30176_);
  and _75808_ (_30179_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  and _75809_ (_30180_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  nor _75810_ (_30181_, _30180_, _30179_);
  and _75811_ (_30182_, _30181_, _30178_);
  and _75812_ (_30183_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and _75813_ (_30184_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  nor _75814_ (_30185_, _30184_, _30183_);
  and _75815_ (_30186_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  and _75816_ (_30187_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  nor _75817_ (_30188_, _30187_, _30186_);
  and _75818_ (_30189_, _30188_, _30185_);
  and _75819_ (_30190_, _30189_, _30182_);
  and _75820_ (_30191_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  and _75821_ (_30192_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  nor _75822_ (_30193_, _30192_, _30191_);
  and _75823_ (_30194_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and _75824_ (_30195_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  nor _75825_ (_30196_, _30195_, _30194_);
  and _75826_ (_30197_, _30196_, _30193_);
  and _75827_ (_30198_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  and _75828_ (_30199_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  nor _75829_ (_30200_, _30199_, _30198_);
  and _75830_ (_30201_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and _75831_ (_30202_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  nor _75832_ (_30203_, _30202_, _30201_);
  and _75833_ (_30204_, _30203_, _30200_);
  and _75834_ (_30205_, _30204_, _30197_);
  and _75835_ (_30206_, _30205_, _30190_);
  and _75836_ (_30207_, _30206_, _30175_);
  and _75837_ (_30208_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and _75838_ (_30209_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  nor _75839_ (_30210_, _30209_, _30208_);
  and _75840_ (_30211_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  and _75841_ (_30212_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  nor _75842_ (_30213_, _30212_, _30211_);
  and _75843_ (_30214_, _30213_, _30210_);
  and _75844_ (_30215_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and _75845_ (_30216_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  nor _75846_ (_30217_, _30216_, _30215_);
  and _75847_ (_30218_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  and _75848_ (_30219_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  nor _75849_ (_30220_, _30219_, _30218_);
  and _75850_ (_30221_, _30220_, _30217_);
  and _75851_ (_30222_, _30221_, _30214_);
  and _75852_ (_30223_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  and _75853_ (_30224_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  nor _75854_ (_30225_, _30224_, _30223_);
  and _75855_ (_30226_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and _75856_ (_30227_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  nor _75857_ (_30228_, _30227_, _30226_);
  and _75858_ (_30229_, _30228_, _30225_);
  and _75859_ (_30230_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  and _75860_ (_30231_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  nor _75861_ (_30232_, _30231_, _30230_);
  and _75862_ (_30233_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and _75863_ (_30234_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  nor _75864_ (_30235_, _30234_, _30233_);
  and _75865_ (_30236_, _30235_, _30232_);
  and _75866_ (_30237_, _30236_, _30229_);
  and _75867_ (_30238_, _30237_, _30222_);
  and _75868_ (_30239_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and _75869_ (_30240_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  nor _75870_ (_30241_, _30240_, _30239_);
  and _75871_ (_30242_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  and _75872_ (_30243_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  nor _75873_ (_30244_, _30243_, _30242_);
  and _75874_ (_30245_, _30244_, _30241_);
  and _75875_ (_30246_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  and _75876_ (_30247_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  nor _75877_ (_30248_, _30247_, _30246_);
  and _75878_ (_30249_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and _75879_ (_30250_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  nor _75880_ (_30251_, _30250_, _30249_);
  and _75881_ (_30252_, _30251_, _30248_);
  and _75882_ (_30253_, _30252_, _30245_);
  and _75883_ (_30254_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  and _75884_ (_30255_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  nor _75885_ (_30256_, _30255_, _30254_);
  and _75886_ (_30257_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  and _75887_ (_30258_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  nor _75888_ (_30259_, _30258_, _30257_);
  and _75889_ (_30260_, _30259_, _30256_);
  and _75890_ (_30261_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  and _75891_ (_30262_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  nor _75892_ (_30263_, _30262_, _30261_);
  and _75893_ (_30264_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and _75894_ (_30265_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  nor _75895_ (_30266_, _30265_, _30264_);
  and _75896_ (_30267_, _30266_, _30263_);
  and _75897_ (_30268_, _30267_, _30260_);
  and _75898_ (_30269_, _30268_, _30253_);
  and _75899_ (_30270_, _30269_, _30238_);
  and _75900_ (_30271_, _30270_, _30207_);
  and _75901_ (_30272_, _30271_, _30144_);
  and _75902_ (_30273_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and _75903_ (_30274_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  nor _75904_ (_30275_, _30274_, _30273_);
  and _75905_ (_30276_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and _75906_ (_30277_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  nor _75907_ (_30278_, _30277_, _30276_);
  and _75908_ (_30279_, _30278_, _30275_);
  and _75909_ (_30280_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and _75910_ (_30281_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  nor _75911_ (_30282_, _30281_, _30280_);
  and _75912_ (_30283_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  and _75913_ (_30284_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  nor _75914_ (_30285_, _30284_, _30283_);
  and _75915_ (_30286_, _30285_, _30282_);
  and _75916_ (_30287_, _30286_, _30279_);
  and _75917_ (_30288_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  and _75918_ (_30289_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  nor _75919_ (_30290_, _30289_, _30288_);
  and _75920_ (_30291_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and _75921_ (_30292_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  nor _75922_ (_30293_, _30292_, _30291_);
  and _75923_ (_30294_, _30293_, _30290_);
  and _75924_ (_30295_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  and _75925_ (_30296_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  nor _75926_ (_30297_, _30296_, _30295_);
  and _75927_ (_30298_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and _75928_ (_30299_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  nor _75929_ (_30300_, _30299_, _30298_);
  and _75930_ (_30301_, _30300_, _30297_);
  and _75931_ (_30302_, _30301_, _30294_);
  and _75932_ (_30303_, _30302_, _30287_);
  and _75933_ (_30304_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and _75934_ (_30305_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  nor _75935_ (_30306_, _30305_, _30304_);
  and _75936_ (_30307_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  and _75937_ (_30308_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  nor _75938_ (_30309_, _30308_, _30307_);
  and _75939_ (_30310_, _30309_, _30306_);
  and _75940_ (_30311_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and _75941_ (_30312_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  nor _75942_ (_30313_, _30312_, _30311_);
  and _75943_ (_30314_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  and _75944_ (_30315_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  nor _75945_ (_30316_, _30315_, _30314_);
  and _75946_ (_30317_, _30316_, _30313_);
  and _75947_ (_30318_, _30317_, _30310_);
  and _75948_ (_30319_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  and _75949_ (_30320_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  nor _75950_ (_30321_, _30320_, _30319_);
  and _75951_ (_30322_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and _75952_ (_30323_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  nor _75953_ (_30324_, _30323_, _30322_);
  and _75954_ (_30325_, _30324_, _30321_);
  and _75955_ (_30326_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  and _75956_ (_30327_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  nor _75957_ (_30328_, _30327_, _30326_);
  and _75958_ (_30329_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and _75959_ (_30330_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  nor _75960_ (_30331_, _30330_, _30329_);
  and _75961_ (_30332_, _30331_, _30328_);
  and _75962_ (_30333_, _30332_, _30325_);
  and _75963_ (_30334_, _30333_, _30318_);
  and _75964_ (_30335_, _30334_, _30303_);
  and _75965_ (_30336_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and _75966_ (_30337_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  nor _75967_ (_30338_, _30337_, _30336_);
  and _75968_ (_30339_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  and _75969_ (_30340_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  nor _75970_ (_30341_, _30340_, _30339_);
  and _75971_ (_30342_, _30341_, _30338_);
  and _75972_ (_30343_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and _75973_ (_30344_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  nor _75974_ (_30345_, _30344_, _30343_);
  and _75975_ (_30346_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and _75976_ (_30347_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  nor _75977_ (_30348_, _30347_, _30346_);
  and _75978_ (_30349_, _30348_, _30345_);
  and _75979_ (_30350_, _30349_, _30342_);
  and _75980_ (_30351_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  and _75981_ (_30352_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  nor _75982_ (_30353_, _30352_, _30351_);
  and _75983_ (_30354_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and _75984_ (_30355_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  nor _75985_ (_30356_, _30355_, _30354_);
  and _75986_ (_30357_, _30356_, _30353_);
  and _75987_ (_30358_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  and _75988_ (_30359_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  nor _75989_ (_30360_, _30359_, _30358_);
  and _75990_ (_30361_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and _75991_ (_30362_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  nor _75992_ (_30363_, _30362_, _30361_);
  and _75993_ (_30364_, _30363_, _30360_);
  and _75994_ (_30365_, _30364_, _30357_);
  and _75995_ (_30366_, _30365_, _30350_);
  and _75996_ (_30367_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  and _75997_ (_30368_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  nor _75998_ (_30369_, _30368_, _30367_);
  and _75999_ (_30370_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and _76000_ (_30371_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  nor _76001_ (_30372_, _30371_, _30370_);
  and _76002_ (_30373_, _30372_, _30369_);
  and _76003_ (_30374_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  and _76004_ (_30375_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  nor _76005_ (_30376_, _30375_, _30374_);
  and _76006_ (_30377_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  and _76007_ (_30378_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  nor _76008_ (_30379_, _30378_, _30377_);
  and _76009_ (_30380_, _30379_, _30376_);
  and _76010_ (_30381_, _30380_, _30373_);
  and _76011_ (_30382_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and _76012_ (_30383_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  nor _76013_ (_30384_, _30383_, _30382_);
  and _76014_ (_30385_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  and _76015_ (_30386_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  nor _76016_ (_30387_, _30386_, _30385_);
  and _76017_ (_30388_, _30387_, _30384_);
  and _76018_ (_30389_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and _76019_ (_30390_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  nor _76020_ (_30391_, _30390_, _30389_);
  and _76021_ (_30392_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  and _76022_ (_30393_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  nor _76023_ (_30394_, _30393_, _30392_);
  and _76024_ (_30395_, _30394_, _30391_);
  and _76025_ (_30396_, _30395_, _30388_);
  and _76026_ (_30397_, _30396_, _30381_);
  and _76027_ (_30398_, _30397_, _30366_);
  and _76028_ (_30399_, _30398_, _30335_);
  and _76029_ (_30400_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  and _76030_ (_30401_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  nor _76031_ (_30402_, _30401_, _30400_);
  and _76032_ (_30403_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and _76033_ (_30404_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  nor _76034_ (_30405_, _30404_, _30403_);
  and _76035_ (_30406_, _30405_, _30402_);
  and _76036_ (_30407_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  and _76037_ (_30408_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  nor _76038_ (_30409_, _30408_, _30407_);
  and _76039_ (_30410_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and _76040_ (_30411_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  nor _76041_ (_30412_, _30411_, _30410_);
  and _76042_ (_30413_, _30412_, _30409_);
  and _76043_ (_30414_, _30413_, _30406_);
  and _76044_ (_30415_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and _76045_ (_30416_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  nor _76046_ (_30417_, _30416_, _30415_);
  and _76047_ (_30418_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  and _76048_ (_30419_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  nor _76049_ (_30420_, _30419_, _30418_);
  and _76050_ (_30421_, _30420_, _30417_);
  and _76051_ (_30422_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and _76052_ (_30423_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  nor _76053_ (_30424_, _30423_, _30422_);
  and _76054_ (_30425_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  and _76055_ (_30426_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  nor _76056_ (_30427_, _30426_, _30425_);
  and _76057_ (_30428_, _30427_, _30424_);
  and _76058_ (_30429_, _30428_, _30421_);
  and _76059_ (_30430_, _30429_, _30414_);
  and _76060_ (_30431_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and _76061_ (_30432_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  nor _76062_ (_30433_, _30432_, _30431_);
  and _76063_ (_30434_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  and _76064_ (_30435_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  nor _76065_ (_30436_, _30435_, _30434_);
  and _76066_ (_30437_, _30436_, _30433_);
  and _76067_ (_30438_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  and _76068_ (_30439_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  nor _76069_ (_30440_, _30439_, _30438_);
  and _76070_ (_30441_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and _76071_ (_30442_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  nor _76072_ (_30443_, _30442_, _30441_);
  and _76073_ (_30444_, _30443_, _30440_);
  and _76074_ (_30445_, _30444_, _30437_);
  and _76075_ (_30446_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  and _76076_ (_30447_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  nor _76077_ (_30448_, _30447_, _30446_);
  and _76078_ (_30449_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and _76079_ (_30450_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  nor _76080_ (_30451_, _30450_, _30449_);
  and _76081_ (_30452_, _30451_, _30448_);
  and _76082_ (_30453_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  and _76083_ (_30454_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  nor _76084_ (_30455_, _30454_, _30453_);
  and _76085_ (_30456_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and _76086_ (_30457_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  nor _76087_ (_30458_, _30457_, _30456_);
  and _76088_ (_30459_, _30458_, _30455_);
  and _76089_ (_30460_, _30459_, _30452_);
  and _76090_ (_30461_, _30460_, _30445_);
  and _76091_ (_30462_, _30461_, _30430_);
  and _76092_ (_30463_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and _76093_ (_30464_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  nor _76094_ (_30465_, _30464_, _30463_);
  and _76095_ (_30466_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  and _76096_ (_30467_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  nor _76097_ (_30468_, _30467_, _30466_);
  and _76098_ (_30469_, _30468_, _30465_);
  and _76099_ (_30470_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and _76100_ (_30471_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  nor _76101_ (_30472_, _30471_, _30470_);
  and _76102_ (_30473_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  and _76103_ (_30474_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  nor _76104_ (_30475_, _30474_, _30473_);
  and _76105_ (_30476_, _30475_, _30472_);
  and _76106_ (_30477_, _30476_, _30469_);
  and _76107_ (_30478_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  and _76108_ (_30479_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  nor _76109_ (_30480_, _30479_, _30478_);
  and _76110_ (_30481_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and _76111_ (_30482_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  nor _76112_ (_30483_, _30482_, _30481_);
  and _76113_ (_30484_, _30483_, _30480_);
  and _76114_ (_30485_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  and _76115_ (_30486_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  nor _76116_ (_30487_, _30486_, _30485_);
  and _76117_ (_30488_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and _76118_ (_30489_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor _76119_ (_30490_, _30489_, _30488_);
  and _76120_ (_30491_, _30490_, _30487_);
  and _76121_ (_30492_, _30491_, _30484_);
  and _76122_ (_30493_, _30492_, _30477_);
  and _76123_ (_30494_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and _76124_ (_30495_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor _76125_ (_30496_, _30495_, _30494_);
  and _76126_ (_30497_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and _76127_ (_30498_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor _76128_ (_30499_, _30498_, _30497_);
  and _76129_ (_30500_, _30499_, _30496_);
  and _76130_ (_30501_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and _76131_ (_30502_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor _76132_ (_30503_, _30502_, _30501_);
  and _76133_ (_30504_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and _76134_ (_30505_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor _76135_ (_30506_, _30505_, _30504_);
  and _76136_ (_30507_, _30506_, _30503_);
  and _76137_ (_30508_, _30507_, _30500_);
  and _76138_ (_30509_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and _76139_ (_30510_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and _76140_ (_30511_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _76141_ (_30512_, _30511_, _30510_);
  nor _76142_ (_30513_, _30512_, _30509_);
  and _76143_ (_30514_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and _76144_ (_30515_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor _76145_ (_30516_, _30515_, _30514_);
  and _76146_ (_30517_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and _76147_ (_30518_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor _76148_ (_30519_, _30518_, _30517_);
  and _76149_ (_30520_, _30519_, _30516_);
  and _76150_ (_30521_, _30520_, _30513_);
  and _76151_ (_30522_, _30521_, _30508_);
  and _76152_ (_30523_, _30522_, _30493_);
  and _76153_ (_30524_, _30523_, _30462_);
  and _76154_ (_30525_, _30524_, _30399_);
  and _76155_ (_30526_, _30525_, _30272_);
  and _76156_ (_30527_, _30526_, _30017_);
  nor _76157_ (_30528_, _29491_, iram_op1_reg[3]);
  nor _76158_ (_30529_, _30528_, _30009_);
  and _76159_ (_30530_, _30529_, _30527_);
  and _76160_ (_30531_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  not _76161_ (_30532_, _30531_);
  and _76162_ (_30533_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and _76163_ (_30534_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or _76164_ (_30535_, _30534_, _30533_);
  and _76165_ (_30536_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  and _76166_ (_30537_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  or _76167_ (_30538_, _30537_, _30536_);
  or _76168_ (_30539_, _30538_, _30535_);
  and _76169_ (_30540_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  and _76170_ (_30541_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or _76171_ (_30542_, _30541_, _30540_);
  and _76172_ (_30543_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and _76173_ (_30544_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  or _76174_ (_30545_, _30544_, _30543_);
  or _76175_ (_30546_, _30545_, _30542_);
  or _76176_ (_30547_, _30546_, _30539_);
  and _76177_ (_30548_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and _76178_ (_30549_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or _76179_ (_30550_, _30549_, _30548_);
  and _76180_ (_30551_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  and _76181_ (_30552_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or _76182_ (_30553_, _30552_, _30551_);
  or _76183_ (_30554_, _30553_, _30550_);
  and _76184_ (_30555_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and _76185_ (_30556_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  or _76186_ (_30557_, _30556_, _30555_);
  and _76187_ (_30558_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and _76188_ (_30559_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or _76189_ (_30560_, _30559_, _30558_);
  or _76190_ (_30561_, _30560_, _30557_);
  or _76191_ (_30562_, _30561_, _30554_);
  or _76192_ (_30563_, _30562_, _30547_);
  and _76193_ (_30564_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and _76194_ (_30565_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or _76195_ (_30566_, _30565_, _30564_);
  and _76196_ (_30567_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  and _76197_ (_30568_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  or _76198_ (_30569_, _30568_, _30567_);
  or _76199_ (_30570_, _30569_, _30566_);
  and _76200_ (_30571_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and _76201_ (_30572_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  or _76202_ (_30573_, _30572_, _30571_);
  and _76203_ (_30574_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  and _76204_ (_30575_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or _76205_ (_30576_, _30575_, _30574_);
  or _76206_ (_30577_, _30576_, _30573_);
  or _76207_ (_30578_, _30577_, _30570_);
  and _76208_ (_30579_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  and _76209_ (_30580_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or _76210_ (_30581_, _30580_, _30579_);
  and _76211_ (_30582_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  and _76212_ (_30583_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or _76213_ (_30584_, _30583_, _30582_);
  or _76214_ (_30585_, _30584_, _30581_);
  and _76215_ (_30586_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and _76216_ (_30587_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or _76217_ (_30588_, _30587_, _30586_);
  and _76218_ (_30589_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  and _76219_ (_30590_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or _76220_ (_30591_, _30590_, _30589_);
  or _76221_ (_30592_, _30591_, _30588_);
  or _76222_ (_30593_, _30592_, _30585_);
  or _76223_ (_30594_, _30593_, _30578_);
  or _76224_ (_30595_, _30594_, _30563_);
  and _76225_ (_30596_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and _76226_ (_30597_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  or _76227_ (_30598_, _30597_, _30596_);
  and _76228_ (_30599_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and _76229_ (_30600_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or _76230_ (_30601_, _30600_, _30599_);
  or _76231_ (_30602_, _30601_, _30598_);
  and _76232_ (_30603_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and _76233_ (_30604_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor _76234_ (_30605_, _30604_, _30603_);
  and _76235_ (_30606_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and _76236_ (_30607_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  nor _76237_ (_30608_, _30607_, _30606_);
  nand _76238_ (_30609_, _30608_, _30605_);
  or _76239_ (_30610_, _30609_, _30602_);
  and _76240_ (_30611_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  and _76241_ (_30612_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or _76242_ (_30613_, _30612_, _30611_);
  and _76243_ (_30614_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  and _76244_ (_30615_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or _76245_ (_30616_, _30615_, _30614_);
  or _76246_ (_30617_, _30616_, _30613_);
  and _76247_ (_30618_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  and _76248_ (_30619_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or _76249_ (_30620_, _30619_, _30618_);
  and _76250_ (_30621_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and _76251_ (_30622_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or _76252_ (_30623_, _30622_, _30621_);
  or _76253_ (_30624_, _30623_, _30620_);
  or _76254_ (_30625_, _30624_, _30617_);
  or _76255_ (_30626_, _30625_, _30610_);
  and _76256_ (_30627_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  and _76257_ (_30628_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  or _76258_ (_30629_, _30628_, _30627_);
  and _76259_ (_30630_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and _76260_ (_30631_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or _76261_ (_30632_, _30631_, _30630_);
  or _76262_ (_30633_, _30632_, _30629_);
  and _76263_ (_30634_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  and _76264_ (_30635_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  nor _76265_ (_30636_, _30635_, _30634_);
  and _76266_ (_30637_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and _76267_ (_30638_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  nor _76268_ (_30639_, _30638_, _30637_);
  nand _76269_ (_30640_, _30639_, _30636_);
  or _76270_ (_30641_, _30640_, _30633_);
  and _76271_ (_30642_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and _76272_ (_30643_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or _76273_ (_30644_, _30643_, _30642_);
  and _76274_ (_30645_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and _76275_ (_30646_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or _76276_ (_30647_, _30646_, _30645_);
  or _76277_ (_30648_, _30647_, _30644_);
  and _76278_ (_30649_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and _76279_ (_30650_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or _76280_ (_30651_, _30650_, _30649_);
  and _76281_ (_30652_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  and _76282_ (_30653_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or _76283_ (_30654_, _30653_, _30652_);
  or _76284_ (_30655_, _30654_, _30651_);
  or _76285_ (_30656_, _30655_, _30648_);
  or _76286_ (_30657_, _30656_, _30641_);
  or _76287_ (_30658_, _30657_, _30626_);
  or _76288_ (_30659_, _30658_, _30595_);
  and _76289_ (_30660_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and _76290_ (_30661_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  or _76291_ (_30662_, _30661_, _30660_);
  and _76292_ (_30663_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and _76293_ (_30664_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or _76294_ (_30665_, _30664_, _30663_);
  or _76295_ (_30666_, _30665_, _30662_);
  and _76296_ (_30667_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  and _76297_ (_30668_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or _76298_ (_30669_, _30668_, _30667_);
  and _76299_ (_30670_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and _76300_ (_30671_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or _76301_ (_30672_, _30671_, _30670_);
  or _76302_ (_30673_, _30672_, _30669_);
  or _76303_ (_30674_, _30673_, _30666_);
  and _76304_ (_30675_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and _76305_ (_30676_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or _76306_ (_30677_, _30676_, _30675_);
  and _76307_ (_30678_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and _76308_ (_30679_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  or _76309_ (_30680_, _30679_, _30678_);
  or _76310_ (_30681_, _30680_, _30677_);
  and _76311_ (_30682_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and _76312_ (_30683_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  nor _76313_ (_30684_, _30683_, _30682_);
  and _76314_ (_30685_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  and _76315_ (_30686_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  nor _76316_ (_30687_, _30686_, _30685_);
  nand _76317_ (_30688_, _30687_, _30684_);
  or _76318_ (_30689_, _30688_, _30681_);
  or _76319_ (_30690_, _30689_, _30674_);
  and _76320_ (_30691_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and _76321_ (_30692_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or _76322_ (_30693_, _30692_, _30691_);
  and _76323_ (_30694_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and _76324_ (_30695_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or _76325_ (_30696_, _30695_, _30694_);
  or _76326_ (_30697_, _30696_, _30693_);
  and _76327_ (_30698_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  and _76328_ (_30699_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  nor _76329_ (_30700_, _30699_, _30698_);
  and _76330_ (_30701_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and _76331_ (_30702_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  nor _76332_ (_30703_, _30702_, _30701_);
  nand _76333_ (_30704_, _30703_, _30700_);
  or _76334_ (_30705_, _30704_, _30697_);
  and _76335_ (_30706_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and _76336_ (_30707_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or _76337_ (_30708_, _30707_, _30706_);
  and _76338_ (_30709_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  and _76339_ (_30710_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or _76340_ (_30711_, _30710_, _30709_);
  or _76341_ (_30712_, _30711_, _30708_);
  and _76342_ (_30713_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  and _76343_ (_30714_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  or _76344_ (_30715_, _30714_, _30713_);
  and _76345_ (_30716_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  and _76346_ (_30717_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or _76347_ (_30718_, _30717_, _30716_);
  or _76348_ (_30719_, _30718_, _30715_);
  or _76349_ (_30720_, _30719_, _30712_);
  or _76350_ (_30721_, _30720_, _30705_);
  or _76351_ (_30722_, _30721_, _30690_);
  and _76352_ (_30723_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and _76353_ (_30724_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor _76354_ (_30725_, _30724_, _30723_);
  and _76355_ (_30726_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  and _76356_ (_30727_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  nor _76357_ (_30728_, _30727_, _30726_);
  nand _76358_ (_30729_, _30728_, _30725_);
  and _76359_ (_30730_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and _76360_ (_30731_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  nor _76361_ (_30732_, _30731_, _30730_);
  and _76362_ (_30733_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  and _76363_ (_30734_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  nor _76364_ (_30735_, _30734_, _30733_);
  nand _76365_ (_30736_, _30735_, _30732_);
  or _76366_ (_30737_, _30736_, _30729_);
  and _76367_ (_30738_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  and _76368_ (_30739_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or _76369_ (_30740_, _30739_, _30738_);
  and _76370_ (_30741_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  and _76371_ (_30742_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or _76372_ (_30743_, _30742_, _30741_);
  or _76373_ (_30744_, _30743_, _30740_);
  and _76374_ (_30745_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  and _76375_ (_30746_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  or _76376_ (_30747_, _30746_, _30745_);
  and _76377_ (_30748_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and _76378_ (_30749_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or _76379_ (_30750_, _30749_, _30748_);
  or _76380_ (_30751_, _30750_, _30747_);
  or _76381_ (_30752_, _30751_, _30744_);
  or _76382_ (_30753_, _30752_, _30737_);
  and _76383_ (_30754_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and _76384_ (_30755_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or _76385_ (_30756_, _30755_, _30754_);
  and _76386_ (_30757_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and _76387_ (_30758_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or _76388_ (_30759_, _30758_, _30757_);
  or _76389_ (_30760_, _30759_, _30756_);
  and _76390_ (_30761_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and _76391_ (_30762_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or _76392_ (_30763_, _30762_, _30761_);
  and _76393_ (_30764_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and _76394_ (_30765_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  or _76395_ (_30766_, _30765_, _30764_);
  or _76396_ (_30767_, _30766_, _30763_);
  or _76397_ (_30768_, _30767_, _30760_);
  and _76398_ (_30769_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  and _76399_ (_30770_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  or _76400_ (_30771_, _30770_, _30769_);
  and _76401_ (_30772_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and _76402_ (_30773_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or _76403_ (_30774_, _30773_, _30772_);
  or _76404_ (_30775_, _30774_, _30771_);
  and _76405_ (_30776_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and _76406_ (_30777_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  or _76407_ (_30778_, _30777_, _30776_);
  and _76408_ (_30779_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  and _76409_ (_30780_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or _76410_ (_30781_, _30780_, _30779_);
  or _76411_ (_30782_, _30781_, _30778_);
  or _76412_ (_30783_, _30782_, _30775_);
  or _76413_ (_30784_, _30783_, _30768_);
  or _76414_ (_30785_, _30784_, _30753_);
  or _76415_ (_30786_, _30785_, _30722_);
  or _76416_ (_30787_, _30786_, _30659_);
  and _76417_ (_30788_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and _76418_ (_30789_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or _76419_ (_30790_, _30789_, _30788_);
  and _76420_ (_30791_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  and _76421_ (_30792_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or _76422_ (_30793_, _30792_, _30791_);
  or _76423_ (_30794_, _30793_, _30790_);
  and _76424_ (_30795_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  and _76425_ (_30796_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or _76426_ (_30797_, _30796_, _30795_);
  and _76427_ (_30798_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and _76428_ (_30799_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or _76429_ (_30800_, _30799_, _30798_);
  or _76430_ (_30801_, _30800_, _30797_);
  or _76431_ (_30802_, _30801_, _30794_);
  and _76432_ (_30803_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  and _76433_ (_30804_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  or _76434_ (_30805_, _30804_, _30803_);
  and _76435_ (_30806_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and _76436_ (_30807_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  or _76437_ (_30808_, _30807_, _30806_);
  or _76438_ (_30809_, _30808_, _30805_);
  and _76439_ (_30810_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and _76440_ (_30811_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  or _76441_ (_30812_, _30811_, _30810_);
  and _76442_ (_30813_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  and _76443_ (_30814_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or _76444_ (_30815_, _30814_, _30813_);
  or _76445_ (_30816_, _30815_, _30812_);
  or _76446_ (_30817_, _30816_, _30809_);
  or _76447_ (_30818_, _30817_, _30802_);
  and _76448_ (_30819_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  and _76449_ (_30820_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  or _76450_ (_30821_, _30820_, _30819_);
  and _76451_ (_30822_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and _76452_ (_30823_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or _76453_ (_30824_, _30823_, _30822_);
  or _76454_ (_30825_, _30824_, _30821_);
  and _76455_ (_30826_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  and _76456_ (_30827_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  or _76457_ (_30828_, _30827_, _30826_);
  and _76458_ (_30829_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  and _76459_ (_30830_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or _76460_ (_30831_, _30830_, _30829_);
  or _76461_ (_30832_, _30831_, _30828_);
  or _76462_ (_30833_, _30832_, _30825_);
  and _76463_ (_30834_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and _76464_ (_30835_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  or _76465_ (_30836_, _30835_, _30834_);
  and _76466_ (_30837_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and _76467_ (_30838_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or _76468_ (_30839_, _30838_, _30837_);
  or _76469_ (_30840_, _30839_, _30836_);
  and _76470_ (_30841_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  and _76471_ (_30842_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  nor _76472_ (_30843_, _30842_, _30841_);
  and _76473_ (_30844_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and _76474_ (_30845_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor _76475_ (_30846_, _30845_, _30844_);
  nand _76476_ (_30847_, _30846_, _30843_);
  or _76477_ (_30848_, _30847_, _30840_);
  or _76478_ (_30849_, _30848_, _30833_);
  or _76479_ (_30850_, _30849_, _30818_);
  and _76480_ (_30851_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and _76481_ (_30852_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  nor _76482_ (_30853_, _30852_, _30851_);
  and _76483_ (_30854_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  and _76484_ (_30855_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  nor _76485_ (_30856_, _30855_, _30854_);
  nand _76486_ (_30857_, _30856_, _30853_);
  and _76487_ (_30858_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  and _76488_ (_30859_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  or _76489_ (_30860_, _30859_, _30858_);
  and _76490_ (_30861_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and _76491_ (_30862_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  or _76492_ (_30863_, _30862_, _30861_);
  or _76493_ (_30864_, _30863_, _30860_);
  or _76494_ (_30865_, _30864_, _30857_);
  and _76495_ (_30866_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  and _76496_ (_30867_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  and _76497_ (_30868_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or _76498_ (_30869_, _30868_, _30867_);
  or _76499_ (_30870_, _30869_, _30866_);
  and _76500_ (_30871_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and _76501_ (_30872_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  nor _76502_ (_30873_, _30872_, _30871_);
  and _76503_ (_30874_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  and _76504_ (_30875_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  nor _76505_ (_30876_, _30875_, _30874_);
  nand _76506_ (_30877_, _30876_, _30873_);
  or _76507_ (_30878_, _30877_, _30870_);
  or _76508_ (_30879_, _30878_, _30865_);
  and _76509_ (_30880_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and _76510_ (_30881_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or _76511_ (_30882_, _30881_, _30880_);
  and _76512_ (_30883_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  and _76513_ (_30884_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or _76514_ (_30885_, _30884_, _30883_);
  or _76515_ (_30886_, _30885_, _30882_);
  and _76516_ (_30887_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  and _76517_ (_30888_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or _76518_ (_30889_, _30888_, _30887_);
  and _76519_ (_30890_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  and _76520_ (_30891_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  or _76521_ (_30892_, _30891_, _30890_);
  or _76522_ (_30893_, _30892_, _30889_);
  or _76523_ (_30894_, _30893_, _30886_);
  and _76524_ (_30895_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  and _76525_ (_30896_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or _76526_ (_30897_, _30896_, _30895_);
  and _76527_ (_30898_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  and _76528_ (_30899_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or _76529_ (_30900_, _30899_, _30898_);
  or _76530_ (_30901_, _30900_, _30897_);
  and _76531_ (_30902_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and _76532_ (_30903_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or _76533_ (_30904_, _30903_, _30902_);
  and _76534_ (_30905_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and _76535_ (_30906_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  or _76536_ (_30907_, _30906_, _30905_);
  or _76537_ (_30908_, _30907_, _30904_);
  or _76538_ (_30909_, _30908_, _30901_);
  or _76539_ (_30910_, _30909_, _30894_);
  or _76540_ (_30911_, _30910_, _30879_);
  or _76541_ (_30912_, _30911_, _30850_);
  and _76542_ (_30913_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  and _76543_ (_30914_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or _76544_ (_30915_, _30914_, _30913_);
  and _76545_ (_30916_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and _76546_ (_30917_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or _76547_ (_30918_, _30917_, _30916_);
  or _76548_ (_30919_, _30918_, _30915_);
  and _76549_ (_30920_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and _76550_ (_30921_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or _76551_ (_30922_, _30921_, _30920_);
  and _76552_ (_30923_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  and _76553_ (_30924_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  or _76554_ (_30925_, _30924_, _30923_);
  or _76555_ (_30926_, _30925_, _30922_);
  or _76556_ (_30927_, _30926_, _30919_);
  and _76557_ (_30928_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and _76558_ (_30929_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or _76559_ (_30930_, _30929_, _30928_);
  and _76560_ (_30931_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  and _76561_ (_30932_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or _76562_ (_30933_, _30932_, _30931_);
  or _76563_ (_30934_, _30933_, _30930_);
  and _76564_ (_30935_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and _76565_ (_30936_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or _76566_ (_30937_, _30936_, _30935_);
  and _76567_ (_30938_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and _76568_ (_30939_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or _76569_ (_30940_, _30939_, _30938_);
  or _76570_ (_30941_, _30940_, _30937_);
  or _76571_ (_30942_, _30941_, _30934_);
  or _76572_ (_30943_, _30942_, _30927_);
  and _76573_ (_30944_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and _76574_ (_30945_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or _76575_ (_30946_, _30945_, _30944_);
  and _76576_ (_30947_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  and _76577_ (_30948_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or _76578_ (_30949_, _30948_, _30947_);
  or _76579_ (_30950_, _30949_, _30946_);
  and _76580_ (_30951_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and _76581_ (_30952_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or _76582_ (_30953_, _30952_, _30951_);
  and _76583_ (_30954_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and _76584_ (_30955_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  or _76585_ (_30956_, _30955_, _30954_);
  or _76586_ (_30957_, _30956_, _30953_);
  or _76587_ (_30958_, _30957_, _30950_);
  and _76588_ (_30959_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  and _76589_ (_30960_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or _76590_ (_30961_, _30960_, _30959_);
  and _76591_ (_30962_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  and _76592_ (_30963_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or _76593_ (_30964_, _30963_, _30962_);
  or _76594_ (_30965_, _30964_, _30961_);
  and _76595_ (_30966_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  and _76596_ (_30967_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or _76597_ (_30968_, _30967_, _30966_);
  and _76598_ (_30969_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and _76599_ (_30970_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or _76600_ (_30971_, _30970_, _30969_);
  or _76601_ (_30972_, _30971_, _30968_);
  or _76602_ (_30973_, _30972_, _30965_);
  or _76603_ (_30974_, _30973_, _30958_);
  or _76604_ (_30975_, _30974_, _30943_);
  and _76605_ (_30976_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and _76606_ (_30977_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or _76607_ (_30978_, _30977_, _30976_);
  and _76608_ (_30979_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  and _76609_ (_30980_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or _76610_ (_30981_, _30980_, _30979_);
  or _76611_ (_30982_, _30981_, _30978_);
  and _76612_ (_30983_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and _76613_ (_30984_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or _76614_ (_30985_, _30984_, _30983_);
  and _76615_ (_30986_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  and _76616_ (_30987_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or _76617_ (_30988_, _30987_, _30986_);
  or _76618_ (_30989_, _30988_, _30985_);
  or _76619_ (_30990_, _30989_, _30982_);
  and _76620_ (_30991_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and _76621_ (_30992_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  or _76622_ (_30993_, _30992_, _30991_);
  and _76623_ (_30994_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  and _76624_ (_30995_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or _76625_ (_30996_, _30995_, _30994_);
  or _76626_ (_30997_, _30996_, _30993_);
  and _76627_ (_30998_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  and _76628_ (_30999_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  or _76629_ (_31000_, _30999_, _30998_);
  and _76630_ (_31001_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and _76631_ (_31002_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or _76632_ (_31003_, _31002_, _31001_);
  or _76633_ (_31004_, _31003_, _31000_);
  or _76634_ (_31005_, _31004_, _30997_);
  or _76635_ (_31006_, _31005_, _30990_);
  and _76636_ (_31007_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and _76637_ (_31008_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  or _76638_ (_31009_, _31008_, _31007_);
  and _76639_ (_31010_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  and _76640_ (_31011_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or _76641_ (_31012_, _31011_, _31010_);
  or _76642_ (_31013_, _31012_, _31009_);
  and _76643_ (_31014_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  and _76644_ (_31015_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  nor _76645_ (_31016_, _31015_, _31014_);
  and _76646_ (_31017_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and _76647_ (_31018_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  nor _76648_ (_31019_, _31018_, _31017_);
  nand _76649_ (_31020_, _31019_, _31016_);
  or _76650_ (_31021_, _31020_, _31013_);
  and _76651_ (_31022_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and _76652_ (_31023_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  or _76653_ (_31024_, _31023_, _31022_);
  and _76654_ (_31025_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and _76655_ (_31026_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or _76656_ (_31027_, _31026_, _31025_);
  or _76657_ (_31028_, _31027_, _31024_);
  and _76658_ (_31029_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and _76659_ (_31030_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or _76660_ (_31031_, _31030_, _31029_);
  and _76661_ (_31032_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and _76662_ (_31033_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or _76663_ (_31034_, _31033_, _31032_);
  or _76664_ (_31035_, _31034_, _31031_);
  or _76665_ (_31036_, _31035_, _31028_);
  or _76666_ (_31037_, _31036_, _31021_);
  or _76667_ (_31038_, _31037_, _31006_);
  or _76668_ (_31039_, _31038_, _30975_);
  or _76669_ (_31040_, _31039_, _30912_);
  nor _76670_ (_31041_, _31040_, _30787_);
  and _76671_ (_31042_, _31041_, _30532_);
  and _76672_ (_31043_, _30010_, iram_op1_reg[5]);
  and _76673_ (_31044_, _31043_, iram_op1_reg[6]);
  nor _76674_ (_31045_, _31044_, iram_op1_reg[7]);
  and _76675_ (_31046_, _31044_, iram_op1_reg[7]);
  nor _76676_ (_31047_, _31046_, _31045_);
  nor _76677_ (_31048_, _31047_, _31042_);
  or _76678_ (_31049_, _31048_, _30530_);
  or _76679_ (_31050_, _31049_, _30015_);
  or _76680_ (_31051_, _31050_, _29496_);
  and _76681_ (_31052_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  not _76682_ (_31053_, _31052_);
  and _76683_ (_31054_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  and _76684_ (_31055_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  nor _76685_ (_31056_, _31055_, _31054_);
  and _76686_ (_31057_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and _76687_ (_31058_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  nor _76688_ (_31059_, _31058_, _31057_);
  and _76689_ (_31060_, _31059_, _31056_);
  and _76690_ (_31061_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  and _76691_ (_31062_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  nor _76692_ (_31063_, _31062_, _31061_);
  and _76693_ (_31064_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and _76694_ (_31065_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  nor _76695_ (_31066_, _31065_, _31064_);
  and _76696_ (_31067_, _31066_, _31063_);
  and _76697_ (_31068_, _31067_, _31060_);
  and _76698_ (_31069_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and _76699_ (_31070_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  nor _76700_ (_31071_, _31070_, _31069_);
  and _76701_ (_31072_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  and _76702_ (_31073_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  nor _76703_ (_31074_, _31073_, _31072_);
  and _76704_ (_31075_, _31074_, _31071_);
  and _76705_ (_31076_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and _76706_ (_31077_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  nor _76707_ (_31078_, _31077_, _31076_);
  and _76708_ (_31079_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  and _76709_ (_31080_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  nor _76710_ (_31081_, _31080_, _31079_);
  and _76711_ (_31082_, _31081_, _31078_);
  and _76712_ (_31083_, _31082_, _31075_);
  and _76713_ (_31084_, _31083_, _31068_);
  and _76714_ (_31085_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  and _76715_ (_31086_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  nor _76716_ (_31087_, _31086_, _31085_);
  and _76717_ (_31088_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and _76718_ (_31089_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  nor _76719_ (_31090_, _31089_, _31088_);
  and _76720_ (_31091_, _31090_, _31087_);
  and _76721_ (_31092_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  and _76722_ (_31093_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  nor _76723_ (_31094_, _31093_, _31092_);
  and _76724_ (_31095_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and _76725_ (_31096_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  nor _76726_ (_31097_, _31096_, _31095_);
  and _76727_ (_31098_, _31097_, _31094_);
  and _76728_ (_31099_, _31098_, _31091_);
  and _76729_ (_31100_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and _76730_ (_31101_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  nor _76731_ (_31102_, _31101_, _31100_);
  and _76732_ (_31103_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  and _76733_ (_31104_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  nor _76734_ (_31105_, _31104_, _31103_);
  and _76735_ (_31106_, _31105_, _31102_);
  and _76736_ (_31107_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and _76737_ (_31108_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  nor _76738_ (_31109_, _31108_, _31107_);
  and _76739_ (_31110_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  and _76740_ (_31111_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  nor _76741_ (_31112_, _31111_, _31110_);
  and _76742_ (_31113_, _31112_, _31109_);
  and _76743_ (_31114_, _31113_, _31106_);
  and _76744_ (_31115_, _31114_, _31099_);
  and _76745_ (_31116_, _31115_, _31084_);
  and _76746_ (_31117_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and _76747_ (_31118_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  nor _76748_ (_31119_, _31118_, _31117_);
  and _76749_ (_31120_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  and _76750_ (_31121_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  nor _76751_ (_31122_, _31121_, _31120_);
  and _76752_ (_31123_, _31122_, _31119_);
  and _76753_ (_31124_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and _76754_ (_31125_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  nor _76755_ (_31126_, _31125_, _31124_);
  and _76756_ (_31127_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  and _76757_ (_31128_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  nor _76758_ (_31129_, _31128_, _31127_);
  and _76759_ (_31130_, _31129_, _31126_);
  and _76760_ (_31131_, _31130_, _31123_);
  and _76761_ (_31132_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  and _76762_ (_31133_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  nor _76763_ (_31134_, _31133_, _31132_);
  and _76764_ (_31135_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and _76765_ (_31136_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  nor _76766_ (_31137_, _31136_, _31135_);
  and _76767_ (_31138_, _31137_, _31134_);
  and _76768_ (_31139_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  and _76769_ (_31140_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  nor _76770_ (_31141_, _31140_, _31139_);
  and _76771_ (_31142_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and _76772_ (_31143_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  nor _76773_ (_31144_, _31143_, _31142_);
  and _76774_ (_31145_, _31144_, _31141_);
  and _76775_ (_31146_, _31145_, _31138_);
  and _76776_ (_31147_, _31146_, _31131_);
  and _76777_ (_31148_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and _76778_ (_31149_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  nor _76779_ (_31150_, _31149_, _31148_);
  and _76780_ (_31151_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  and _76781_ (_31152_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  nor _76782_ (_31153_, _31152_, _31151_);
  and _76783_ (_31154_, _31153_, _31150_);
  and _76784_ (_31155_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  and _76785_ (_31156_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  nor _76786_ (_31157_, _31156_, _31155_);
  and _76787_ (_31158_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  and _76788_ (_31159_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  nor _76789_ (_31160_, _31159_, _31158_);
  and _76790_ (_31161_, _31160_, _31157_);
  and _76791_ (_31162_, _31161_, _31154_);
  and _76792_ (_31163_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and _76793_ (_31164_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  nor _76794_ (_31165_, _31164_, _31163_);
  and _76795_ (_31166_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  and _76796_ (_31167_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  nor _76797_ (_31168_, _31167_, _31166_);
  and _76798_ (_31169_, _31168_, _31165_);
  and _76799_ (_31170_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and _76800_ (_31171_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  nor _76801_ (_31172_, _31171_, _31170_);
  and _76802_ (_31173_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  and _76803_ (_31174_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  nor _76804_ (_31175_, _31174_, _31173_);
  and _76805_ (_31176_, _31175_, _31172_);
  and _76806_ (_31177_, _31176_, _31169_);
  and _76807_ (_31178_, _31177_, _31162_);
  and _76808_ (_31179_, _31178_, _31147_);
  and _76809_ (_31180_, _31179_, _31116_);
  and _76810_ (_31181_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and _76811_ (_31182_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  nor _76812_ (_31183_, _31182_, _31181_);
  and _76813_ (_31184_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  and _76814_ (_31185_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  nor _76815_ (_31186_, _31185_, _31184_);
  and _76816_ (_31187_, _31186_, _31183_);
  and _76817_ (_31188_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and _76818_ (_31189_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  nor _76819_ (_31190_, _31189_, _31188_);
  and _76820_ (_31191_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  and _76821_ (_31192_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  nor _76822_ (_31193_, _31192_, _31191_);
  and _76823_ (_31194_, _31193_, _31190_);
  and _76824_ (_31195_, _31194_, _31187_);
  and _76825_ (_31196_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  and _76826_ (_31197_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  nor _76827_ (_31198_, _31197_, _31196_);
  and _76828_ (_31199_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and _76829_ (_31200_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  nor _76830_ (_31201_, _31200_, _31199_);
  and _76831_ (_31202_, _31201_, _31198_);
  and _76832_ (_31203_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  and _76833_ (_31204_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  nor _76834_ (_31205_, _31204_, _31203_);
  and _76835_ (_31206_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and _76836_ (_31207_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  nor _76837_ (_31208_, _31207_, _31206_);
  and _76838_ (_31209_, _31208_, _31205_);
  and _76839_ (_31210_, _31209_, _31202_);
  and _76840_ (_31211_, _31210_, _31195_);
  and _76841_ (_31212_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  and _76842_ (_31213_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  nor _76843_ (_31214_, _31213_, _31212_);
  and _76844_ (_31215_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and _76845_ (_31216_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  nor _76846_ (_31217_, _31216_, _31215_);
  and _76847_ (_31218_, _31217_, _31214_);
  and _76848_ (_31219_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  and _76849_ (_31220_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  nor _76850_ (_31221_, _31220_, _31219_);
  and _76851_ (_31222_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and _76852_ (_31223_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  nor _76853_ (_31224_, _31223_, _31222_);
  and _76854_ (_31225_, _31224_, _31221_);
  and _76855_ (_31226_, _31225_, _31218_);
  and _76856_ (_31227_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and _76857_ (_31228_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  nor _76858_ (_31229_, _31228_, _31227_);
  and _76859_ (_31230_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  and _76860_ (_31231_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  nor _76861_ (_31232_, _31231_, _31230_);
  and _76862_ (_31233_, _31232_, _31229_);
  and _76863_ (_31234_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and _76864_ (_31235_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  nor _76865_ (_31236_, _31235_, _31234_);
  and _76866_ (_31237_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  and _76867_ (_31238_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  nor _76868_ (_31239_, _31238_, _31237_);
  and _76869_ (_31240_, _31239_, _31236_);
  and _76870_ (_31241_, _31240_, _31233_);
  and _76871_ (_31242_, _31241_, _31226_);
  and _76872_ (_31243_, _31242_, _31211_);
  and _76873_ (_31244_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and _76874_ (_31245_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  nor _76875_ (_31246_, _31245_, _31244_);
  and _76876_ (_31247_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  and _76877_ (_31248_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  nor _76878_ (_31249_, _31248_, _31247_);
  and _76879_ (_31250_, _31249_, _31246_);
  and _76880_ (_31251_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  and _76881_ (_31252_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  nor _76882_ (_31253_, _31252_, _31251_);
  and _76883_ (_31254_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and _76884_ (_31255_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  nor _76885_ (_31256_, _31255_, _31254_);
  and _76886_ (_31257_, _31256_, _31253_);
  and _76887_ (_31258_, _31257_, _31250_);
  and _76888_ (_31259_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and _76889_ (_31260_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  nor _76890_ (_31261_, _31260_, _31259_);
  and _76891_ (_31262_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  and _76892_ (_31263_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  nor _76893_ (_31264_, _31263_, _31262_);
  and _76894_ (_31265_, _31264_, _31261_);
  and _76895_ (_31266_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and _76896_ (_31267_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  nor _76897_ (_31268_, _31267_, _31266_);
  and _76898_ (_31269_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  and _76899_ (_31270_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  nor _76900_ (_31271_, _31270_, _31269_);
  and _76901_ (_31272_, _31271_, _31268_);
  and _76902_ (_31273_, _31272_, _31265_);
  and _76903_ (_31274_, _31273_, _31258_);
  and _76904_ (_31275_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and _76905_ (_31276_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  nor _76906_ (_31277_, _31276_, _31275_);
  and _76907_ (_31278_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  and _76908_ (_31279_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  nor _76909_ (_31280_, _31279_, _31278_);
  and _76910_ (_31281_, _31280_, _31277_);
  and _76911_ (_31282_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and _76912_ (_31283_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  nor _76913_ (_31284_, _31283_, _31282_);
  and _76914_ (_31285_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  and _76915_ (_31286_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  nor _76916_ (_31287_, _31286_, _31285_);
  and _76917_ (_31288_, _31287_, _31284_);
  and _76918_ (_31289_, _31288_, _31281_);
  and _76919_ (_31290_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  and _76920_ (_31291_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  nor _76921_ (_31292_, _31291_, _31290_);
  and _76922_ (_31293_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and _76923_ (_31294_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  nor _76924_ (_31295_, _31294_, _31293_);
  and _76925_ (_31296_, _31295_, _31292_);
  and _76926_ (_31297_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  and _76927_ (_31298_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  nor _76928_ (_31299_, _31298_, _31297_);
  and _76929_ (_31300_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  and _76930_ (_31301_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  nor _76931_ (_31302_, _31301_, _31300_);
  and _76932_ (_31303_, _31302_, _31299_);
  and _76933_ (_31304_, _31303_, _31296_);
  and _76934_ (_31305_, _31304_, _31289_);
  and _76935_ (_31306_, _31305_, _31274_);
  and _76936_ (_31307_, _31306_, _31243_);
  and _76937_ (_31308_, _31307_, _31180_);
  and _76938_ (_31309_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and _76939_ (_31310_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  nor _76940_ (_31311_, _31310_, _31309_);
  and _76941_ (_31312_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  and _76942_ (_31313_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  nor _76943_ (_31314_, _31313_, _31312_);
  and _76944_ (_31315_, _31314_, _31311_);
  and _76945_ (_31316_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and _76946_ (_31317_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  nor _76947_ (_31318_, _31317_, _31316_);
  and _76948_ (_31319_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  and _76949_ (_31320_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  nor _76950_ (_31321_, _31320_, _31319_);
  and _76951_ (_31322_, _31321_, _31318_);
  and _76952_ (_31323_, _31322_, _31315_);
  and _76953_ (_31324_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  and _76954_ (_31325_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  nor _76955_ (_31326_, _31325_, _31324_);
  and _76956_ (_31327_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and _76957_ (_31328_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  nor _76958_ (_31329_, _31328_, _31327_);
  and _76959_ (_31330_, _31329_, _31326_);
  and _76960_ (_31331_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  and _76961_ (_31332_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  nor _76962_ (_31333_, _31332_, _31331_);
  and _76963_ (_31334_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and _76964_ (_31335_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  nor _76965_ (_31336_, _31335_, _31334_);
  and _76966_ (_31337_, _31336_, _31333_);
  and _76967_ (_31338_, _31337_, _31330_);
  and _76968_ (_31339_, _31338_, _31323_);
  and _76969_ (_31340_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  and _76970_ (_31341_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  nor _76971_ (_31342_, _31341_, _31340_);
  and _76972_ (_31343_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and _76973_ (_31344_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  nor _76974_ (_31345_, _31344_, _31343_);
  and _76975_ (_31346_, _31345_, _31342_);
  and _76976_ (_31347_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  and _76977_ (_31348_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  nor _76978_ (_31349_, _31348_, _31347_);
  and _76979_ (_31350_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  and _76980_ (_31351_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  nor _76981_ (_31352_, _31351_, _31350_);
  and _76982_ (_31353_, _31352_, _31349_);
  and _76983_ (_31354_, _31353_, _31346_);
  and _76984_ (_31355_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and _76985_ (_31356_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  nor _76986_ (_31357_, _31356_, _31355_);
  and _76987_ (_31358_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  and _76988_ (_31359_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  nor _76989_ (_31360_, _31359_, _31358_);
  and _76990_ (_31361_, _31360_, _31357_);
  and _76991_ (_31362_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and _76992_ (_31363_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  nor _76993_ (_31364_, _31363_, _31362_);
  and _76994_ (_31365_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  and _76995_ (_31366_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  nor _76996_ (_31367_, _31366_, _31365_);
  and _76997_ (_31368_, _31367_, _31364_);
  and _76998_ (_31369_, _31368_, _31361_);
  and _76999_ (_31370_, _31369_, _31354_);
  and _77000_ (_31371_, _31370_, _31339_);
  and _77001_ (_31372_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and _77002_ (_31373_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  nor _77003_ (_31374_, _31373_, _31372_);
  and _77004_ (_31375_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  and _77005_ (_31376_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  nor _77006_ (_31377_, _31376_, _31375_);
  and _77007_ (_31378_, _31377_, _31374_);
  and _77008_ (_31379_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  and _77009_ (_31380_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  nor _77010_ (_31381_, _31380_, _31379_);
  and _77011_ (_31382_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and _77012_ (_31383_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  nor _77013_ (_31384_, _31383_, _31382_);
  and _77014_ (_31385_, _31384_, _31381_);
  and _77015_ (_31386_, _31385_, _31378_);
  and _77016_ (_31387_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and _77017_ (_31388_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  nor _77018_ (_31389_, _31388_, _31387_);
  and _77019_ (_31390_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  and _77020_ (_31391_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  nor _77021_ (_31392_, _31391_, _31390_);
  and _77022_ (_31393_, _31392_, _31389_);
  and _77023_ (_31394_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and _77024_ (_31395_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  nor _77025_ (_31396_, _31395_, _31394_);
  and _77026_ (_31397_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  and _77027_ (_31398_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  nor _77028_ (_31399_, _31398_, _31397_);
  and _77029_ (_31400_, _31399_, _31396_);
  and _77030_ (_31401_, _31400_, _31393_);
  and _77031_ (_31402_, _31401_, _31386_);
  and _77032_ (_31403_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and _77033_ (_31404_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  nor _77034_ (_31405_, _31404_, _31403_);
  and _77035_ (_31406_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  and _77036_ (_31407_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  nor _77037_ (_31408_, _31407_, _31406_);
  and _77038_ (_31409_, _31408_, _31405_);
  and _77039_ (_31410_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  and _77040_ (_31411_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  nor _77041_ (_31412_, _31411_, _31410_);
  and _77042_ (_31413_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  and _77043_ (_31414_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  nor _77044_ (_31415_, _31414_, _31413_);
  and _77045_ (_31416_, _31415_, _31412_);
  and _77046_ (_31417_, _31416_, _31409_);
  and _77047_ (_31418_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  and _77048_ (_31419_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  nor _77049_ (_31420_, _31419_, _31418_);
  and _77050_ (_31421_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and _77051_ (_31422_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  nor _77052_ (_31423_, _31422_, _31421_);
  and _77053_ (_31424_, _31423_, _31420_);
  and _77054_ (_31425_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  and _77055_ (_31426_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  nor _77056_ (_31427_, _31426_, _31425_);
  and _77057_ (_31428_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  and _77058_ (_31429_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  nor _77059_ (_31430_, _31429_, _31428_);
  and _77060_ (_31431_, _31430_, _31427_);
  and _77061_ (_31432_, _31431_, _31424_);
  and _77062_ (_31433_, _31432_, _31417_);
  and _77063_ (_31434_, _31433_, _31402_);
  and _77064_ (_31435_, _31434_, _31371_);
  and _77065_ (_31436_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and _77066_ (_31437_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  nor _77067_ (_31438_, _31437_, _31436_);
  and _77068_ (_31439_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  and _77069_ (_31440_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  nor _77070_ (_31441_, _31440_, _31439_);
  and _77071_ (_31442_, _31441_, _31438_);
  and _77072_ (_31443_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and _77073_ (_31444_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  nor _77074_ (_31445_, _31444_, _31443_);
  and _77075_ (_31446_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  and _77076_ (_31447_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  nor _77077_ (_31448_, _31447_, _31446_);
  and _77078_ (_31449_, _31448_, _31445_);
  and _77079_ (_31450_, _31449_, _31442_);
  and _77080_ (_31451_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  and _77081_ (_31452_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  nor _77082_ (_31453_, _31452_, _31451_);
  and _77083_ (_31454_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and _77084_ (_31455_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  nor _77085_ (_31456_, _31455_, _31454_);
  and _77086_ (_31457_, _31456_, _31453_);
  and _77087_ (_31458_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  and _77088_ (_31459_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  nor _77089_ (_31460_, _31459_, _31458_);
  and _77090_ (_31461_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and _77091_ (_31462_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  nor _77092_ (_31463_, _31462_, _31461_);
  and _77093_ (_31464_, _31463_, _31460_);
  and _77094_ (_31465_, _31464_, _31457_);
  and _77095_ (_31466_, _31465_, _31450_);
  and _77096_ (_31467_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  and _77097_ (_31468_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  nor _77098_ (_31469_, _31468_, _31467_);
  and _77099_ (_31470_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and _77100_ (_31471_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  nor _77101_ (_31472_, _31471_, _31470_);
  and _77102_ (_31473_, _31472_, _31469_);
  and _77103_ (_31474_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  and _77104_ (_31475_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  nor _77105_ (_31476_, _31475_, _31474_);
  and _77106_ (_31477_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and _77107_ (_31478_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  nor _77108_ (_31479_, _31478_, _31477_);
  and _77109_ (_31480_, _31479_, _31476_);
  and _77110_ (_31481_, _31480_, _31473_);
  and _77111_ (_31482_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and _77112_ (_31483_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  nor _77113_ (_31484_, _31483_, _31482_);
  and _77114_ (_31485_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  and _77115_ (_31486_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  nor _77116_ (_31487_, _31486_, _31485_);
  and _77117_ (_31488_, _31487_, _31484_);
  and _77118_ (_31489_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and _77119_ (_31490_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  nor _77120_ (_31491_, _31490_, _31489_);
  and _77121_ (_31492_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  and _77122_ (_31493_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  nor _77123_ (_31494_, _31493_, _31492_);
  and _77124_ (_31495_, _31494_, _31491_);
  and _77125_ (_31496_, _31495_, _31488_);
  and _77126_ (_31497_, _31496_, _31481_);
  and _77127_ (_31498_, _31497_, _31466_);
  and _77128_ (_31499_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  and _77129_ (_31500_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  nor _77130_ (_31501_, _31500_, _31499_);
  and _77131_ (_31502_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and _77132_ (_31503_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  nor _77133_ (_31504_, _31503_, _31502_);
  and _77134_ (_31505_, _31504_, _31501_);
  and _77135_ (_31506_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and _77136_ (_31507_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  nor _77137_ (_31508_, _31507_, _31506_);
  and _77138_ (_31509_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and _77139_ (_31510_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  nor _77140_ (_31511_, _31510_, _31509_);
  and _77141_ (_31512_, _31511_, _31508_);
  and _77142_ (_31513_, _31512_, _31505_);
  and _77143_ (_31514_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  and _77144_ (_31515_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  nor _77145_ (_31516_, _31515_, _31514_);
  and _77146_ (_31517_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and _77147_ (_31518_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  nor _77148_ (_31519_, _31518_, _31517_);
  and _77149_ (_31520_, _31519_, _31516_);
  and _77150_ (_31521_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  and _77151_ (_31522_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  nor _77152_ (_31523_, _31522_, _31521_);
  and _77153_ (_31524_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and _77154_ (_31525_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  nor _77155_ (_31526_, _31525_, _31524_);
  and _77156_ (_31527_, _31526_, _31523_);
  and _77157_ (_31528_, _31527_, _31520_);
  and _77158_ (_31529_, _31528_, _31513_);
  and _77159_ (_31530_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and _77160_ (_31531_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor _77161_ (_31532_, _31531_, _31530_);
  and _77162_ (_31533_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and _77163_ (_31534_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor _77164_ (_31535_, _31534_, _31533_);
  and _77165_ (_31536_, _31535_, _31532_);
  and _77166_ (_31537_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and _77167_ (_31538_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and _77168_ (_31539_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _77169_ (_31540_, _31539_, _31538_);
  nor _77170_ (_31541_, _31540_, _31537_);
  and _77171_ (_31542_, _31541_, _31536_);
  and _77172_ (_31543_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _77173_ (_31544_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor _77174_ (_31545_, _31544_, _31543_);
  and _77175_ (_31546_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and _77176_ (_31547_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor _77177_ (_31548_, _31547_, _31546_);
  and _77178_ (_31549_, _31548_, _31545_);
  and _77179_ (_31550_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and _77180_ (_31551_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor _77181_ (_31552_, _31551_, _31550_);
  and _77182_ (_31553_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and _77183_ (_31554_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor _77184_ (_31555_, _31554_, _31553_);
  and _77185_ (_31556_, _31555_, _31552_);
  and _77186_ (_31557_, _31556_, _31549_);
  and _77187_ (_31558_, _31557_, _31542_);
  and _77188_ (_31559_, _31558_, _31529_);
  and _77189_ (_31560_, _31559_, _31498_);
  and _77190_ (_31561_, _31560_, _31435_);
  and _77191_ (_31562_, _31561_, _31308_);
  and _77192_ (_31563_, _31562_, _31053_);
  nor _77193_ (_31564_, _31563_, _21566_);
  and _77194_ (_31565_, _31563_, _21566_);
  or _77195_ (_31566_, _31565_, _31564_);
  and _77196_ (_31567_, _31566_, iram_op1_reg[0]);
  and _77197_ (_31568_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  not _77198_ (_31569_, _31568_);
  and _77199_ (_31570_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  and _77200_ (_31571_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  nor _77201_ (_31572_, _31571_, _31570_);
  and _77202_ (_31573_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and _77203_ (_31574_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  nor _77204_ (_31575_, _31574_, _31573_);
  and _77205_ (_31576_, _31575_, _31572_);
  and _77206_ (_31577_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and _77207_ (_31578_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  nor _77208_ (_31579_, _31578_, _31577_);
  and _77209_ (_31580_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and _77210_ (_31581_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  nor _77211_ (_31582_, _31581_, _31580_);
  and _77212_ (_31583_, _31582_, _31579_);
  and _77213_ (_31584_, _31583_, _31576_);
  and _77214_ (_31585_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and _77215_ (_31586_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  nor _77216_ (_31587_, _31586_, _31585_);
  and _77217_ (_31588_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  and _77218_ (_31589_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  nor _77219_ (_31590_, _31589_, _31588_);
  and _77220_ (_31591_, _31590_, _31587_);
  and _77221_ (_31592_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  and _77222_ (_31593_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  nor _77223_ (_31594_, _31593_, _31592_);
  and _77224_ (_31595_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and _77225_ (_31596_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  nor _77226_ (_31597_, _31596_, _31595_);
  and _77227_ (_31598_, _31597_, _31594_);
  and _77228_ (_31599_, _31598_, _31591_);
  and _77229_ (_31600_, _31599_, _31584_);
  and _77230_ (_31601_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  and _77231_ (_31602_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  nor _77232_ (_31603_, _31602_, _31601_);
  and _77233_ (_31604_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and _77234_ (_31605_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  nor _77235_ (_31606_, _31605_, _31604_);
  and _77236_ (_31607_, _31606_, _31603_);
  and _77237_ (_31608_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and _77238_ (_31609_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  nor _77239_ (_31610_, _31609_, _31608_);
  and _77240_ (_31611_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  and _77241_ (_31612_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  nor _77242_ (_31613_, _31612_, _31611_);
  and _77243_ (_31614_, _31613_, _31610_);
  and _77244_ (_31615_, _31614_, _31607_);
  and _77245_ (_31616_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  and _77246_ (_31617_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  nor _77247_ (_31618_, _31617_, _31616_);
  and _77248_ (_31619_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  and _77249_ (_31620_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  nor _77250_ (_31621_, _31620_, _31619_);
  and _77251_ (_31622_, _31621_, _31618_);
  and _77252_ (_31623_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  and _77253_ (_31624_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  nor _77254_ (_31625_, _31624_, _31623_);
  and _77255_ (_31626_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and _77256_ (_31627_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  nor _77257_ (_31628_, _31627_, _31626_);
  and _77258_ (_31629_, _31628_, _31625_);
  and _77259_ (_31630_, _31629_, _31622_);
  and _77260_ (_31631_, _31630_, _31615_);
  and _77261_ (_31632_, _31631_, _31600_);
  and _77262_ (_31633_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and _77263_ (_31634_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  nor _77264_ (_31635_, _31634_, _31633_);
  and _77265_ (_31636_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  and _77266_ (_31637_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  nor _77267_ (_31638_, _31637_, _31636_);
  and _77268_ (_31639_, _31638_, _31635_);
  and _77269_ (_31640_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and _77270_ (_31641_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  nor _77271_ (_31642_, _31641_, _31640_);
  and _77272_ (_31643_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  and _77273_ (_31644_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  nor _77274_ (_31645_, _31644_, _31643_);
  and _77275_ (_31646_, _31645_, _31642_);
  and _77276_ (_31647_, _31646_, _31639_);
  and _77277_ (_31648_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  and _77278_ (_31649_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  nor _77279_ (_31650_, _31649_, _31648_);
  and _77280_ (_31651_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and _77281_ (_31652_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  nor _77282_ (_31653_, _31652_, _31651_);
  and _77283_ (_31654_, _31653_, _31650_);
  and _77284_ (_31655_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  and _77285_ (_31656_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  nor _77286_ (_31657_, _31656_, _31655_);
  and _77287_ (_31658_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and _77288_ (_31659_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  nor _77289_ (_31660_, _31659_, _31658_);
  and _77290_ (_31661_, _31660_, _31657_);
  and _77291_ (_31662_, _31661_, _31654_);
  and _77292_ (_31663_, _31662_, _31647_);
  and _77293_ (_31664_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and _77294_ (_31665_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  nor _77295_ (_31666_, _31665_, _31664_);
  and _77296_ (_31667_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  and _77297_ (_31668_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  nor _77298_ (_31669_, _31668_, _31667_);
  and _77299_ (_31670_, _31669_, _31666_);
  and _77300_ (_31671_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  and _77301_ (_31672_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  nor _77302_ (_31673_, _31672_, _31671_);
  and _77303_ (_31674_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  and _77304_ (_31675_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  nor _77305_ (_31676_, _31675_, _31674_);
  and _77306_ (_31677_, _31676_, _31673_);
  and _77307_ (_31678_, _31677_, _31670_);
  and _77308_ (_31679_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  and _77309_ (_31680_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  nor _77310_ (_31681_, _31680_, _31679_);
  and _77311_ (_31682_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and _77312_ (_31683_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  nor _77313_ (_31684_, _31683_, _31682_);
  and _77314_ (_31685_, _31684_, _31681_);
  and _77315_ (_31686_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  and _77316_ (_31687_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  nor _77317_ (_31688_, _31687_, _31686_);
  and _77318_ (_31689_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  and _77319_ (_31690_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  nor _77320_ (_31691_, _31690_, _31689_);
  and _77321_ (_31692_, _31691_, _31688_);
  and _77322_ (_31693_, _31692_, _31685_);
  and _77323_ (_31694_, _31693_, _31678_);
  and _77324_ (_31695_, _31694_, _31663_);
  and _77325_ (_31696_, _31695_, _31632_);
  and _77326_ (_31697_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  and _77327_ (_31698_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  nor _77328_ (_31699_, _31698_, _31697_);
  and _77329_ (_31700_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and _77330_ (_31701_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  nor _77331_ (_31702_, _31701_, _31700_);
  and _77332_ (_31703_, _31702_, _31699_);
  and _77333_ (_31704_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and _77334_ (_31705_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  nor _77335_ (_31706_, _31705_, _31704_);
  and _77336_ (_31707_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  and _77337_ (_31708_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  nor _77338_ (_31709_, _31708_, _31707_);
  and _77339_ (_31710_, _31709_, _31706_);
  and _77340_ (_31711_, _31710_, _31703_);
  and _77341_ (_31712_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and _77342_ (_31713_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  nor _77343_ (_31714_, _31713_, _31712_);
  and _77344_ (_31715_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  and _77345_ (_31716_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  nor _77346_ (_31717_, _31716_, _31715_);
  and _77347_ (_31718_, _31717_, _31714_);
  and _77348_ (_31719_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and _77349_ (_31720_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  nor _77350_ (_31721_, _31720_, _31719_);
  and _77351_ (_31722_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and _77352_ (_31723_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  nor _77353_ (_31724_, _31723_, _31722_);
  and _77354_ (_31725_, _31724_, _31721_);
  and _77355_ (_31726_, _31725_, _31718_);
  and _77356_ (_31727_, _31726_, _31711_);
  and _77357_ (_31728_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and _77358_ (_31729_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  nor _77359_ (_31730_, _31729_, _31728_);
  and _77360_ (_31731_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  and _77361_ (_31732_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  nor _77362_ (_31733_, _31732_, _31731_);
  and _77363_ (_31734_, _31733_, _31730_);
  and _77364_ (_31735_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and _77365_ (_31736_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  nor _77366_ (_31737_, _31736_, _31735_);
  and _77367_ (_31738_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and _77368_ (_31739_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  nor _77369_ (_31740_, _31739_, _31738_);
  and _77370_ (_31741_, _31740_, _31737_);
  and _77371_ (_31742_, _31741_, _31734_);
  and _77372_ (_31743_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  and _77373_ (_31744_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  nor _77374_ (_31745_, _31744_, _31743_);
  and _77375_ (_31746_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and _77376_ (_31747_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  nor _77377_ (_31748_, _31747_, _31746_);
  and _77378_ (_31749_, _31748_, _31745_);
  and _77379_ (_31750_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and _77380_ (_31751_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  nor _77381_ (_31752_, _31751_, _31750_);
  and _77382_ (_31753_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  and _77383_ (_31754_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  nor _77384_ (_31755_, _31754_, _31753_);
  and _77385_ (_31756_, _31755_, _31752_);
  and _77386_ (_31757_, _31756_, _31749_);
  and _77387_ (_31758_, _31757_, _31742_);
  and _77388_ (_31759_, _31758_, _31727_);
  and _77389_ (_31760_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and _77390_ (_31761_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  nor _77391_ (_31762_, _31761_, _31760_);
  and _77392_ (_31763_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  and _77393_ (_31764_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  nor _77394_ (_31765_, _31764_, _31763_);
  and _77395_ (_31766_, _31765_, _31762_);
  and _77396_ (_31767_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and _77397_ (_31768_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  nor _77398_ (_31769_, _31768_, _31767_);
  and _77399_ (_31770_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  and _77400_ (_31771_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  nor _77401_ (_31772_, _31771_, _31770_);
  and _77402_ (_31773_, _31772_, _31769_);
  and _77403_ (_31774_, _31773_, _31766_);
  and _77404_ (_31775_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  and _77405_ (_31776_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  nor _77406_ (_31777_, _31776_, _31775_);
  and _77407_ (_31778_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and _77408_ (_31779_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  nor _77409_ (_31780_, _31779_, _31778_);
  and _77410_ (_31781_, _31780_, _31777_);
  and _77411_ (_31782_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  and _77412_ (_31783_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  nor _77413_ (_31784_, _31783_, _31782_);
  and _77414_ (_31785_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and _77415_ (_31786_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  nor _77416_ (_31787_, _31786_, _31785_);
  and _77417_ (_31788_, _31787_, _31784_);
  and _77418_ (_31789_, _31788_, _31781_);
  and _77419_ (_31790_, _31789_, _31774_);
  and _77420_ (_31791_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  and _77421_ (_31792_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  nor _77422_ (_31793_, _31792_, _31791_);
  and _77423_ (_31794_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and _77424_ (_31795_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  nor _77425_ (_31796_, _31795_, _31794_);
  and _77426_ (_31797_, _31796_, _31793_);
  and _77427_ (_31798_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  and _77428_ (_31799_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  nor _77429_ (_31800_, _31799_, _31798_);
  and _77430_ (_31801_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  and _77431_ (_31802_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  nor _77432_ (_31803_, _31802_, _31801_);
  and _77433_ (_31804_, _31803_, _31800_);
  and _77434_ (_31805_, _31804_, _31797_);
  and _77435_ (_31806_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and _77436_ (_31807_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  nor _77437_ (_31808_, _31807_, _31806_);
  and _77438_ (_31809_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  and _77439_ (_31810_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  nor _77440_ (_31811_, _31810_, _31809_);
  and _77441_ (_31812_, _31811_, _31808_);
  and _77442_ (_31813_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  and _77443_ (_31814_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  nor _77444_ (_31815_, _31814_, _31813_);
  and _77445_ (_31816_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and _77446_ (_31817_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  nor _77447_ (_31818_, _31817_, _31816_);
  and _77448_ (_31819_, _31818_, _31815_);
  and _77449_ (_31820_, _31819_, _31812_);
  and _77450_ (_31821_, _31820_, _31805_);
  and _77451_ (_31822_, _31821_, _31790_);
  and _77452_ (_31823_, _31822_, _31759_);
  and _77453_ (_31824_, _31823_, _31696_);
  and _77454_ (_31825_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and _77455_ (_31826_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  nor _77456_ (_31827_, _31826_, _31825_);
  and _77457_ (_31828_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and _77458_ (_31829_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  nor _77459_ (_31830_, _31829_, _31828_);
  and _77460_ (_31831_, _31830_, _31827_);
  and _77461_ (_31832_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and _77462_ (_31833_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  nor _77463_ (_31834_, _31833_, _31832_);
  and _77464_ (_31835_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  and _77465_ (_31836_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  nor _77466_ (_31837_, _31836_, _31835_);
  and _77467_ (_31838_, _31837_, _31834_);
  and _77468_ (_31839_, _31838_, _31831_);
  and _77469_ (_31840_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  and _77470_ (_31841_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  nor _77471_ (_31842_, _31841_, _31840_);
  and _77472_ (_31843_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and _77473_ (_31844_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  nor _77474_ (_31845_, _31844_, _31843_);
  and _77475_ (_31846_, _31845_, _31842_);
  and _77476_ (_31847_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and _77477_ (_31848_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  nor _77478_ (_31849_, _31848_, _31847_);
  and _77479_ (_31850_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  and _77480_ (_31851_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  nor _77481_ (_31852_, _31851_, _31850_);
  and _77482_ (_31853_, _31852_, _31849_);
  and _77483_ (_31854_, _31853_, _31846_);
  and _77484_ (_31855_, _31854_, _31839_);
  and _77485_ (_31856_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  and _77486_ (_31857_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  nor _77487_ (_31858_, _31857_, _31856_);
  and _77488_ (_31859_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and _77489_ (_31860_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  nor _77490_ (_31861_, _31860_, _31859_);
  and _77491_ (_31862_, _31861_, _31858_);
  and _77492_ (_31863_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and _77493_ (_31864_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  nor _77494_ (_31865_, _31864_, _31863_);
  and _77495_ (_31866_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  and _77496_ (_31867_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  nor _77497_ (_31868_, _31867_, _31866_);
  and _77498_ (_31869_, _31868_, _31865_);
  and _77499_ (_31870_, _31869_, _31862_);
  and _77500_ (_31871_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  and _77501_ (_31872_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  nor _77502_ (_31873_, _31872_, _31871_);
  and _77503_ (_31874_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and _77504_ (_31875_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  nor _77505_ (_31876_, _31875_, _31874_);
  and _77506_ (_31877_, _31876_, _31873_);
  and _77507_ (_31878_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and _77508_ (_31879_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  nor _77509_ (_31880_, _31879_, _31878_);
  and _77510_ (_31881_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  and _77511_ (_31882_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  nor _77512_ (_31883_, _31882_, _31881_);
  and _77513_ (_31884_, _31883_, _31880_);
  and _77514_ (_31885_, _31884_, _31877_);
  and _77515_ (_31886_, _31885_, _31870_);
  and _77516_ (_31887_, _31886_, _31855_);
  and _77517_ (_31888_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  and _77518_ (_31889_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  nor _77519_ (_31890_, _31889_, _31888_);
  and _77520_ (_31891_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and _77521_ (_31892_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  nor _77522_ (_31893_, _31892_, _31891_);
  and _77523_ (_31894_, _31893_, _31890_);
  and _77524_ (_31895_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  and _77525_ (_31896_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  nor _77526_ (_31897_, _31896_, _31895_);
  and _77527_ (_31898_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and _77528_ (_31899_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  nor _77529_ (_31900_, _31899_, _31898_);
  and _77530_ (_31901_, _31900_, _31897_);
  and _77531_ (_31902_, _31901_, _31894_);
  and _77532_ (_31903_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and _77533_ (_31904_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  nor _77534_ (_31905_, _31904_, _31903_);
  and _77535_ (_31906_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  and _77536_ (_31907_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  nor _77537_ (_31908_, _31907_, _31906_);
  and _77538_ (_31909_, _31908_, _31905_);
  and _77539_ (_31910_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and _77540_ (_31911_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  nor _77541_ (_31912_, _31911_, _31910_);
  and _77542_ (_31913_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  and _77543_ (_31914_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  nor _77544_ (_31915_, _31914_, _31913_);
  and _77545_ (_31916_, _31915_, _31912_);
  and _77546_ (_31917_, _31916_, _31909_);
  and _77547_ (_31918_, _31917_, _31902_);
  and _77548_ (_31919_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  and _77549_ (_31920_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  nor _77550_ (_31921_, _31920_, _31919_);
  and _77551_ (_31922_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and _77552_ (_31923_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  nor _77553_ (_31924_, _31923_, _31922_);
  and _77554_ (_31925_, _31924_, _31921_);
  and _77555_ (_31926_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  and _77556_ (_31927_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  nor _77557_ (_31928_, _31927_, _31926_);
  and _77558_ (_31929_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  and _77559_ (_31930_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  nor _77560_ (_31931_, _31930_, _31929_);
  and _77561_ (_31932_, _31931_, _31928_);
  and _77562_ (_31933_, _31932_, _31925_);
  and _77563_ (_31934_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and _77564_ (_31935_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  nor _77565_ (_31936_, _31935_, _31934_);
  and _77566_ (_31937_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  and _77567_ (_31938_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  nor _77568_ (_31939_, _31938_, _31937_);
  and _77569_ (_31940_, _31939_, _31936_);
  and _77570_ (_31941_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and _77571_ (_31942_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  nor _77572_ (_31943_, _31942_, _31941_);
  and _77573_ (_31944_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  and _77574_ (_31945_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  nor _77575_ (_31946_, _31945_, _31944_);
  and _77576_ (_31947_, _31946_, _31943_);
  and _77577_ (_31948_, _31947_, _31940_);
  and _77578_ (_31949_, _31948_, _31933_);
  and _77579_ (_31950_, _31949_, _31918_);
  and _77580_ (_31951_, _31950_, _31887_);
  and _77581_ (_31952_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  and _77582_ (_31953_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  nor _77583_ (_31954_, _31953_, _31952_);
  and _77584_ (_31955_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and _77585_ (_31956_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  nor _77586_ (_31957_, _31956_, _31955_);
  and _77587_ (_31958_, _31957_, _31954_);
  and _77588_ (_31959_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  and _77589_ (_31960_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  nor _77590_ (_31961_, _31960_, _31959_);
  and _77591_ (_31962_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and _77592_ (_31963_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  nor _77593_ (_31964_, _31963_, _31962_);
  and _77594_ (_31965_, _31964_, _31961_);
  and _77595_ (_31966_, _31965_, _31958_);
  and _77596_ (_31967_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and _77597_ (_31968_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  nor _77598_ (_31969_, _31968_, _31967_);
  and _77599_ (_31970_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and _77600_ (_31971_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  nor _77601_ (_31972_, _31971_, _31970_);
  and _77602_ (_31973_, _31972_, _31969_);
  and _77603_ (_31974_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and _77604_ (_31975_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  nor _77605_ (_31976_, _31975_, _31974_);
  and _77606_ (_31977_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  and _77607_ (_31978_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  nor _77608_ (_31979_, _31978_, _31977_);
  and _77609_ (_31980_, _31979_, _31976_);
  and _77610_ (_31981_, _31980_, _31973_);
  and _77611_ (_31982_, _31981_, _31966_);
  and _77612_ (_31983_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  and _77613_ (_31984_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  nor _77614_ (_31985_, _31984_, _31983_);
  and _77615_ (_31986_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and _77616_ (_31987_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  nor _77617_ (_31988_, _31987_, _31986_);
  and _77618_ (_31989_, _31988_, _31985_);
  and _77619_ (_31990_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  and _77620_ (_31991_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  nor _77621_ (_31992_, _31991_, _31990_);
  and _77622_ (_31993_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and _77623_ (_31994_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  nor _77624_ (_31995_, _31994_, _31993_);
  and _77625_ (_31996_, _31995_, _31992_);
  and _77626_ (_31997_, _31996_, _31989_);
  and _77627_ (_31998_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and _77628_ (_31999_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  nor _77629_ (_32000_, _31999_, _31998_);
  and _77630_ (_32001_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  and _77631_ (_32002_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  nor _77632_ (_32003_, _32002_, _32001_);
  and _77633_ (_32004_, _32003_, _32000_);
  and _77634_ (_32005_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and _77635_ (_32006_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  nor _77636_ (_32007_, _32006_, _32005_);
  and _77637_ (_32008_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  and _77638_ (_32009_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  nor _77639_ (_32010_, _32009_, _32008_);
  and _77640_ (_32011_, _32010_, _32007_);
  and _77641_ (_32012_, _32011_, _32004_);
  and _77642_ (_32013_, _32012_, _31997_);
  and _77643_ (_32014_, _32013_, _31982_);
  and _77644_ (_32015_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  and _77645_ (_32016_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  nor _77646_ (_32017_, _32016_, _32015_);
  and _77647_ (_32018_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and _77648_ (_32019_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  nor _77649_ (_32020_, _32019_, _32018_);
  and _77650_ (_32021_, _32020_, _32017_);
  and _77651_ (_32022_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  and _77652_ (_32023_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  nor _77653_ (_32024_, _32023_, _32022_);
  and _77654_ (_32025_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and _77655_ (_32026_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  nor _77656_ (_32027_, _32026_, _32025_);
  and _77657_ (_32028_, _32027_, _32024_);
  and _77658_ (_32029_, _32028_, _32021_);
  and _77659_ (_32030_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and _77660_ (_32031_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  nor _77661_ (_32032_, _32031_, _32030_);
  and _77662_ (_32033_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  and _77663_ (_32034_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  nor _77664_ (_32035_, _32034_, _32033_);
  and _77665_ (_32036_, _32035_, _32032_);
  and _77666_ (_32037_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and _77667_ (_32038_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  nor _77668_ (_32039_, _32038_, _32037_);
  and _77669_ (_32040_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  and _77670_ (_32041_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  nor _77671_ (_32042_, _32041_, _32040_);
  and _77672_ (_32043_, _32042_, _32039_);
  and _77673_ (_32044_, _32043_, _32036_);
  and _77674_ (_32045_, _32044_, _32029_);
  and _77675_ (_32046_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and _77676_ (_32047_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor _77677_ (_32048_, _32047_, _32046_);
  and _77678_ (_32049_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and _77679_ (_32050_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor _77680_ (_32051_, _32050_, _32049_);
  and _77681_ (_32052_, _32051_, _32048_);
  and _77682_ (_32053_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and _77683_ (_32054_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and _77684_ (_32055_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or _77685_ (_32056_, _32055_, _32054_);
  nor _77686_ (_32057_, _32056_, _32053_);
  and _77687_ (_32058_, _32057_, _32052_);
  and _77688_ (_32059_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and _77689_ (_32060_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor _77690_ (_32061_, _32060_, _32059_);
  and _77691_ (_32062_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and _77692_ (_32063_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor _77693_ (_32064_, _32063_, _32062_);
  and _77694_ (_32065_, _32064_, _32061_);
  and _77695_ (_32066_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and _77696_ (_32067_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor _77697_ (_32068_, _32067_, _32066_);
  and _77698_ (_32069_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and _77699_ (_32070_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor _77700_ (_32071_, _32070_, _32069_);
  and _77701_ (_32072_, _32071_, _32068_);
  and _77702_ (_32073_, _32072_, _32065_);
  and _77703_ (_32074_, _32073_, _32058_);
  and _77704_ (_32075_, _32074_, _32045_);
  and _77705_ (_32076_, _32075_, _32014_);
  and _77706_ (_32077_, _32076_, _31951_);
  and _77707_ (_32078_, _32077_, _31824_);
  and _77708_ (_32079_, _32078_, _31569_);
  nor _77709_ (_32080_, _32079_, _31566_);
  or _77710_ (_32081_, _32080_, _31567_);
  nor _77711_ (_32082_, _30529_, _30527_);
  and _77712_ (_32083_, _32079_, _21570_);
  and _77713_ (_32084_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  not _77714_ (_32085_, _32084_);
  and _77715_ (_32086_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  and _77716_ (_32087_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or _77717_ (_32088_, _32087_, _32086_);
  and _77718_ (_32089_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and _77719_ (_32090_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  or _77720_ (_32091_, _32090_, _32089_);
  or _77721_ (_32092_, _32091_, _32088_);
  and _77722_ (_32093_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  and _77723_ (_32094_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or _77724_ (_32095_, _32094_, _32093_);
  and _77725_ (_32096_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and _77726_ (_32097_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or _77727_ (_32098_, _32097_, _32096_);
  or _77728_ (_32099_, _32098_, _32095_);
  or _77729_ (_32100_, _32099_, _32092_);
  and _77730_ (_32101_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  and _77731_ (_32102_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or _77732_ (_32103_, _32102_, _32101_);
  and _77733_ (_32104_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  and _77734_ (_32105_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or _77735_ (_32106_, _32105_, _32104_);
  or _77736_ (_32107_, _32106_, _32103_);
  and _77737_ (_32108_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and _77738_ (_32109_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or _77739_ (_32110_, _32109_, _32108_);
  and _77740_ (_32111_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  and _77741_ (_32112_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or _77742_ (_32113_, _32112_, _32111_);
  or _77743_ (_32114_, _32113_, _32110_);
  or _77744_ (_32115_, _32114_, _32107_);
  or _77745_ (_32116_, _32115_, _32100_);
  and _77746_ (_32117_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  and _77747_ (_32118_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or _77748_ (_32119_, _32118_, _32117_);
  and _77749_ (_32120_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  and _77750_ (_32121_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or _77751_ (_32122_, _32121_, _32120_);
  or _77752_ (_32123_, _32122_, _32119_);
  and _77753_ (_32124_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  and _77754_ (_32125_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  or _77755_ (_32126_, _32125_, _32124_);
  and _77756_ (_32127_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  and _77757_ (_32128_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  or _77758_ (_32129_, _32128_, _32127_);
  or _77759_ (_32130_, _32129_, _32126_);
  or _77760_ (_32131_, _32130_, _32123_);
  and _77761_ (_32132_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and _77762_ (_32133_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  or _77763_ (_32134_, _32133_, _32132_);
  and _77764_ (_32135_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and _77765_ (_32136_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or _77766_ (_32137_, _32136_, _32135_);
  or _77767_ (_32138_, _32137_, _32134_);
  and _77768_ (_32139_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  and _77769_ (_32140_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  or _77770_ (_32141_, _32140_, _32139_);
  and _77771_ (_32142_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and _77772_ (_32143_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or _77773_ (_32144_, _32143_, _32142_);
  or _77774_ (_32145_, _32144_, _32141_);
  or _77775_ (_32146_, _32145_, _32138_);
  or _77776_ (_32147_, _32146_, _32131_);
  or _77777_ (_32148_, _32147_, _32116_);
  and _77778_ (_32149_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  and _77779_ (_32150_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or _77780_ (_32151_, _32150_, _32149_);
  and _77781_ (_32152_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and _77782_ (_32153_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or _77783_ (_32154_, _32153_, _32152_);
  or _77784_ (_32155_, _32154_, _32151_);
  and _77785_ (_32156_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  and _77786_ (_32157_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  nor _77787_ (_32158_, _32157_, _32156_);
  and _77788_ (_32159_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and _77789_ (_32160_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  nor _77790_ (_32161_, _32160_, _32159_);
  nand _77791_ (_32162_, _32161_, _32158_);
  or _77792_ (_32163_, _32162_, _32155_);
  and _77793_ (_32164_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and _77794_ (_32165_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or _77795_ (_32166_, _32165_, _32164_);
  and _77796_ (_32167_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  and _77797_ (_32168_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  or _77798_ (_32169_, _32168_, _32167_);
  or _77799_ (_32170_, _32169_, _32166_);
  and _77800_ (_32171_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  and _77801_ (_32172_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or _77802_ (_32173_, _32172_, _32171_);
  and _77803_ (_32174_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and _77804_ (_32175_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  or _77805_ (_32176_, _32175_, _32174_);
  or _77806_ (_32177_, _32176_, _32173_);
  or _77807_ (_32178_, _32177_, _32170_);
  or _77808_ (_32179_, _32178_, _32163_);
  and _77809_ (_32180_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and _77810_ (_32181_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  or _77811_ (_32182_, _32181_, _32180_);
  and _77812_ (_32183_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and _77813_ (_32184_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or _77814_ (_32185_, _32184_, _32183_);
  or _77815_ (_32186_, _32185_, _32182_);
  and _77816_ (_32187_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and _77817_ (_32188_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  or _77818_ (_32189_, _32188_, _32187_);
  and _77819_ (_32190_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  and _77820_ (_32191_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or _77821_ (_32192_, _32191_, _32190_);
  or _77822_ (_32193_, _32192_, _32189_);
  or _77823_ (_32194_, _32193_, _32186_);
  and _77824_ (_32195_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and _77825_ (_32196_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  or _77826_ (_32197_, _32196_, _32195_);
  and _77827_ (_32198_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and _77828_ (_32199_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  or _77829_ (_32200_, _32199_, _32198_);
  or _77830_ (_32201_, _32200_, _32197_);
  and _77831_ (_32202_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  and _77832_ (_32203_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or _77833_ (_32204_, _32203_, _32202_);
  and _77834_ (_32205_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and _77835_ (_32206_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  or _77836_ (_32207_, _32206_, _32205_);
  or _77837_ (_32208_, _32207_, _32204_);
  or _77838_ (_32209_, _32208_, _32201_);
  or _77839_ (_32210_, _32209_, _32194_);
  or _77840_ (_32211_, _32210_, _32179_);
  or _77841_ (_32212_, _32211_, _32148_);
  and _77842_ (_32213_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and _77843_ (_32214_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  nor _77844_ (_32215_, _32214_, _32213_);
  and _77845_ (_32216_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  and _77846_ (_32217_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor _77847_ (_32218_, _32217_, _32216_);
  nand _77848_ (_32219_, _32218_, _32215_);
  and _77849_ (_32220_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and _77850_ (_32221_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or _77851_ (_32222_, _32221_, _32220_);
  and _77852_ (_32223_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  and _77853_ (_32224_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or _77854_ (_32225_, _32224_, _32223_);
  or _77855_ (_32226_, _32225_, _32222_);
  or _77856_ (_32227_, _32226_, _32219_);
  and _77857_ (_32228_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and _77858_ (_32229_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or _77859_ (_32230_, _32229_, _32228_);
  and _77860_ (_32231_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  and _77861_ (_32232_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or _77862_ (_32233_, _32232_, _32231_);
  or _77863_ (_32234_, _32233_, _32230_);
  and _77864_ (_32235_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and _77865_ (_32236_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or _77866_ (_32237_, _32236_, _32235_);
  and _77867_ (_32238_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and _77868_ (_32239_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or _77869_ (_32240_, _32239_, _32238_);
  or _77870_ (_32241_, _32240_, _32237_);
  or _77871_ (_32242_, _32241_, _32234_);
  or _77872_ (_32243_, _32242_, _32227_);
  and _77873_ (_32244_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and _77874_ (_32245_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or _77875_ (_32246_, _32245_, _32244_);
  and _77876_ (_32247_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and _77877_ (_32248_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or _77878_ (_32249_, _32248_, _32247_);
  or _77879_ (_32250_, _32249_, _32246_);
  and _77880_ (_32251_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  and _77881_ (_32252_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or _77882_ (_32253_, _32252_, _32251_);
  and _77883_ (_32254_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and _77884_ (_32255_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or _77885_ (_32256_, _32255_, _32254_);
  or _77886_ (_32257_, _32256_, _32253_);
  or _77887_ (_32258_, _32257_, _32250_);
  and _77888_ (_32259_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and _77889_ (_32260_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or _77890_ (_32261_, _32260_, _32259_);
  and _77891_ (_32262_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and _77892_ (_32263_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or _77893_ (_32264_, _32263_, _32262_);
  or _77894_ (_32265_, _32264_, _32261_);
  and _77895_ (_32266_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  and _77896_ (_32267_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or _77897_ (_32268_, _32267_, _32266_);
  and _77898_ (_32269_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and _77899_ (_32270_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or _77900_ (_32271_, _32270_, _32269_);
  or _77901_ (_32272_, _32271_, _32268_);
  or _77902_ (_32273_, _32272_, _32265_);
  or _77903_ (_32274_, _32273_, _32258_);
  or _77904_ (_32275_, _32274_, _32243_);
  and _77905_ (_32276_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and _77906_ (_32277_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  or _77907_ (_32278_, _32277_, _32276_);
  and _77908_ (_32279_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  and _77909_ (_32280_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  or _77910_ (_32281_, _32280_, _32279_);
  or _77911_ (_32282_, _32281_, _32278_);
  and _77912_ (_32283_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  and _77913_ (_32284_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or _77914_ (_32285_, _32284_, _32283_);
  and _77915_ (_32286_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  and _77916_ (_32287_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  or _77917_ (_32288_, _32287_, _32286_);
  or _77918_ (_32289_, _32288_, _32285_);
  or _77919_ (_32290_, _32289_, _32282_);
  and _77920_ (_32291_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and _77921_ (_32292_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  nor _77922_ (_32293_, _32292_, _32291_);
  and _77923_ (_32294_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  and _77924_ (_32295_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  nor _77925_ (_32296_, _32295_, _32294_);
  nand _77926_ (_32297_, _32296_, _32293_);
  and _77927_ (_32298_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and _77928_ (_32299_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or _77929_ (_32300_, _32299_, _32298_);
  and _77930_ (_32301_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and _77931_ (_32302_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or _77932_ (_32303_, _32302_, _32301_);
  or _77933_ (_32304_, _32303_, _32300_);
  or _77934_ (_32305_, _32304_, _32297_);
  or _77935_ (_32306_, _32305_, _32290_);
  and _77936_ (_32307_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and _77937_ (_32308_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or _77938_ (_32309_, _32308_, _32307_);
  and _77939_ (_32310_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and _77940_ (_32311_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  or _77941_ (_32312_, _32311_, _32310_);
  or _77942_ (_32313_, _32312_, _32309_);
  and _77943_ (_32314_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and _77944_ (_32315_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  or _77945_ (_32316_, _32315_, _32314_);
  and _77946_ (_32317_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and _77947_ (_32318_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or _77948_ (_32319_, _32318_, _32317_);
  or _77949_ (_32320_, _32319_, _32316_);
  or _77950_ (_32321_, _32320_, _32313_);
  and _77951_ (_32322_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and _77952_ (_32323_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or _77953_ (_32324_, _32323_, _32322_);
  and _77954_ (_32325_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  and _77955_ (_32326_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  or _77956_ (_32327_, _32326_, _32325_);
  or _77957_ (_32328_, _32327_, _32324_);
  and _77958_ (_32329_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  and _77959_ (_32330_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or _77960_ (_32331_, _32330_, _32329_);
  and _77961_ (_32332_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and _77962_ (_32333_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or _77963_ (_32334_, _32333_, _32332_);
  or _77964_ (_32335_, _32334_, _32331_);
  or _77965_ (_32336_, _32335_, _32328_);
  or _77966_ (_32337_, _32336_, _32321_);
  or _77967_ (_32338_, _32337_, _32306_);
  or _77968_ (_32339_, _32338_, _32275_);
  or _77969_ (_32340_, _32339_, _32212_);
  and _77970_ (_32341_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and _77971_ (_32342_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or _77972_ (_32343_, _32342_, _32341_);
  and _77973_ (_32344_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and _77974_ (_32345_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or _77975_ (_32346_, _32345_, _32344_);
  or _77976_ (_32347_, _32346_, _32343_);
  and _77977_ (_32348_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  and _77978_ (_32349_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _77979_ (_32350_, _32349_, _32348_);
  and _77980_ (_32351_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and _77981_ (_32352_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or _77982_ (_32353_, _32352_, _32351_);
  or _77983_ (_32354_, _32353_, _32350_);
  or _77984_ (_32355_, _32354_, _32347_);
  and _77985_ (_32356_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  and _77986_ (_32357_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  or _77987_ (_32358_, _32357_, _32356_);
  and _77988_ (_32359_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  and _77989_ (_32360_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  or _77990_ (_32361_, _32360_, _32359_);
  or _77991_ (_32362_, _32361_, _32358_);
  and _77992_ (_32363_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  and _77993_ (_32364_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or _77994_ (_32365_, _32364_, _32363_);
  and _77995_ (_32366_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  and _77996_ (_32367_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  or _77997_ (_32368_, _32367_, _32366_);
  or _77998_ (_32369_, _32368_, _32365_);
  or _77999_ (_32370_, _32369_, _32362_);
  or _78000_ (_32371_, _32370_, _32355_);
  and _78001_ (_32372_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and _78002_ (_32373_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or _78003_ (_32374_, _32373_, _32372_);
  and _78004_ (_32375_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and _78005_ (_32376_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or _78006_ (_32377_, _32376_, _32375_);
  or _78007_ (_32378_, _32377_, _32374_);
  and _78008_ (_32379_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and _78009_ (_32380_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  nor _78010_ (_32381_, _32380_, _32379_);
  and _78011_ (_32382_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  and _78012_ (_32383_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  nor _78013_ (_32384_, _32383_, _32382_);
  nand _78014_ (_32385_, _32384_, _32381_);
  or _78015_ (_32386_, _32385_, _32378_);
  and _78016_ (_32387_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  and _78017_ (_32388_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or _78018_ (_32389_, _32388_, _32387_);
  and _78019_ (_32390_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and _78020_ (_32391_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or _78021_ (_32392_, _32391_, _32390_);
  or _78022_ (_32393_, _32392_, _32389_);
  and _78023_ (_32394_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and _78024_ (_32395_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or _78025_ (_32396_, _32395_, _32394_);
  and _78026_ (_32397_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  and _78027_ (_32398_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or _78028_ (_32399_, _32398_, _32397_);
  or _78029_ (_32400_, _32399_, _32396_);
  or _78030_ (_32401_, _32400_, _32393_);
  or _78031_ (_32402_, _32401_, _32386_);
  or _78032_ (_32403_, _32402_, _32371_);
  and _78033_ (_32404_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and _78034_ (_32405_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or _78035_ (_32406_, _32405_, _32404_);
  and _78036_ (_32407_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  and _78037_ (_32408_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or _78038_ (_32409_, _32408_, _32407_);
  or _78039_ (_32410_, _32409_, _32406_);
  and _78040_ (_32411_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and _78041_ (_32412_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  nor _78042_ (_32413_, _32412_, _32411_);
  and _78043_ (_32414_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  and _78044_ (_32415_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  nor _78045_ (_32416_, _32415_, _32414_);
  nand _78046_ (_32417_, _32416_, _32413_);
  or _78047_ (_32418_, _32417_, _32410_);
  and _78048_ (_32419_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and _78049_ (_32420_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  and _78050_ (_32421_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  or _78051_ (_32422_, _32421_, _32420_);
  or _78052_ (_32423_, _32422_, _32419_);
  and _78053_ (_32424_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  and _78054_ (_32425_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or _78055_ (_32426_, _32425_, _32424_);
  and _78056_ (_32427_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and _78057_ (_32428_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  or _78058_ (_32429_, _32428_, _32427_);
  or _78059_ (_32430_, _32429_, _32426_);
  or _78060_ (_32431_, _32430_, _32423_);
  or _78061_ (_32432_, _32431_, _32418_);
  and _78062_ (_32433_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  and _78063_ (_32434_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  nor _78064_ (_32435_, _32434_, _32433_);
  and _78065_ (_32436_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  and _78066_ (_32437_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  nor _78067_ (_32438_, _32437_, _32436_);
  nand _78068_ (_32439_, _32438_, _32435_);
  and _78069_ (_32440_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and _78070_ (_32441_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  or _78071_ (_32442_, _32441_, _32440_);
  and _78072_ (_32443_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and _78073_ (_32444_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or _78074_ (_32445_, _32444_, _32443_);
  or _78075_ (_32446_, _32445_, _32442_);
  or _78076_ (_32447_, _32446_, _32439_);
  and _78077_ (_32448_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  and _78078_ (_32449_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or _78079_ (_32450_, _32449_, _32448_);
  and _78080_ (_32451_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  and _78081_ (_32452_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or _78082_ (_32453_, _32452_, _32451_);
  or _78083_ (_32454_, _32453_, _32450_);
  and _78084_ (_32455_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  and _78085_ (_32456_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or _78086_ (_32457_, _32456_, _32455_);
  and _78087_ (_32458_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  and _78088_ (_32459_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or _78089_ (_32460_, _32459_, _32458_);
  or _78090_ (_32461_, _32460_, _32457_);
  or _78091_ (_32462_, _32461_, _32454_);
  or _78092_ (_32463_, _32462_, _32447_);
  or _78093_ (_32464_, _32463_, _32432_);
  or _78094_ (_32465_, _32464_, _32403_);
  and _78095_ (_32466_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  and _78096_ (_32467_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  nor _78097_ (_32468_, _32467_, _32466_);
  and _78098_ (_32469_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  and _78099_ (_32470_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  nor _78100_ (_32471_, _32470_, _32469_);
  nand _78101_ (_32472_, _32471_, _32468_);
  and _78102_ (_32473_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  and _78103_ (_32474_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or _78104_ (_32475_, _32474_, _32473_);
  and _78105_ (_32476_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and _78106_ (_32477_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  or _78107_ (_32478_, _32477_, _32476_);
  or _78108_ (_32479_, _32478_, _32475_);
  or _78109_ (_32480_, _32479_, _32472_);
  and _78110_ (_32481_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and _78111_ (_32482_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  nor _78112_ (_32483_, _32482_, _32481_);
  and _78113_ (_32484_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and _78114_ (_32485_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  nor _78115_ (_32486_, _32485_, _32484_);
  nand _78116_ (_32487_, _32486_, _32483_);
  and _78117_ (_32488_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  and _78118_ (_32489_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or _78119_ (_32490_, _32489_, _32488_);
  and _78120_ (_32491_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and _78121_ (_32492_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or _78122_ (_32493_, _32492_, _32491_);
  or _78123_ (_32494_, _32493_, _32490_);
  or _78124_ (_32495_, _32494_, _32487_);
  or _78125_ (_32496_, _32495_, _32480_);
  and _78126_ (_32497_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  and _78127_ (_32498_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  nor _78128_ (_32499_, _32498_, _32497_);
  and _78129_ (_32500_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  and _78130_ (_32501_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor _78131_ (_32502_, _32501_, _32500_);
  nand _78132_ (_32503_, _32502_, _32499_);
  and _78133_ (_32504_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and _78134_ (_32505_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  or _78135_ (_32506_, _32505_, _32504_);
  and _78136_ (_32507_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  and _78137_ (_32508_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  or _78138_ (_32509_, _32508_, _32507_);
  or _78139_ (_32510_, _32509_, _32506_);
  or _78140_ (_32511_, _32510_, _32503_);
  and _78141_ (_32512_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  and _78142_ (_32513_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  nor _78143_ (_32514_, _32513_, _32512_);
  and _78144_ (_32515_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and _78145_ (_32516_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  nor _78146_ (_32517_, _32516_, _32515_);
  nand _78147_ (_32518_, _32517_, _32514_);
  and _78148_ (_32519_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  and _78149_ (_32520_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or _78150_ (_32521_, _32520_, _32519_);
  and _78151_ (_32522_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  and _78152_ (_32523_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or _78153_ (_32524_, _32523_, _32522_);
  or _78154_ (_32525_, _32524_, _32521_);
  or _78155_ (_32526_, _32525_, _32518_);
  or _78156_ (_32527_, _32526_, _32511_);
  or _78157_ (_32528_, _32527_, _32496_);
  and _78158_ (_32529_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and _78159_ (_32530_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or _78160_ (_32531_, _32530_, _32529_);
  and _78161_ (_32532_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and _78162_ (_32533_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or _78163_ (_32534_, _32533_, _32532_);
  or _78164_ (_32535_, _32534_, _32531_);
  and _78165_ (_32536_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  and _78166_ (_32537_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or _78167_ (_32538_, _32537_, _32536_);
  and _78168_ (_32539_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and _78169_ (_32540_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  or _78170_ (_32541_, _32540_, _32539_);
  or _78171_ (_32542_, _32541_, _32538_);
  or _78172_ (_32543_, _32542_, _32535_);
  and _78173_ (_32544_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  and _78174_ (_32545_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or _78175_ (_32546_, _32545_, _32544_);
  and _78176_ (_32547_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  and _78177_ (_32548_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or _78178_ (_32549_, _32548_, _32547_);
  or _78179_ (_32550_, _32549_, _32546_);
  and _78180_ (_32551_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  and _78181_ (_32552_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  nor _78182_ (_32553_, _32552_, _32551_);
  and _78183_ (_32554_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and _78184_ (_32555_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  nor _78185_ (_32556_, _32555_, _32554_);
  nand _78186_ (_32557_, _32556_, _32553_);
  or _78187_ (_32558_, _32557_, _32550_);
  or _78188_ (_32559_, _32558_, _32543_);
  and _78189_ (_32560_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  and _78190_ (_32561_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or _78191_ (_32562_, _32561_, _32560_);
  and _78192_ (_32563_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  and _78193_ (_32564_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  or _78194_ (_32565_, _32564_, _32563_);
  or _78195_ (_32566_, _32565_, _32562_);
  and _78196_ (_32567_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and _78197_ (_32568_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  or _78198_ (_32569_, _32568_, _32567_);
  and _78199_ (_32570_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and _78200_ (_32571_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  or _78201_ (_32572_, _32571_, _32570_);
  or _78202_ (_32573_, _32572_, _32569_);
  or _78203_ (_32574_, _32573_, _32566_);
  and _78204_ (_32575_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  and _78205_ (_32576_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  or _78206_ (_32577_, _32576_, _32575_);
  and _78207_ (_32578_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  and _78208_ (_32579_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  or _78209_ (_32580_, _32579_, _32578_);
  or _78210_ (_32581_, _32580_, _32577_);
  and _78211_ (_32582_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and _78212_ (_32583_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or _78213_ (_32584_, _32583_, _32582_);
  and _78214_ (_32585_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  and _78215_ (_32586_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or _78216_ (_32587_, _32586_, _32585_);
  or _78217_ (_32588_, _32587_, _32584_);
  or _78218_ (_32589_, _32588_, _32581_);
  or _78219_ (_32590_, _32589_, _32574_);
  or _78220_ (_32591_, _32590_, _32559_);
  or _78221_ (_32592_, _32591_, _32528_);
  or _78222_ (_32593_, _32592_, _32465_);
  nor _78223_ (_32594_, _32593_, _32340_);
  and _78224_ (_32595_, _32594_, _32085_);
  nor _78225_ (_32596_, _30010_, iram_op1_reg[5]);
  nor _78226_ (_32597_, _32596_, _31043_);
  and _78227_ (_32598_, _32597_, _32595_);
  or _78228_ (_32599_, _32598_, _32083_);
  or _78229_ (_32600_, _32599_, _32082_);
  nor _78230_ (_32601_, _32597_, _32595_);
  and _78231_ (_32602_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  not _78232_ (_32603_, _32602_);
  and _78233_ (_32604_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and _78234_ (_32605_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  nor _78235_ (_32606_, _32605_, _32604_);
  and _78236_ (_32607_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  and _78237_ (_32608_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  nor _78238_ (_32609_, _32608_, _32607_);
  and _78239_ (_32610_, _32609_, _32606_);
  and _78240_ (_32611_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and _78241_ (_32612_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  nor _78242_ (_32613_, _32612_, _32611_);
  and _78243_ (_32614_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and _78244_ (_32615_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  nor _78245_ (_32616_, _32615_, _32614_);
  and _78246_ (_32617_, _32616_, _32613_);
  and _78247_ (_32618_, _32617_, _32610_);
  and _78248_ (_32619_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  and _78249_ (_32620_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  nor _78250_ (_32621_, _32620_, _32619_);
  and _78251_ (_32622_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and _78252_ (_32623_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  nor _78253_ (_32624_, _32623_, _32622_);
  and _78254_ (_32625_, _32624_, _32621_);
  and _78255_ (_32626_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  and _78256_ (_32627_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  nor _78257_ (_32628_, _32627_, _32626_);
  and _78258_ (_32629_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and _78259_ (_32630_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  nor _78260_ (_32631_, _32630_, _32629_);
  and _78261_ (_32632_, _32631_, _32628_);
  and _78262_ (_32633_, _32632_, _32625_);
  and _78263_ (_32634_, _32633_, _32618_);
  and _78264_ (_32635_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  and _78265_ (_32636_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  nor _78266_ (_32637_, _32636_, _32635_);
  and _78267_ (_32638_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and _78268_ (_32639_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  nor _78269_ (_32640_, _32639_, _32638_);
  and _78270_ (_32641_, _32640_, _32637_);
  and _78271_ (_32642_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  and _78272_ (_32643_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  nor _78273_ (_32644_, _32643_, _32642_);
  and _78274_ (_32645_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  and _78275_ (_32646_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  nor _78276_ (_32647_, _32646_, _32645_);
  and _78277_ (_32648_, _32647_, _32644_);
  and _78278_ (_32649_, _32648_, _32641_);
  and _78279_ (_32650_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and _78280_ (_32651_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  nor _78281_ (_32652_, _32651_, _32650_);
  and _78282_ (_32653_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  and _78283_ (_32654_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  nor _78284_ (_32655_, _32654_, _32653_);
  and _78285_ (_32656_, _32655_, _32652_);
  and _78286_ (_32657_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and _78287_ (_32658_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  nor _78288_ (_32659_, _32658_, _32657_);
  and _78289_ (_32660_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  and _78290_ (_32661_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  nor _78291_ (_32662_, _32661_, _32660_);
  and _78292_ (_32663_, _32662_, _32659_);
  and _78293_ (_32664_, _32663_, _32656_);
  and _78294_ (_32665_, _32664_, _32649_);
  and _78295_ (_32666_, _32665_, _32634_);
  and _78296_ (_32667_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and _78297_ (_32668_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  nor _78298_ (_32669_, _32668_, _32667_);
  and _78299_ (_32670_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  and _78300_ (_32671_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  nor _78301_ (_32672_, _32671_, _32670_);
  and _78302_ (_32673_, _32672_, _32669_);
  and _78303_ (_32674_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and _78304_ (_32675_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  nor _78305_ (_32676_, _32675_, _32674_);
  and _78306_ (_32677_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  and _78307_ (_32678_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  nor _78308_ (_32679_, _32678_, _32677_);
  and _78309_ (_32680_, _32679_, _32676_);
  and _78310_ (_32681_, _32680_, _32673_);
  and _78311_ (_32682_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  and _78312_ (_32683_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  nor _78313_ (_32684_, _32683_, _32682_);
  and _78314_ (_32685_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and _78315_ (_32686_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  nor _78316_ (_32687_, _32686_, _32685_);
  and _78317_ (_32688_, _32687_, _32684_);
  and _78318_ (_32689_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  and _78319_ (_32690_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  nor _78320_ (_32691_, _32690_, _32689_);
  and _78321_ (_32692_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and _78322_ (_32693_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  nor _78323_ (_32694_, _32693_, _32692_);
  and _78324_ (_32695_, _32694_, _32691_);
  and _78325_ (_32696_, _32695_, _32688_);
  and _78326_ (_32697_, _32696_, _32681_);
  and _78327_ (_32698_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  and _78328_ (_32699_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  nor _78329_ (_32700_, _32699_, _32698_);
  and _78330_ (_32701_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and _78331_ (_32702_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  nor _78332_ (_32703_, _32702_, _32701_);
  and _78333_ (_32704_, _32703_, _32700_);
  and _78334_ (_32705_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and _78335_ (_32706_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  nor _78336_ (_32707_, _32706_, _32705_);
  and _78337_ (_32708_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  and _78338_ (_32709_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  nor _78339_ (_32710_, _32709_, _32708_);
  and _78340_ (_32711_, _32710_, _32707_);
  and _78341_ (_32712_, _32711_, _32704_);
  and _78342_ (_32713_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  and _78343_ (_32714_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  nor _78344_ (_32715_, _32714_, _32713_);
  and _78345_ (_32716_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and _78346_ (_32717_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  nor _78347_ (_32718_, _32717_, _32716_);
  and _78348_ (_32719_, _32718_, _32715_);
  and _78349_ (_32720_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  and _78350_ (_32721_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  nor _78351_ (_32722_, _32721_, _32720_);
  and _78352_ (_32723_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and _78353_ (_32724_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  nor _78354_ (_32725_, _32724_, _32723_);
  and _78355_ (_32726_, _32725_, _32722_);
  and _78356_ (_32727_, _32726_, _32719_);
  and _78357_ (_32728_, _32727_, _32712_);
  and _78358_ (_32729_, _32728_, _32697_);
  and _78359_ (_32730_, _32729_, _32666_);
  and _78360_ (_32731_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  and _78361_ (_32732_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  nor _78362_ (_32733_, _32732_, _32731_);
  and _78363_ (_32734_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and _78364_ (_32735_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  nor _78365_ (_32736_, _32735_, _32734_);
  and _78366_ (_32737_, _32736_, _32733_);
  and _78367_ (_32738_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  and _78368_ (_32739_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  nor _78369_ (_32740_, _32739_, _32738_);
  and _78370_ (_32741_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and _78371_ (_32742_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  nor _78372_ (_32743_, _32742_, _32741_);
  and _78373_ (_32744_, _32743_, _32740_);
  and _78374_ (_32745_, _32744_, _32737_);
  and _78375_ (_32746_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and _78376_ (_32747_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  nor _78377_ (_32748_, _32747_, _32746_);
  and _78378_ (_32749_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  and _78379_ (_32750_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  nor _78380_ (_32751_, _32750_, _32749_);
  and _78381_ (_32752_, _32751_, _32748_);
  and _78382_ (_32753_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and _78383_ (_32754_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  nor _78384_ (_32755_, _32754_, _32753_);
  and _78385_ (_32756_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and _78386_ (_32757_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  nor _78387_ (_32758_, _32757_, _32756_);
  and _78388_ (_32759_, _32758_, _32755_);
  and _78389_ (_32760_, _32759_, _32752_);
  and _78390_ (_32761_, _32760_, _32745_);
  and _78391_ (_32762_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  and _78392_ (_32763_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  nor _78393_ (_32764_, _32763_, _32762_);
  and _78394_ (_32765_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and _78395_ (_32766_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  nor _78396_ (_32767_, _32766_, _32765_);
  and _78397_ (_32768_, _32767_, _32764_);
  and _78398_ (_32769_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  and _78399_ (_32770_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  nor _78400_ (_32771_, _32770_, _32769_);
  and _78401_ (_32772_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  and _78402_ (_32773_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  nor _78403_ (_32774_, _32773_, _32772_);
  and _78404_ (_32775_, _32774_, _32771_);
  and _78405_ (_32776_, _32775_, _32768_);
  and _78406_ (_32777_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and _78407_ (_32778_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  nor _78408_ (_32779_, _32778_, _32777_);
  and _78409_ (_32780_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  and _78410_ (_32781_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  nor _78411_ (_32782_, _32781_, _32780_);
  and _78412_ (_32783_, _32782_, _32779_);
  and _78413_ (_32784_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and _78414_ (_32785_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  nor _78415_ (_32786_, _32785_, _32784_);
  and _78416_ (_32787_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  and _78417_ (_32788_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  nor _78418_ (_32789_, _32788_, _32787_);
  and _78419_ (_32790_, _32789_, _32786_);
  and _78420_ (_32791_, _32790_, _32783_);
  and _78421_ (_32792_, _32791_, _32776_);
  and _78422_ (_32793_, _32792_, _32761_);
  and _78423_ (_32794_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and _78424_ (_32795_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  nor _78425_ (_32796_, _32795_, _32794_);
  and _78426_ (_32797_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  and _78427_ (_32798_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  nor _78428_ (_32799_, _32798_, _32797_);
  and _78429_ (_32800_, _32799_, _32796_);
  and _78430_ (_32801_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  and _78431_ (_32802_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  nor _78432_ (_32803_, _32802_, _32801_);
  and _78433_ (_32804_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and _78434_ (_32805_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  nor _78435_ (_32806_, _32805_, _32804_);
  and _78436_ (_32807_, _32806_, _32803_);
  and _78437_ (_32808_, _32807_, _32800_);
  and _78438_ (_32809_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  and _78439_ (_32810_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  nor _78440_ (_32811_, _32810_, _32809_);
  and _78441_ (_32812_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and _78442_ (_32813_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  nor _78443_ (_32814_, _32813_, _32812_);
  and _78444_ (_32815_, _32814_, _32811_);
  and _78445_ (_32816_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  and _78446_ (_32817_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  nor _78447_ (_32818_, _32817_, _32816_);
  and _78448_ (_32819_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and _78449_ (_32820_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  nor _78450_ (_32821_, _32820_, _32819_);
  and _78451_ (_32822_, _32821_, _32818_);
  and _78452_ (_32823_, _32822_, _32815_);
  and _78453_ (_32824_, _32823_, _32808_);
  and _78454_ (_32825_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  and _78455_ (_32826_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  nor _78456_ (_32827_, _32826_, _32825_);
  and _78457_ (_32828_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and _78458_ (_32829_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  nor _78459_ (_32830_, _32829_, _32828_);
  and _78460_ (_32831_, _32830_, _32827_);
  and _78461_ (_32832_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  and _78462_ (_32833_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  nor _78463_ (_32834_, _32833_, _32832_);
  and _78464_ (_32835_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  and _78465_ (_32836_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  nor _78466_ (_32837_, _32836_, _32835_);
  and _78467_ (_32838_, _32837_, _32834_);
  and _78468_ (_32839_, _32838_, _32831_);
  and _78469_ (_32840_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and _78470_ (_32841_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  nor _78471_ (_32842_, _32841_, _32840_);
  and _78472_ (_32843_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  and _78473_ (_32844_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  nor _78474_ (_32845_, _32844_, _32843_);
  and _78475_ (_32846_, _32845_, _32842_);
  and _78476_ (_32847_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and _78477_ (_32848_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  nor _78478_ (_32849_, _32848_, _32847_);
  and _78479_ (_32850_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  and _78480_ (_32851_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  nor _78481_ (_32852_, _32851_, _32850_);
  and _78482_ (_32853_, _32852_, _32849_);
  and _78483_ (_32854_, _32853_, _32846_);
  and _78484_ (_32855_, _32854_, _32839_);
  and _78485_ (_32856_, _32855_, _32824_);
  and _78486_ (_32857_, _32856_, _32793_);
  and _78487_ (_32858_, _32857_, _32730_);
  and _78488_ (_32859_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  and _78489_ (_32860_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  nor _78490_ (_32861_, _32860_, _32859_);
  and _78491_ (_32862_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and _78492_ (_32863_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  nor _78493_ (_32864_, _32863_, _32862_);
  and _78494_ (_32865_, _32864_, _32861_);
  and _78495_ (_32866_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  and _78496_ (_32867_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  nor _78497_ (_32868_, _32867_, _32866_);
  and _78498_ (_32869_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  and _78499_ (_32870_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  nor _78500_ (_32871_, _32870_, _32869_);
  and _78501_ (_32872_, _32871_, _32868_);
  and _78502_ (_32873_, _32872_, _32865_);
  and _78503_ (_32874_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and _78504_ (_32875_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  nor _78505_ (_32876_, _32875_, _32874_);
  and _78506_ (_32877_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  and _78507_ (_32878_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  nor _78508_ (_32879_, _32878_, _32877_);
  and _78509_ (_32880_, _32879_, _32876_);
  and _78510_ (_32881_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and _78511_ (_32882_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  nor _78512_ (_32883_, _32882_, _32881_);
  and _78513_ (_32884_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  and _78514_ (_32885_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  nor _78515_ (_32886_, _32885_, _32884_);
  and _78516_ (_32887_, _32886_, _32883_);
  and _78517_ (_32888_, _32887_, _32880_);
  and _78518_ (_32889_, _32888_, _32873_);
  and _78519_ (_32890_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and _78520_ (_32891_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  nor _78521_ (_32892_, _32891_, _32890_);
  and _78522_ (_32893_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  and _78523_ (_32894_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  nor _78524_ (_32895_, _32894_, _32893_);
  and _78525_ (_32896_, _32895_, _32892_);
  and _78526_ (_32897_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and _78527_ (_32898_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  nor _78528_ (_32899_, _32898_, _32897_);
  and _78529_ (_32900_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and _78530_ (_32901_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  nor _78531_ (_32902_, _32901_, _32900_);
  and _78532_ (_32903_, _32902_, _32899_);
  and _78533_ (_32904_, _32903_, _32896_);
  and _78534_ (_32905_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  and _78535_ (_32906_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  nor _78536_ (_32907_, _32906_, _32905_);
  and _78537_ (_32908_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and _78538_ (_32909_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  nor _78539_ (_32910_, _32909_, _32908_);
  and _78540_ (_32911_, _32910_, _32907_);
  and _78541_ (_32912_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  and _78542_ (_32913_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  nor _78543_ (_32914_, _32913_, _32912_);
  and _78544_ (_32915_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and _78545_ (_32916_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  nor _78546_ (_32917_, _32916_, _32915_);
  and _78547_ (_32918_, _32917_, _32914_);
  and _78548_ (_32919_, _32918_, _32911_);
  and _78549_ (_32920_, _32919_, _32904_);
  and _78550_ (_32921_, _32920_, _32889_);
  and _78551_ (_32922_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and _78552_ (_32923_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  nor _78553_ (_32924_, _32923_, _32922_);
  and _78554_ (_32925_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  and _78555_ (_32926_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  nor _78556_ (_32927_, _32926_, _32925_);
  and _78557_ (_32928_, _32927_, _32924_);
  and _78558_ (_32929_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and _78559_ (_32930_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  nor _78560_ (_32931_, _32930_, _32929_);
  and _78561_ (_32932_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  and _78562_ (_32933_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  nor _78563_ (_32934_, _32933_, _32932_);
  and _78564_ (_32935_, _32934_, _32931_);
  and _78565_ (_32936_, _32935_, _32928_);
  and _78566_ (_32937_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  and _78567_ (_32938_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  nor _78568_ (_32939_, _32938_, _32937_);
  and _78569_ (_32940_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and _78570_ (_32941_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  nor _78571_ (_32942_, _32941_, _32940_);
  and _78572_ (_32943_, _32942_, _32939_);
  and _78573_ (_32944_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  and _78574_ (_32945_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  nor _78575_ (_32946_, _32945_, _32944_);
  and _78576_ (_32947_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and _78577_ (_32948_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  nor _78578_ (_32949_, _32948_, _32947_);
  and _78579_ (_32950_, _32949_, _32946_);
  and _78580_ (_32951_, _32950_, _32943_);
  and _78581_ (_32952_, _32951_, _32936_);
  and _78582_ (_32953_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and _78583_ (_32954_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  nor _78584_ (_32955_, _32954_, _32953_);
  and _78585_ (_32956_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  and _78586_ (_32957_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  nor _78587_ (_32958_, _32957_, _32956_);
  and _78588_ (_32959_, _32958_, _32955_);
  and _78589_ (_32960_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  and _78590_ (_32961_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  nor _78591_ (_32962_, _32961_, _32960_);
  and _78592_ (_32963_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  and _78593_ (_32964_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  nor _78594_ (_32965_, _32964_, _32963_);
  and _78595_ (_32966_, _32965_, _32962_);
  and _78596_ (_32967_, _32966_, _32959_);
  and _78597_ (_32968_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  and _78598_ (_32969_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  nor _78599_ (_32970_, _32969_, _32968_);
  and _78600_ (_32971_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and _78601_ (_32972_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  nor _78602_ (_32973_, _32972_, _32971_);
  and _78603_ (_32974_, _32973_, _32970_);
  and _78604_ (_32975_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and _78605_ (_32976_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  nor _78606_ (_32977_, _32976_, _32975_);
  and _78607_ (_32978_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  and _78608_ (_32979_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  nor _78609_ (_32980_, _32979_, _32978_);
  and _78610_ (_32981_, _32980_, _32977_);
  and _78611_ (_32982_, _32981_, _32974_);
  and _78612_ (_32983_, _32982_, _32967_);
  and _78613_ (_32984_, _32983_, _32952_);
  and _78614_ (_32985_, _32984_, _32921_);
  and _78615_ (_32986_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and _78616_ (_32987_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  nor _78617_ (_32988_, _32987_, _32986_);
  and _78618_ (_32989_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  and _78619_ (_32990_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  nor _78620_ (_32991_, _32990_, _32989_);
  and _78621_ (_32992_, _32991_, _32988_);
  and _78622_ (_32993_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and _78623_ (_32994_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  nor _78624_ (_32995_, _32994_, _32993_);
  and _78625_ (_32996_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  and _78626_ (_32997_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  nor _78627_ (_32998_, _32997_, _32996_);
  and _78628_ (_32999_, _32998_, _32995_);
  and _78629_ (_33000_, _32999_, _32992_);
  and _78630_ (_33001_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  and _78631_ (_33002_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  nor _78632_ (_33003_, _33002_, _33001_);
  and _78633_ (_33004_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and _78634_ (_33005_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  nor _78635_ (_33006_, _33005_, _33004_);
  and _78636_ (_33007_, _33006_, _33003_);
  and _78637_ (_33008_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  and _78638_ (_33009_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  nor _78639_ (_33010_, _33009_, _33008_);
  and _78640_ (_33011_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and _78641_ (_33012_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  nor _78642_ (_33013_, _33012_, _33011_);
  and _78643_ (_33014_, _33013_, _33010_);
  and _78644_ (_33015_, _33014_, _33007_);
  and _78645_ (_33016_, _33015_, _33000_);
  and _78646_ (_33017_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and _78647_ (_33018_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  nor _78648_ (_33019_, _33018_, _33017_);
  and _78649_ (_33020_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  and _78650_ (_33021_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  nor _78651_ (_33022_, _33021_, _33020_);
  and _78652_ (_33023_, _33022_, _33019_);
  and _78653_ (_33024_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and _78654_ (_33025_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  nor _78655_ (_33026_, _33025_, _33024_);
  and _78656_ (_33027_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  and _78657_ (_33028_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  nor _78658_ (_33029_, _33028_, _33027_);
  and _78659_ (_33030_, _33029_, _33026_);
  and _78660_ (_33031_, _33030_, _33023_);
  and _78661_ (_33032_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  and _78662_ (_33033_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  nor _78663_ (_33034_, _33033_, _33032_);
  and _78664_ (_33035_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and _78665_ (_33036_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  nor _78666_ (_33037_, _33036_, _33035_);
  and _78667_ (_33038_, _33037_, _33034_);
  and _78668_ (_33039_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  and _78669_ (_33040_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  nor _78670_ (_33041_, _33040_, _33039_);
  and _78671_ (_33042_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and _78672_ (_33043_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  nor _78673_ (_33044_, _33043_, _33042_);
  and _78674_ (_33045_, _33044_, _33041_);
  and _78675_ (_33046_, _33045_, _33038_);
  and _78676_ (_33047_, _33046_, _33031_);
  and _78677_ (_33048_, _33047_, _33016_);
  and _78678_ (_33049_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  and _78679_ (_33050_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  nor _78680_ (_33051_, _33050_, _33049_);
  and _78681_ (_33052_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and _78682_ (_33053_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  nor _78683_ (_33054_, _33053_, _33052_);
  and _78684_ (_33055_, _33054_, _33051_);
  and _78685_ (_33056_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  and _78686_ (_33057_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  nor _78687_ (_33058_, _33057_, _33056_);
  and _78688_ (_33059_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and _78689_ (_33060_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  nor _78690_ (_33061_, _33060_, _33059_);
  and _78691_ (_33062_, _33061_, _33058_);
  and _78692_ (_33063_, _33062_, _33055_);
  and _78693_ (_33064_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and _78694_ (_33065_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  nor _78695_ (_33066_, _33065_, _33064_);
  and _78696_ (_33067_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  and _78697_ (_33068_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  nor _78698_ (_33069_, _33068_, _33067_);
  and _78699_ (_33070_, _33069_, _33066_);
  and _78700_ (_33071_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and _78701_ (_33072_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  nor _78702_ (_33073_, _33072_, _33071_);
  and _78703_ (_33074_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  and _78704_ (_33075_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  nor _78705_ (_33076_, _33075_, _33074_);
  and _78706_ (_33077_, _33076_, _33073_);
  and _78707_ (_33078_, _33077_, _33070_);
  and _78708_ (_33079_, _33078_, _33063_);
  and _78709_ (_33080_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and _78710_ (_33081_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor _78711_ (_33082_, _33081_, _33080_);
  and _78712_ (_33083_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and _78713_ (_33084_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor _78714_ (_33085_, _33084_, _33083_);
  and _78715_ (_33086_, _33085_, _33082_);
  and _78716_ (_33087_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and _78717_ (_33088_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and _78718_ (_33089_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or _78719_ (_33090_, _33089_, _33088_);
  nor _78720_ (_33091_, _33090_, _33087_);
  and _78721_ (_33092_, _33091_, _33086_);
  and _78722_ (_33093_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and _78723_ (_33094_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor _78724_ (_33095_, _33094_, _33093_);
  and _78725_ (_33096_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and _78726_ (_33097_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor _78727_ (_33098_, _33097_, _33096_);
  and _78728_ (_33099_, _33098_, _33095_);
  and _78729_ (_33100_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and _78730_ (_33101_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor _78731_ (_33102_, _33101_, _33100_);
  and _78732_ (_33103_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and _78733_ (_33104_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor _78734_ (_33105_, _33104_, _33103_);
  and _78735_ (_33106_, _33105_, _33102_);
  and _78736_ (_33107_, _33106_, _33099_);
  and _78737_ (_33108_, _33107_, _33092_);
  and _78738_ (_33109_, _33108_, _33079_);
  and _78739_ (_33110_, _33109_, _33048_);
  and _78740_ (_33111_, _33110_, _32985_);
  and _78741_ (_33112_, _33111_, _32858_);
  and _78742_ (_33113_, _33112_, _32603_);
  nor _78743_ (_33114_, _31043_, iram_op1_reg[6]);
  nor _78744_ (_33115_, _33114_, _31044_);
  nor _78745_ (_33116_, _33115_, _33113_);
  or _78746_ (_33117_, _33116_, _32601_);
  and _78747_ (_33118_, _31047_, _31042_);
  and _78748_ (_33119_, _33115_, _33113_);
  or _78749_ (_33120_, _33119_, _33118_);
  or _78750_ (_33121_, _33120_, _33117_);
  or _78751_ (_33122_, _33121_, _32600_);
  or _78752_ (_33123_, _33122_, _32081_);
  or _78753_ (_33124_, _33123_, _31051_);
  and _78754_ (_33125_, pc_inc_dir_r, _28439_);
  and _78755_ (_33126_, _33125_, _28364_);
  and _78756_ (property_invalid_inc_dir_iram, _33126_, _33124_);
  buf _78757_ (_38319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [7]);
  buf _78758_ (_38312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [0]);
  buf _78759_ (_38313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [1]);
  buf _78760_ (_38314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [2]);
  buf _78761_ (_38315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [3]);
  buf _78762_ (_38316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [4]);
  buf _78763_ (_38317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [5]);
  buf _78764_ (_38318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [6]);
  buf _78765_ (_38996_, _39040_);
  buf _78766_ (_36894_[7], _36865_[7]);
  buf _78767_ (_36895_[7], _36866_[7]);
  buf _78768_ (_36906_[7], _36865_[7]);
  buf _78769_ (_36907_[7], _36866_[7]);
  buf _78770_ (_36894_[0], _36865_[0]);
  buf _78771_ (_36894_[1], _36865_[1]);
  buf _78772_ (_36894_[2], _36865_[2]);
  buf _78773_ (_36894_[3], _36865_[3]);
  buf _78774_ (_36894_[4], _36865_[4]);
  buf _78775_ (_36894_[5], _36865_[5]);
  buf _78776_ (_36894_[6], _36865_[6]);
  buf _78777_ (_36895_[0], _36866_[0]);
  buf _78778_ (_36895_[1], _36866_[1]);
  buf _78779_ (_36895_[2], _36866_[2]);
  buf _78780_ (_36895_[3], _36866_[3]);
  buf _78781_ (_36895_[4], _36866_[4]);
  buf _78782_ (_36895_[5], _36866_[5]);
  buf _78783_ (_36895_[6], _36866_[6]);
  buf _78784_ (_36906_[0], _36865_[0]);
  buf _78785_ (_36906_[1], _36865_[1]);
  buf _78786_ (_36906_[2], _36865_[2]);
  buf _78787_ (_36906_[3], _36865_[3]);
  buf _78788_ (_36906_[4], _36865_[4]);
  buf _78789_ (_36906_[5], _36865_[5]);
  buf _78790_ (_36906_[6], _36865_[6]);
  buf _78791_ (_36907_[0], _36866_[0]);
  buf _78792_ (_36907_[1], _36866_[1]);
  buf _78793_ (_36907_[2], _36866_[2]);
  buf _78794_ (_36907_[3], _36866_[3]);
  buf _78795_ (_36907_[4], _36866_[4]);
  buf _78796_ (_36907_[5], _36866_[5]);
  buf _78797_ (_36907_[6], _36866_[6]);
  buf _78798_ (_38990_, _36880_);
  buf _78799_ (_36926_, _36880_);
  dff _78800_ (iram_op1[0], _00003_[0], clk);
  dff _78801_ (iram_op1[1], _00003_[1], clk);
  dff _78802_ (iram_op1[2], _00003_[2], clk);
  dff _78803_ (iram_op1[3], _00003_[3], clk);
  dff _78804_ (iram_op1[4], _00003_[4], clk);
  dff _78805_ (iram_op1[5], _00003_[5], clk);
  dff _78806_ (iram_op1[6], _00003_[6], clk);
  dff _78807_ (iram_op1[7], _00003_[7], clk);
  dff _78808_ (op1_out_r[0], _00005_[0], clk);
  dff _78809_ (op1_out_r[1], _00005_[1], clk);
  dff _78810_ (op1_out_r[2], _00005_[2], clk);
  dff _78811_ (op1_out_r[3], _00005_[3], clk);
  dff _78812_ (op1_out_r[4], _00005_[4], clk);
  dff _78813_ (op1_out_r[5], _00005_[5], clk);
  dff _78814_ (op1_out_r[6], _00005_[6], clk);
  dff _78815_ (op1_out_r[7], _00005_[7], clk);
  dff _78816_ (cy_reg, _00001_, clk);
  dff _78817_ (acc_reg[0], _00000_[0], clk);
  dff _78818_ (acc_reg[1], _00000_[1], clk);
  dff _78819_ (acc_reg[2], _00000_[2], clk);
  dff _78820_ (acc_reg[3], _00000_[3], clk);
  dff _78821_ (acc_reg[4], _00000_[4], clk);
  dff _78822_ (acc_reg[5], _00000_[5], clk);
  dff _78823_ (acc_reg[6], _00000_[6], clk);
  dff _78824_ (acc_reg[7], _00000_[7], clk);
  dff _78825_ (iram_op1_reg[0], _00004_[0], clk);
  dff _78826_ (iram_op1_reg[1], _00004_[1], clk);
  dff _78827_ (iram_op1_reg[2], _00004_[2], clk);
  dff _78828_ (iram_op1_reg[3], _00004_[3], clk);
  dff _78829_ (iram_op1_reg[4], _00004_[4], clk);
  dff _78830_ (iram_op1_reg[5], _00004_[5], clk);
  dff _78831_ (iram_op1_reg[6], _00004_[6], clk);
  dff _78832_ (iram_op1_reg[7], _00004_[7], clk);
  dff _78833_ (pc_change_r, _00006_, clk);
  dff _78834_ (pc_inc_acc_r, _00007_, clk);
  dff _78835_ (pc_inc_dir_r, _00008_, clk);
  dff _78836_ (first_instr, _00002_, clk);
  dff _78837_ (\oc8051_symbolic_cxrom1.regarray[0] [0], _36730_, clk);
  dff _78838_ (\oc8051_symbolic_cxrom1.regarray[0] [1], _36731_, clk);
  dff _78839_ (\oc8051_symbolic_cxrom1.regarray[0] [2], _36732_, clk);
  dff _78840_ (\oc8051_symbolic_cxrom1.regarray[0] [3], _36733_, clk);
  dff _78841_ (\oc8051_symbolic_cxrom1.regarray[0] [4], _36734_, clk);
  dff _78842_ (\oc8051_symbolic_cxrom1.regarray[0] [5], _36735_, clk);
  dff _78843_ (\oc8051_symbolic_cxrom1.regarray[0] [6], _36736_, clk);
  dff _78844_ (\oc8051_symbolic_cxrom1.regarray[0] [7], _36737_, clk);
  dff _78845_ (\oc8051_symbolic_cxrom1.regvalid [0], _36858_, clk);
  dff _78846_ (\oc8051_symbolic_cxrom1.regvalid [1], _36729_[1], clk);
  dff _78847_ (\oc8051_symbolic_cxrom1.regvalid [2], _36729_[2], clk);
  dff _78848_ (\oc8051_symbolic_cxrom1.regvalid [3], _36729_[3], clk);
  dff _78849_ (\oc8051_symbolic_cxrom1.regvalid [4], _36729_[4], clk);
  dff _78850_ (\oc8051_symbolic_cxrom1.regvalid [5], _36729_[5], clk);
  dff _78851_ (\oc8051_symbolic_cxrom1.regvalid [6], _36729_[6], clk);
  dff _78852_ (\oc8051_symbolic_cxrom1.regvalid [7], _36729_[7], clk);
  dff _78853_ (\oc8051_symbolic_cxrom1.regvalid [8], _36729_[8], clk);
  dff _78854_ (\oc8051_symbolic_cxrom1.regvalid [9], _36729_[9], clk);
  dff _78855_ (\oc8051_symbolic_cxrom1.regvalid [10], _36729_[10], clk);
  dff _78856_ (\oc8051_symbolic_cxrom1.regvalid [11], _36729_[11], clk);
  dff _78857_ (\oc8051_symbolic_cxrom1.regvalid [12], _36729_[12], clk);
  dff _78858_ (\oc8051_symbolic_cxrom1.regvalid [13], _36729_[13], clk);
  dff _78859_ (\oc8051_symbolic_cxrom1.regvalid [14], _36729_[14], clk);
  dff _78860_ (\oc8051_symbolic_cxrom1.regvalid [15], _36729_[15], clk);
  dff _78861_ (\oc8051_symbolic_cxrom1.regarray[1] [0], _36786_, clk);
  dff _78862_ (\oc8051_symbolic_cxrom1.regarray[1] [1], _36787_, clk);
  dff _78863_ (\oc8051_symbolic_cxrom1.regarray[1] [2], _36788_, clk);
  dff _78864_ (\oc8051_symbolic_cxrom1.regarray[1] [3], _36789_, clk);
  dff _78865_ (\oc8051_symbolic_cxrom1.regarray[1] [4], _36790_, clk);
  dff _78866_ (\oc8051_symbolic_cxrom1.regarray[1] [5], _36791_, clk);
  dff _78867_ (\oc8051_symbolic_cxrom1.regarray[1] [6], _36792_, clk);
  dff _78868_ (\oc8051_symbolic_cxrom1.regarray[1] [7], _36793_, clk);
  dff _78869_ (\oc8051_symbolic_cxrom1.regarray[2] [0], _36794_, clk);
  dff _78870_ (\oc8051_symbolic_cxrom1.regarray[2] [1], _36795_, clk);
  dff _78871_ (\oc8051_symbolic_cxrom1.regarray[2] [2], _36796_, clk);
  dff _78872_ (\oc8051_symbolic_cxrom1.regarray[2] [3], _36797_, clk);
  dff _78873_ (\oc8051_symbolic_cxrom1.regarray[2] [4], _36798_, clk);
  dff _78874_ (\oc8051_symbolic_cxrom1.regarray[2] [5], _36799_, clk);
  dff _78875_ (\oc8051_symbolic_cxrom1.regarray[2] [6], _36800_, clk);
  dff _78876_ (\oc8051_symbolic_cxrom1.regarray[2] [7], _36801_, clk);
  dff _78877_ (\oc8051_symbolic_cxrom1.regarray[3] [0], _36802_, clk);
  dff _78878_ (\oc8051_symbolic_cxrom1.regarray[3] [1], _36803_, clk);
  dff _78879_ (\oc8051_symbolic_cxrom1.regarray[3] [2], _36804_, clk);
  dff _78880_ (\oc8051_symbolic_cxrom1.regarray[3] [3], _36805_, clk);
  dff _78881_ (\oc8051_symbolic_cxrom1.regarray[3] [4], _36806_, clk);
  dff _78882_ (\oc8051_symbolic_cxrom1.regarray[3] [5], _36807_, clk);
  dff _78883_ (\oc8051_symbolic_cxrom1.regarray[3] [6], _36808_, clk);
  dff _78884_ (\oc8051_symbolic_cxrom1.regarray[3] [7], _36809_, clk);
  dff _78885_ (\oc8051_symbolic_cxrom1.regarray[4] [0], _36810_, clk);
  dff _78886_ (\oc8051_symbolic_cxrom1.regarray[4] [1], _36811_, clk);
  dff _78887_ (\oc8051_symbolic_cxrom1.regarray[4] [2], _36812_, clk);
  dff _78888_ (\oc8051_symbolic_cxrom1.regarray[4] [3], _36813_, clk);
  dff _78889_ (\oc8051_symbolic_cxrom1.regarray[4] [4], _36814_, clk);
  dff _78890_ (\oc8051_symbolic_cxrom1.regarray[4] [5], _36815_, clk);
  dff _78891_ (\oc8051_symbolic_cxrom1.regarray[4] [6], _36816_, clk);
  dff _78892_ (\oc8051_symbolic_cxrom1.regarray[4] [7], _36857_[7], clk);
  dff _78893_ (\oc8051_symbolic_cxrom1.regarray[5] [0], _36817_, clk);
  dff _78894_ (\oc8051_symbolic_cxrom1.regarray[5] [1], _36818_, clk);
  dff _78895_ (\oc8051_symbolic_cxrom1.regarray[5] [2], _36819_, clk);
  dff _78896_ (\oc8051_symbolic_cxrom1.regarray[5] [3], _36820_, clk);
  dff _78897_ (\oc8051_symbolic_cxrom1.regarray[5] [4], _36821_, clk);
  dff _78898_ (\oc8051_symbolic_cxrom1.regarray[5] [5], _36822_, clk);
  dff _78899_ (\oc8051_symbolic_cxrom1.regarray[5] [6], _36823_, clk);
  dff _78900_ (\oc8051_symbolic_cxrom1.regarray[5] [7], _36824_, clk);
  dff _78901_ (\oc8051_symbolic_cxrom1.regarray[6] [0], _36825_, clk);
  dff _78902_ (\oc8051_symbolic_cxrom1.regarray[6] [1], _36826_, clk);
  dff _78903_ (\oc8051_symbolic_cxrom1.regarray[6] [2], _36827_, clk);
  dff _78904_ (\oc8051_symbolic_cxrom1.regarray[6] [3], _36828_, clk);
  dff _78905_ (\oc8051_symbolic_cxrom1.regarray[6] [4], _36829_, clk);
  dff _78906_ (\oc8051_symbolic_cxrom1.regarray[6] [5], _36830_, clk);
  dff _78907_ (\oc8051_symbolic_cxrom1.regarray[6] [6], _36831_, clk);
  dff _78908_ (\oc8051_symbolic_cxrom1.regarray[6] [7], _36832_, clk);
  dff _78909_ (\oc8051_symbolic_cxrom1.regarray[7] [0], _36833_, clk);
  dff _78910_ (\oc8051_symbolic_cxrom1.regarray[7] [1], _36834_, clk);
  dff _78911_ (\oc8051_symbolic_cxrom1.regarray[7] [2], _36835_, clk);
  dff _78912_ (\oc8051_symbolic_cxrom1.regarray[7] [3], _36836_, clk);
  dff _78913_ (\oc8051_symbolic_cxrom1.regarray[7] [4], _36837_, clk);
  dff _78914_ (\oc8051_symbolic_cxrom1.regarray[7] [5], _36838_, clk);
  dff _78915_ (\oc8051_symbolic_cxrom1.regarray[7] [6], _36839_, clk);
  dff _78916_ (\oc8051_symbolic_cxrom1.regarray[7] [7], _36840_, clk);
  dff _78917_ (\oc8051_symbolic_cxrom1.regarray[8] [0], _36841_, clk);
  dff _78918_ (\oc8051_symbolic_cxrom1.regarray[8] [1], _36842_, clk);
  dff _78919_ (\oc8051_symbolic_cxrom1.regarray[8] [2], _36843_, clk);
  dff _78920_ (\oc8051_symbolic_cxrom1.regarray[8] [3], _36844_, clk);
  dff _78921_ (\oc8051_symbolic_cxrom1.regarray[8] [4], _36845_, clk);
  dff _78922_ (\oc8051_symbolic_cxrom1.regarray[8] [5], _36846_, clk);
  dff _78923_ (\oc8051_symbolic_cxrom1.regarray[8] [6], _36847_, clk);
  dff _78924_ (\oc8051_symbolic_cxrom1.regarray[8] [7], _36848_, clk);
  dff _78925_ (\oc8051_symbolic_cxrom1.regarray[9] [0], _36849_, clk);
  dff _78926_ (\oc8051_symbolic_cxrom1.regarray[9] [1], _36850_, clk);
  dff _78927_ (\oc8051_symbolic_cxrom1.regarray[9] [2], _36851_, clk);
  dff _78928_ (\oc8051_symbolic_cxrom1.regarray[9] [3], _36852_, clk);
  dff _78929_ (\oc8051_symbolic_cxrom1.regarray[9] [4], _36853_, clk);
  dff _78930_ (\oc8051_symbolic_cxrom1.regarray[9] [5], _36854_, clk);
  dff _78931_ (\oc8051_symbolic_cxrom1.regarray[9] [6], _36855_, clk);
  dff _78932_ (\oc8051_symbolic_cxrom1.regarray[9] [7], _36856_, clk);
  dff _78933_ (\oc8051_symbolic_cxrom1.regarray[10] [0], _36738_, clk);
  dff _78934_ (\oc8051_symbolic_cxrom1.regarray[10] [1], _36739_, clk);
  dff _78935_ (\oc8051_symbolic_cxrom1.regarray[10] [2], _36740_, clk);
  dff _78936_ (\oc8051_symbolic_cxrom1.regarray[10] [3], _36741_, clk);
  dff _78937_ (\oc8051_symbolic_cxrom1.regarray[10] [4], _36742_, clk);
  dff _78938_ (\oc8051_symbolic_cxrom1.regarray[10] [5], _36743_, clk);
  dff _78939_ (\oc8051_symbolic_cxrom1.regarray[10] [6], _36744_, clk);
  dff _78940_ (\oc8051_symbolic_cxrom1.regarray[10] [7], _36745_, clk);
  dff _78941_ (\oc8051_symbolic_cxrom1.regarray[11] [0], _36746_, clk);
  dff _78942_ (\oc8051_symbolic_cxrom1.regarray[11] [1], _36747_, clk);
  dff _78943_ (\oc8051_symbolic_cxrom1.regarray[11] [2], _36748_, clk);
  dff _78944_ (\oc8051_symbolic_cxrom1.regarray[11] [3], _36749_, clk);
  dff _78945_ (\oc8051_symbolic_cxrom1.regarray[11] [4], _36750_, clk);
  dff _78946_ (\oc8051_symbolic_cxrom1.regarray[11] [5], _36751_, clk);
  dff _78947_ (\oc8051_symbolic_cxrom1.regarray[11] [6], _36752_, clk);
  dff _78948_ (\oc8051_symbolic_cxrom1.regarray[11] [7], _36753_, clk);
  dff _78949_ (\oc8051_symbolic_cxrom1.regarray[12] [0], _36754_, clk);
  dff _78950_ (\oc8051_symbolic_cxrom1.regarray[12] [1], _36755_, clk);
  dff _78951_ (\oc8051_symbolic_cxrom1.regarray[12] [2], _36756_, clk);
  dff _78952_ (\oc8051_symbolic_cxrom1.regarray[12] [3], _36757_, clk);
  dff _78953_ (\oc8051_symbolic_cxrom1.regarray[12] [4], _36758_, clk);
  dff _78954_ (\oc8051_symbolic_cxrom1.regarray[12] [5], _36759_, clk);
  dff _78955_ (\oc8051_symbolic_cxrom1.regarray[12] [6], _36760_, clk);
  dff _78956_ (\oc8051_symbolic_cxrom1.regarray[12] [7], _36761_, clk);
  dff _78957_ (\oc8051_symbolic_cxrom1.regarray[13] [0], _36762_, clk);
  dff _78958_ (\oc8051_symbolic_cxrom1.regarray[13] [1], _36763_, clk);
  dff _78959_ (\oc8051_symbolic_cxrom1.regarray[13] [2], _36764_, clk);
  dff _78960_ (\oc8051_symbolic_cxrom1.regarray[13] [3], _36765_, clk);
  dff _78961_ (\oc8051_symbolic_cxrom1.regarray[13] [4], _36766_, clk);
  dff _78962_ (\oc8051_symbolic_cxrom1.regarray[13] [5], _36767_, clk);
  dff _78963_ (\oc8051_symbolic_cxrom1.regarray[13] [6], _36768_, clk);
  dff _78964_ (\oc8051_symbolic_cxrom1.regarray[13] [7], _36769_, clk);
  dff _78965_ (\oc8051_symbolic_cxrom1.regarray[14] [0], _36770_, clk);
  dff _78966_ (\oc8051_symbolic_cxrom1.regarray[14] [1], _36771_, clk);
  dff _78967_ (\oc8051_symbolic_cxrom1.regarray[14] [2], _36772_, clk);
  dff _78968_ (\oc8051_symbolic_cxrom1.regarray[14] [3], _36773_, clk);
  dff _78969_ (\oc8051_symbolic_cxrom1.regarray[14] [4], _36774_, clk);
  dff _78970_ (\oc8051_symbolic_cxrom1.regarray[14] [5], _36775_, clk);
  dff _78971_ (\oc8051_symbolic_cxrom1.regarray[14] [6], _36776_, clk);
  dff _78972_ (\oc8051_symbolic_cxrom1.regarray[14] [7], _36777_, clk);
  dff _78973_ (\oc8051_symbolic_cxrom1.regarray[15] [0], _36778_, clk);
  dff _78974_ (\oc8051_symbolic_cxrom1.regarray[15] [1], _36779_, clk);
  dff _78975_ (\oc8051_symbolic_cxrom1.regarray[15] [2], _36780_, clk);
  dff _78976_ (\oc8051_symbolic_cxrom1.regarray[15] [3], _36781_, clk);
  dff _78977_ (\oc8051_symbolic_cxrom1.regarray[15] [4], _36782_, clk);
  dff _78978_ (\oc8051_symbolic_cxrom1.regarray[15] [5], _36783_, clk);
  dff _78979_ (\oc8051_symbolic_cxrom1.regarray[15] [6], _36784_, clk);
  dff _78980_ (\oc8051_symbolic_cxrom1.regarray[15] [7], _36785_, clk);
  dff _78981_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _36860_[0], clk);
  dff _78982_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _36860_[1], clk);
  dff _78983_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _36860_[2], clk);
  dff _78984_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _36860_[3], clk);
  dff _78985_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _36860_[4], clk);
  dff _78986_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _36860_[5], clk);
  dff _78987_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _36859_[0], clk);
  dff _78988_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _36859_[1], clk);
  dff _78989_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _36861_[0], clk);
  dff _78990_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _36861_[1], clk);
  dff _78991_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _36861_[2], clk);
  dff _78992_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _36861_[3], clk);
  dff _78993_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _36861_[4], clk);
  dff _78994_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _36861_[5], clk);
  dff _78995_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _36861_[6], clk);
  dff _78996_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _36861_[7], clk);
  dff _78997_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _36862_[0], clk);
  dff _78998_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _36862_[1], clk);
  dff _78999_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _36863_[0], clk);
  dff _79000_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _36863_[1], clk);
  dff _79001_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _36863_[2], clk);
  dff _79002_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _36863_[3], clk);
  dff _79003_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _36863_[4], clk);
  dff _79004_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _36863_[5], clk);
  dff _79005_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _36863_[6], clk);
  dff _79006_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _36863_[7], clk);
  dff _79007_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _36863_[8], clk);
  dff _79008_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _36863_[9], clk);
  dff _79009_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _36863_[10], clk);
  dff _79010_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _36863_[11], clk);
  dff _79011_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _36863_[12], clk);
  dff _79012_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _36863_[13], clk);
  dff _79013_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _36863_[14], clk);
  dff _79014_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _36863_[15], clk);
  dff _79015_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _36864_[0], clk);
  dff _79016_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _36864_[1], clk);
  dff _79017_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _36864_[2], clk);
  dff _79018_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _36864_[3], clk);
  dff _79019_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _36864_[4], clk);
  dff _79020_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _36864_[5], clk);
  dff _79021_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _36864_[6], clk);
  dff _79022_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _36864_[7], clk);
  dff _79023_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _36865_[0], clk);
  dff _79024_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _36865_[1], clk);
  dff _79025_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _36865_[2], clk);
  dff _79026_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _36865_[3], clk);
  dff _79027_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _36865_[4], clk);
  dff _79028_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _36865_[5], clk);
  dff _79029_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _36865_[6], clk);
  dff _79030_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _36865_[7], clk);
  dff _79031_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _36866_[0], clk);
  dff _79032_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _36866_[1], clk);
  dff _79033_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _36866_[2], clk);
  dff _79034_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _36866_[3], clk);
  dff _79035_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _36866_[4], clk);
  dff _79036_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _36866_[5], clk);
  dff _79037_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _36866_[6], clk);
  dff _79038_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _36866_[7], clk);
  dff _79039_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _36867_[0], clk);
  dff _79040_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _36867_[1], clk);
  dff _79041_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _36867_[2], clk);
  dff _79042_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _36868_[0], clk);
  dff _79043_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _36868_[1], clk);
  dff _79044_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _36868_[2], clk);
  dff _79045_ (\oc8051_top_1.oc8051_decoder1.state [0], _36869_[0], clk);
  dff _79046_ (\oc8051_top_1.oc8051_decoder1.state [1], _36869_[1], clk);
  dff _79047_ (\oc8051_top_1.oc8051_decoder1.op [0], _36870_[0], clk);
  dff _79048_ (\oc8051_top_1.oc8051_decoder1.op [1], _36870_[1], clk);
  dff _79049_ (\oc8051_top_1.oc8051_decoder1.op [2], _36870_[2], clk);
  dff _79050_ (\oc8051_top_1.oc8051_decoder1.op [3], _36870_[3], clk);
  dff _79051_ (\oc8051_top_1.oc8051_decoder1.op [4], _36870_[4], clk);
  dff _79052_ (\oc8051_top_1.oc8051_decoder1.op [5], _36870_[5], clk);
  dff _79053_ (\oc8051_top_1.oc8051_decoder1.op [6], _36870_[6], clk);
  dff _79054_ (\oc8051_top_1.oc8051_decoder1.op [7], _36870_[7], clk);
  dff _79055_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _36871_, clk);
  dff _79056_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _36872_[0], clk);
  dff _79057_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _36872_[1], clk);
  dff _79058_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _36873_[0], clk);
  dff _79059_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _36873_[1], clk);
  dff _79060_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _36874_[0], clk);
  dff _79061_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _36874_[1], clk);
  dff _79062_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _36874_[2], clk);
  dff _79063_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _36875_[0], clk);
  dff _79064_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _36875_[1], clk);
  dff _79065_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _36875_[2], clk);
  dff _79066_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _36876_[0], clk);
  dff _79067_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _36876_[1], clk);
  dff _79068_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _36877_[0], clk);
  dff _79069_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _36877_[1], clk);
  dff _79070_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _36877_[2], clk);
  dff _79071_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _36877_[3], clk);
  dff _79072_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _36878_[0], clk);
  dff _79073_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _36878_[1], clk);
  dff _79074_ (\oc8051_top_1.oc8051_decoder1.wr , _36879_, clk);
  dff _79075_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _36880_, clk);
  dff _79076_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _36881_[0], clk);
  dff _79077_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _36881_[1], clk);
  dff _79078_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _36881_[2], clk);
  dff _79079_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _36881_[3], clk);
  dff _79080_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _36881_[4], clk);
  dff _79081_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _36881_[5], clk);
  dff _79082_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _36881_[6], clk);
  dff _79083_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _36881_[7], clk);
  dff _79084_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _36882_[0], clk);
  dff _79085_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _36882_[1], clk);
  dff _79086_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _36882_[2], clk);
  dff _79087_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _36882_[3], clk);
  dff _79088_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _36882_[4], clk);
  dff _79089_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _36882_[5], clk);
  dff _79090_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _36882_[6], clk);
  dff _79091_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _36882_[7], clk);
  dff _79092_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _36883_[0], clk);
  dff _79093_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _36883_[1], clk);
  dff _79094_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _36883_[2], clk);
  dff _79095_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _36883_[3], clk);
  dff _79096_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _36883_[4], clk);
  dff _79097_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _36883_[5], clk);
  dff _79098_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _36883_[6], clk);
  dff _79099_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _36883_[7], clk);
  dff _79100_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _36884_[0], clk);
  dff _79101_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _36884_[1], clk);
  dff _79102_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _36884_[2], clk);
  dff _79103_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _36884_[3], clk);
  dff _79104_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _36884_[4], clk);
  dff _79105_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _36884_[5], clk);
  dff _79106_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _36884_[6], clk);
  dff _79107_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _36884_[7], clk);
  dff _79108_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _36885_[0], clk);
  dff _79109_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _36885_[1], clk);
  dff _79110_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _36885_[2], clk);
  dff _79111_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _36885_[3], clk);
  dff _79112_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _36885_[4], clk);
  dff _79113_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _36885_[5], clk);
  dff _79114_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _36885_[6], clk);
  dff _79115_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _36885_[7], clk);
  dff _79116_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _36886_[0], clk);
  dff _79117_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _36886_[1], clk);
  dff _79118_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _36886_[2], clk);
  dff _79119_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _36886_[3], clk);
  dff _79120_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _36886_[4], clk);
  dff _79121_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _36886_[5], clk);
  dff _79122_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _36886_[6], clk);
  dff _79123_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _36886_[7], clk);
  dff _79124_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _36887_[0], clk);
  dff _79125_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _36887_[1], clk);
  dff _79126_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _36887_[2], clk);
  dff _79127_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _36887_[3], clk);
  dff _79128_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _36887_[4], clk);
  dff _79129_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _36887_[5], clk);
  dff _79130_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _36887_[6], clk);
  dff _79131_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _36887_[7], clk);
  dff _79132_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _36888_[0], clk);
  dff _79133_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _36888_[1], clk);
  dff _79134_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _36888_[2], clk);
  dff _79135_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _36888_[3], clk);
  dff _79136_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _36888_[4], clk);
  dff _79137_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _36888_[5], clk);
  dff _79138_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _36888_[6], clk);
  dff _79139_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _36888_[7], clk);
  dff _79140_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _36892_[0], clk);
  dff _79141_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _36892_[1], clk);
  dff _79142_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _36892_[2], clk);
  dff _79143_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _36892_[3], clk);
  dff _79144_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _36892_[4], clk);
  dff _79145_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _36889_[0], clk);
  dff _79146_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _36889_[1], clk);
  dff _79147_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _36889_[2], clk);
  dff _79148_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _36889_[3], clk);
  dff _79149_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _36889_[4], clk);
  dff _79150_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _36889_[5], clk);
  dff _79151_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _36889_[6], clk);
  dff _79152_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _36889_[7], clk);
  dff _79153_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _36889_[8], clk);
  dff _79154_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _36889_[9], clk);
  dff _79155_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _36889_[10], clk);
  dff _79156_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _36889_[11], clk);
  dff _79157_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _36889_[12], clk);
  dff _79158_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _36889_[13], clk);
  dff _79159_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _36889_[14], clk);
  dff _79160_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _36889_[15], clk);
  dff _79161_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _36890_[0], clk);
  dff _79162_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _36890_[1], clk);
  dff _79163_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _36890_[2], clk);
  dff _79164_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _36890_[3], clk);
  dff _79165_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _36890_[4], clk);
  dff _79166_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _36890_[5], clk);
  dff _79167_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _36890_[6], clk);
  dff _79168_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _36890_[7], clk);
  dff _79169_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _36890_[8], clk);
  dff _79170_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _36890_[9], clk);
  dff _79171_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _36890_[10], clk);
  dff _79172_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _36890_[11], clk);
  dff _79173_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _36890_[12], clk);
  dff _79174_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _36890_[13], clk);
  dff _79175_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _36890_[14], clk);
  dff _79176_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _36890_[15], clk);
  dff _79177_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _36913_[0], clk);
  dff _79178_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _36913_[1], clk);
  dff _79179_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _36913_[2], clk);
  dff _79180_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _36913_[3], clk);
  dff _79181_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _36913_[4], clk);
  dff _79182_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _36913_[5], clk);
  dff _79183_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _36913_[6], clk);
  dff _79184_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _36913_[7], clk);
  dff _79185_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _36913_[8], clk);
  dff _79186_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _36913_[9], clk);
  dff _79187_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _36913_[10], clk);
  dff _79188_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _36913_[11], clk);
  dff _79189_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _36913_[12], clk);
  dff _79190_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _36913_[13], clk);
  dff _79191_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _36913_[14], clk);
  dff _79192_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _36913_[15], clk);
  dff _79193_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _36913_[16], clk);
  dff _79194_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _36913_[17], clk);
  dff _79195_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _36913_[18], clk);
  dff _79196_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _36913_[19], clk);
  dff _79197_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _36913_[20], clk);
  dff _79198_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _36913_[21], clk);
  dff _79199_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _36913_[22], clk);
  dff _79200_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _36913_[23], clk);
  dff _79201_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _36913_[24], clk);
  dff _79202_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _36913_[25], clk);
  dff _79203_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _36913_[26], clk);
  dff _79204_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _36913_[27], clk);
  dff _79205_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _36913_[28], clk);
  dff _79206_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _36913_[29], clk);
  dff _79207_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _36913_[30], clk);
  dff _79208_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _36913_[31], clk);
  dff _79209_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _36891_, clk);
  dff _79210_ (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0, clk);
  dff _79211_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _36893_[0], clk);
  dff _79212_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _36893_[1], clk);
  dff _79213_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _36893_[2], clk);
  dff _79214_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _36893_[3], clk);
  dff _79215_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _36893_[4], clk);
  dff _79216_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _36893_[5], clk);
  dff _79217_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _36893_[6], clk);
  dff _79218_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _36893_[7], clk);
  dff _79219_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _36894_[0], clk);
  dff _79220_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _36894_[1], clk);
  dff _79221_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _36894_[2], clk);
  dff _79222_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _36894_[3], clk);
  dff _79223_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _36894_[4], clk);
  dff _79224_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _36894_[5], clk);
  dff _79225_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _36894_[6], clk);
  dff _79226_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _36894_[7], clk);
  dff _79227_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _36895_[0], clk);
  dff _79228_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _36895_[1], clk);
  dff _79229_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _36895_[2], clk);
  dff _79230_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _36895_[3], clk);
  dff _79231_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _36895_[4], clk);
  dff _79232_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _36895_[5], clk);
  dff _79233_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _36895_[6], clk);
  dff _79234_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _36895_[7], clk);
  dff _79235_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _36896_, clk);
  dff _79236_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _36897_, clk);
  dff _79237_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _36898_[0], clk);
  dff _79238_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _36898_[1], clk);
  dff _79239_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _36898_[2], clk);
  dff _79240_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _36898_[3], clk);
  dff _79241_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _36898_[4], clk);
  dff _79242_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _36898_[5], clk);
  dff _79243_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _36898_[6], clk);
  dff _79244_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _36898_[7], clk);
  dff _79245_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _36899_[0], clk);
  dff _79246_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _36899_[1], clk);
  dff _79247_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _36899_[2], clk);
  dff _79248_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _36899_[3], clk);
  dff _79249_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _36899_[4], clk);
  dff _79250_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _36899_[5], clk);
  dff _79251_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _36899_[6], clk);
  dff _79252_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _36899_[7], clk);
  dff _79253_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _36899_[8], clk);
  dff _79254_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _36899_[9], clk);
  dff _79255_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _36899_[10], clk);
  dff _79256_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _36899_[11], clk);
  dff _79257_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _36899_[12], clk);
  dff _79258_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _36899_[13], clk);
  dff _79259_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _36899_[14], clk);
  dff _79260_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _36899_[15], clk);
  dff _79261_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _36900_[0], clk);
  dff _79262_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _36900_[1], clk);
  dff _79263_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _36900_[2], clk);
  dff _79264_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _36900_[3], clk);
  dff _79265_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _36900_[4], clk);
  dff _79266_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _36900_[5], clk);
  dff _79267_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _36900_[6], clk);
  dff _79268_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _36900_[7], clk);
  dff _79269_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _36900_[8], clk);
  dff _79270_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _36900_[9], clk);
  dff _79271_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _36900_[10], clk);
  dff _79272_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _36900_[11], clk);
  dff _79273_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _36900_[12], clk);
  dff _79274_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _36900_[13], clk);
  dff _79275_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _36900_[14], clk);
  dff _79276_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _36900_[15], clk);
  dff _79277_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _36901_, clk);
  dff _79278_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _36903_, clk);
  dff _79279_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _36902_, clk);
  dff _79280_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _36904_[0], clk);
  dff _79281_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _36904_[1], clk);
  dff _79282_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _36904_[2], clk);
  dff _79283_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _36904_[3], clk);
  dff _79284_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _36904_[4], clk);
  dff _79285_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _36904_[5], clk);
  dff _79286_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _36904_[6], clk);
  dff _79287_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _36904_[7], clk);
  dff _79288_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _36905_[0], clk);
  dff _79289_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _36905_[1], clk);
  dff _79290_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _36905_[2], clk);
  dff _79291_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _36906_[0], clk);
  dff _79292_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _36906_[1], clk);
  dff _79293_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _36906_[2], clk);
  dff _79294_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _36906_[3], clk);
  dff _79295_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _36906_[4], clk);
  dff _79296_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _36906_[5], clk);
  dff _79297_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _36906_[6], clk);
  dff _79298_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _36906_[7], clk);
  dff _79299_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _36907_[0], clk);
  dff _79300_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _36907_[1], clk);
  dff _79301_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _36907_[2], clk);
  dff _79302_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _36907_[3], clk);
  dff _79303_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _36907_[4], clk);
  dff _79304_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _36907_[5], clk);
  dff _79305_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _36907_[6], clk);
  dff _79306_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _36907_[7], clk);
  dff _79307_ (\oc8051_top_1.oc8051_memory_interface1.reti , _36908_, clk);
  dff _79308_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _36909_[0], clk);
  dff _79309_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _36909_[1], clk);
  dff _79310_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _36909_[2], clk);
  dff _79311_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _36909_[3], clk);
  dff _79312_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _36909_[4], clk);
  dff _79313_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _36909_[5], clk);
  dff _79314_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _36909_[6], clk);
  dff _79315_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _36909_[7], clk);
  dff _79316_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _36910_, clk);
  dff _79317_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _36911_, clk);
  dff _79318_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _36912_[0], clk);
  dff _79319_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _36912_[1], clk);
  dff _79320_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _36912_[2], clk);
  dff _79321_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _36912_[3], clk);
  dff _79322_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _36914_[0], clk);
  dff _79323_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _36914_[1], clk);
  dff _79324_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _36914_[2], clk);
  dff _79325_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _36914_[3], clk);
  dff _79326_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _36914_[4], clk);
  dff _79327_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _36914_[5], clk);
  dff _79328_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _36914_[6], clk);
  dff _79329_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _36914_[7], clk);
  dff _79330_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _36914_[8], clk);
  dff _79331_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _36914_[9], clk);
  dff _79332_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _36914_[10], clk);
  dff _79333_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _36914_[11], clk);
  dff _79334_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _36914_[12], clk);
  dff _79335_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _36914_[13], clk);
  dff _79336_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _36914_[14], clk);
  dff _79337_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _36914_[15], clk);
  dff _79338_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _36914_[16], clk);
  dff _79339_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _36914_[17], clk);
  dff _79340_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _36914_[18], clk);
  dff _79341_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _36914_[19], clk);
  dff _79342_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _36914_[20], clk);
  dff _79343_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _36914_[21], clk);
  dff _79344_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _36914_[22], clk);
  dff _79345_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _36914_[23], clk);
  dff _79346_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _36914_[24], clk);
  dff _79347_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _36914_[25], clk);
  dff _79348_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _36914_[26], clk);
  dff _79349_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _36914_[27], clk);
  dff _79350_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _36914_[28], clk);
  dff _79351_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _36914_[29], clk);
  dff _79352_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _36914_[30], clk);
  dff _79353_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _36914_[31], clk);
  dff _79354_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _36915_[0], clk);
  dff _79355_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _36915_[1], clk);
  dff _79356_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _36915_[2], clk);
  dff _79357_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _36915_[3], clk);
  dff _79358_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _36915_[4], clk);
  dff _79359_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _36915_[5], clk);
  dff _79360_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _36915_[6], clk);
  dff _79361_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _36915_[7], clk);
  dff _79362_ (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _36916_, clk);
  dff _79363_ (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _36917_, clk);
  dff _79364_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _36918_[0], clk);
  dff _79365_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _36918_[1], clk);
  dff _79366_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _36918_[2], clk);
  dff _79367_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _36918_[3], clk);
  dff _79368_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _36918_[4], clk);
  dff _79369_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _36918_[5], clk);
  dff _79370_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _36918_[6], clk);
  dff _79371_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _36918_[7], clk);
  dff _79372_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _36918_[8], clk);
  dff _79373_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _36918_[9], clk);
  dff _79374_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _36918_[10], clk);
  dff _79375_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _36918_[11], clk);
  dff _79376_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _36918_[12], clk);
  dff _79377_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _36918_[13], clk);
  dff _79378_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _36918_[14], clk);
  dff _79379_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _36918_[15], clk);
  dff _79380_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _36919_, clk);
  dff _79381_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _36920_, clk);
  dff _79382_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _36921_, clk);
  dff _79383_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _36922_[0], clk);
  dff _79384_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _36922_[1], clk);
  dff _79385_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _36922_[2], clk);
  dff _79386_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _36922_[3], clk);
  dff _79387_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _36922_[4], clk);
  dff _79388_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _36922_[5], clk);
  dff _79389_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _36922_[6], clk);
  dff _79390_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _36922_[7], clk);
  dff _79391_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _36922_[8], clk);
  dff _79392_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _36922_[9], clk);
  dff _79393_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _36922_[10], clk);
  dff _79394_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _36922_[11], clk);
  dff _79395_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _36922_[12], clk);
  dff _79396_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _36922_[13], clk);
  dff _79397_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _36922_[14], clk);
  dff _79398_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _36922_[15], clk);
  dff _79399_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _36923_, clk);
  dff _79400_ (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _36924_, clk);
  dff _79401_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _36925_[0], clk);
  dff _79402_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _36925_[1], clk);
  dff _79403_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _36925_[2], clk);
  dff _79404_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _36925_[3], clk);
  dff _79405_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _36925_[4], clk);
  dff _79406_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _36925_[5], clk);
  dff _79407_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _36925_[6], clk);
  dff _79408_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _36925_[7], clk);
  dff _79409_ (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _36926_, clk);
  dff _79410_ (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _36927_[0], clk);
  dff _79411_ (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _36927_[1], clk);
  dff _79412_ (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _36927_[2], clk);
  dff _79413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _37136_, clk);
  dff _79414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _37137_, clk);
  dff _79415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _37138_, clk);
  dff _79416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _37139_, clk);
  dff _79417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _37140_, clk);
  dff _79418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _37141_, clk);
  dff _79419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _37142_, clk);
  dff _79420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _37143_, clk);
  dff _79421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _37128_, clk);
  dff _79422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _37129_, clk);
  dff _79423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _37130_, clk);
  dff _79424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _37131_, clk);
  dff _79425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _37132_, clk);
  dff _79426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _37133_, clk);
  dff _79427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _37134_, clk);
  dff _79428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _37135_, clk);
  dff _79429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _37120_, clk);
  dff _79430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _37121_, clk);
  dff _79431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _37122_, clk);
  dff _79432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _37123_, clk);
  dff _79433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _37124_, clk);
  dff _79434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _37125_, clk);
  dff _79435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _37126_, clk);
  dff _79436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _37127_, clk);
  dff _79437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _37112_, clk);
  dff _79438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _37113_, clk);
  dff _79439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _37114_, clk);
  dff _79440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _37115_, clk);
  dff _79441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _37116_, clk);
  dff _79442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _37117_, clk);
  dff _79443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _37118_, clk);
  dff _79444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _37119_, clk);
  dff _79445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _37096_, clk);
  dff _79446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _37097_, clk);
  dff _79447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _37098_, clk);
  dff _79448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _37099_, clk);
  dff _79449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _37100_, clk);
  dff _79450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _37101_, clk);
  dff _79451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _37102_, clk);
  dff _79452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _37103_, clk);
  dff _79453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _37088_, clk);
  dff _79454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _37089_, clk);
  dff _79455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _37090_, clk);
  dff _79456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _37091_, clk);
  dff _79457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _37092_, clk);
  dff _79458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _37093_, clk);
  dff _79459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _37094_, clk);
  dff _79460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _37095_, clk);
  dff _79461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _37080_, clk);
  dff _79462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _37081_, clk);
  dff _79463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _37082_, clk);
  dff _79464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _37083_, clk);
  dff _79465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _37084_, clk);
  dff _79466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _37085_, clk);
  dff _79467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _37086_, clk);
  dff _79468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _37087_, clk);
  dff _79469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _37072_, clk);
  dff _79470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _37073_, clk);
  dff _79471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _37074_, clk);
  dff _79472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _37075_, clk);
  dff _79473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _37076_, clk);
  dff _79474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _37077_, clk);
  dff _79475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _37078_, clk);
  dff _79476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _37079_, clk);
  dff _79477_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _37184_, clk);
  dff _79478_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _37185_, clk);
  dff _79479_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _37186_, clk);
  dff _79480_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _37187_, clk);
  dff _79481_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _37188_, clk);
  dff _79482_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _37189_, clk);
  dff _79483_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _37190_, clk);
  dff _79484_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _37191_, clk);
  dff _79485_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _37064_, clk);
  dff _79486_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _37065_, clk);
  dff _79487_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _37066_, clk);
  dff _79488_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _37067_, clk);
  dff _79489_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _37068_, clk);
  dff _79490_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _37069_, clk);
  dff _79491_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _37070_, clk);
  dff _79492_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _37071_, clk);
  dff _79493_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _37056_, clk);
  dff _79494_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _37057_, clk);
  dff _79495_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _37058_, clk);
  dff _79496_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _37059_, clk);
  dff _79497_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _37060_, clk);
  dff _79498_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _37061_, clk);
  dff _79499_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _37062_, clk);
  dff _79500_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _37063_, clk);
  dff _79501_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _37048_, clk);
  dff _79502_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _37049_, clk);
  dff _79503_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _37050_, clk);
  dff _79504_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _37051_, clk);
  dff _79505_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _37052_, clk);
  dff _79506_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _37053_, clk);
  dff _79507_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _37054_, clk);
  dff _79508_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _37055_, clk);
  dff _79509_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _37040_, clk);
  dff _79510_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _37041_, clk);
  dff _79511_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _37042_, clk);
  dff _79512_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _37043_, clk);
  dff _79513_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _37044_, clk);
  dff _79514_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _37045_, clk);
  dff _79515_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _37046_, clk);
  dff _79516_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _37047_, clk);
  dff _79517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _37032_, clk);
  dff _79518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _37033_, clk);
  dff _79519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _37034_, clk);
  dff _79520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _37035_, clk);
  dff _79521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _37036_, clk);
  dff _79522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _37037_, clk);
  dff _79523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _37038_, clk);
  dff _79524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _37039_, clk);
  dff _79525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _37024_, clk);
  dff _79526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _37025_, clk);
  dff _79527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _37026_, clk);
  dff _79528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _37027_, clk);
  dff _79529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _37028_, clk);
  dff _79530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _37029_, clk);
  dff _79531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _37030_, clk);
  dff _79532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _37031_, clk);
  dff _79533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _37008_, clk);
  dff _79534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _37009_, clk);
  dff _79535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _37010_, clk);
  dff _79536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _37011_, clk);
  dff _79537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _37012_, clk);
  dff _79538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _37013_, clk);
  dff _79539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _37014_, clk);
  dff _79540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _37015_, clk);
  dff _79541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _37000_, clk);
  dff _79542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _37001_, clk);
  dff _79543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _37002_, clk);
  dff _79544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _37003_, clk);
  dff _79545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _37004_, clk);
  dff _79546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _37005_, clk);
  dff _79547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _37006_, clk);
  dff _79548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _37007_, clk);
  dff _79549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _37200_, clk);
  dff _79550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _37201_, clk);
  dff _79551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _37202_, clk);
  dff _79552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _37203_, clk);
  dff _79553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _37204_, clk);
  dff _79554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _37205_, clk);
  dff _79555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _37206_, clk);
  dff _79556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _37207_, clk);
  dff _79557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _37272_, clk);
  dff _79558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _37273_, clk);
  dff _79559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _37274_, clk);
  dff _79560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _37275_, clk);
  dff _79561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _37276_, clk);
  dff _79562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _37277_, clk);
  dff _79563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _37278_, clk);
  dff _79564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _37279_, clk);
  dff _79565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _37264_, clk);
  dff _79566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _37265_, clk);
  dff _79567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _37266_, clk);
  dff _79568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _37267_, clk);
  dff _79569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _37268_, clk);
  dff _79570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _37269_, clk);
  dff _79571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _37270_, clk);
  dff _79572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _37271_, clk);
  dff _79573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _37256_, clk);
  dff _79574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _37257_, clk);
  dff _79575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _37258_, clk);
  dff _79576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _37259_, clk);
  dff _79577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _37260_, clk);
  dff _79578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _37261_, clk);
  dff _79579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _37262_, clk);
  dff _79580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _37263_, clk);
  dff _79581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _37480_, clk);
  dff _79582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _37481_, clk);
  dff _79583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _37482_, clk);
  dff _79584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _37483_, clk);
  dff _79585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _37484_, clk);
  dff _79586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _37485_, clk);
  dff _79587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _37486_, clk);
  dff _79588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _37487_, clk);
  dff _79589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _37472_, clk);
  dff _79590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _37473_, clk);
  dff _79591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _37474_, clk);
  dff _79592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _37475_, clk);
  dff _79593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _37476_, clk);
  dff _79594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _37477_, clk);
  dff _79595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _37478_, clk);
  dff _79596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _37479_, clk);
  dff _79597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _37464_, clk);
  dff _79598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _37465_, clk);
  dff _79599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _37466_, clk);
  dff _79600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _37467_, clk);
  dff _79601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _37468_, clk);
  dff _79602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _37469_, clk);
  dff _79603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _37470_, clk);
  dff _79604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _37471_, clk);
  dff _79605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _37448_, clk);
  dff _79606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _37449_, clk);
  dff _79607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _37450_, clk);
  dff _79608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _37451_, clk);
  dff _79609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _37452_, clk);
  dff _79610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _37453_, clk);
  dff _79611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _37454_, clk);
  dff _79612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _37455_, clk);
  dff _79613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _37440_, clk);
  dff _79614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _37441_, clk);
  dff _79615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _37442_, clk);
  dff _79616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _37443_, clk);
  dff _79617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _37444_, clk);
  dff _79618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _37445_, clk);
  dff _79619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _37446_, clk);
  dff _79620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _37447_, clk);
  dff _79621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _37432_, clk);
  dff _79622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _37433_, clk);
  dff _79623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _37434_, clk);
  dff _79624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _37435_, clk);
  dff _79625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _37436_, clk);
  dff _79626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _37437_, clk);
  dff _79627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _37438_, clk);
  dff _79628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _37439_, clk);
  dff _79629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _37424_, clk);
  dff _79630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _37425_, clk);
  dff _79631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _37426_, clk);
  dff _79632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _37427_, clk);
  dff _79633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _37428_, clk);
  dff _79634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _37429_, clk);
  dff _79635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _37430_, clk);
  dff _79636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _37431_, clk);
  dff _79637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _37416_, clk);
  dff _79638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _37417_, clk);
  dff _79639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _37418_, clk);
  dff _79640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _37419_, clk);
  dff _79641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _37420_, clk);
  dff _79642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _37421_, clk);
  dff _79643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _37422_, clk);
  dff _79644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _37423_, clk);
  dff _79645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _37408_, clk);
  dff _79646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _37409_, clk);
  dff _79647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _37410_, clk);
  dff _79648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _37411_, clk);
  dff _79649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _37412_, clk);
  dff _79650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _37413_, clk);
  dff _79651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _37414_, clk);
  dff _79652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _37415_, clk);
  dff _79653_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _37400_, clk);
  dff _79654_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _37401_, clk);
  dff _79655_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _37402_, clk);
  dff _79656_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _37403_, clk);
  dff _79657_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _37404_, clk);
  dff _79658_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _37405_, clk);
  dff _79659_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _37406_, clk);
  dff _79660_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _37407_, clk);
  dff _79661_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _37928_, clk);
  dff _79662_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _37929_, clk);
  dff _79663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _37930_, clk);
  dff _79664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _37931_, clk);
  dff _79665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _37932_, clk);
  dff _79666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _37933_, clk);
  dff _79667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _37934_, clk);
  dff _79668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _37935_, clk);
  dff _79669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _37920_, clk);
  dff _79670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _37921_, clk);
  dff _79671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _37922_, clk);
  dff _79672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _37923_, clk);
  dff _79673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _37924_, clk);
  dff _79674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _37925_, clk);
  dff _79675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _37926_, clk);
  dff _79676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _37927_, clk);
  dff _79677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _37912_, clk);
  dff _79678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _37913_, clk);
  dff _79679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _37914_, clk);
  dff _79680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _37915_, clk);
  dff _79681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _37916_, clk);
  dff _79682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _37917_, clk);
  dff _79683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _37918_, clk);
  dff _79684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _37919_, clk);
  dff _79685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _37896_, clk);
  dff _79686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _37897_, clk);
  dff _79687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _37898_, clk);
  dff _79688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _37899_, clk);
  dff _79689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _37900_, clk);
  dff _79690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _37901_, clk);
  dff _79691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _37902_, clk);
  dff _79692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _37903_, clk);
  dff _79693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _37888_, clk);
  dff _79694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _37889_, clk);
  dff _79695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _37890_, clk);
  dff _79696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _37891_, clk);
  dff _79697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _37892_, clk);
  dff _79698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _37893_, clk);
  dff _79699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _37894_, clk);
  dff _79700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _37895_, clk);
  dff _79701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _37880_, clk);
  dff _79702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _37881_, clk);
  dff _79703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _37882_, clk);
  dff _79704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _37883_, clk);
  dff _79705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _37884_, clk);
  dff _79706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _37885_, clk);
  dff _79707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _37886_, clk);
  dff _79708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _37887_, clk);
  dff _79709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _37872_, clk);
  dff _79710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _37873_, clk);
  dff _79711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _37874_, clk);
  dff _79712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _37875_, clk);
  dff _79713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _37876_, clk);
  dff _79714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _37877_, clk);
  dff _79715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _37878_, clk);
  dff _79716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _37879_, clk);
  dff _79717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _37864_, clk);
  dff _79718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _37865_, clk);
  dff _79719_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _37866_, clk);
  dff _79720_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _37867_, clk);
  dff _79721_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _37868_, clk);
  dff _79722_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _37869_, clk);
  dff _79723_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _37870_, clk);
  dff _79724_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _37871_, clk);
  dff _79725_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _38016_, clk);
  dff _79726_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _38017_, clk);
  dff _79727_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _38018_, clk);
  dff _79728_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _38019_, clk);
  dff _79729_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _38020_, clk);
  dff _79730_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _38021_, clk);
  dff _79731_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _38022_, clk);
  dff _79732_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _38023_, clk);
  dff _79733_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _38008_, clk);
  dff _79734_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _38009_, clk);
  dff _79735_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _38010_, clk);
  dff _79736_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _38011_, clk);
  dff _79737_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _38012_, clk);
  dff _79738_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _38013_, clk);
  dff _79739_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _38014_, clk);
  dff _79740_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _38015_, clk);
  dff _79741_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _38000_, clk);
  dff _79742_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _38001_, clk);
  dff _79743_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _38002_, clk);
  dff _79744_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _38003_, clk);
  dff _79745_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _38004_, clk);
  dff _79746_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _38005_, clk);
  dff _79747_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _38006_, clk);
  dff _79748_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _38007_, clk);
  dff _79749_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _37984_, clk);
  dff _79750_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _37985_, clk);
  dff _79751_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _37986_, clk);
  dff _79752_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _37987_, clk);
  dff _79753_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _37988_, clk);
  dff _79754_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _37989_, clk);
  dff _79755_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _37990_, clk);
  dff _79756_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _37991_, clk);
  dff _79757_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _37704_, clk);
  dff _79758_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _37705_, clk);
  dff _79759_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _37706_, clk);
  dff _79760_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _37707_, clk);
  dff _79761_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _37708_, clk);
  dff _79762_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _37709_, clk);
  dff _79763_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _37710_, clk);
  dff _79764_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _37711_, clk);
  dff _79765_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _38064_, clk);
  dff _79766_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _38065_, clk);
  dff _79767_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _38066_, clk);
  dff _79768_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _38067_, clk);
  dff _79769_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _38068_, clk);
  dff _79770_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _38069_, clk);
  dff _79771_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _38070_, clk);
  dff _79772_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _38071_, clk);
  dff _79773_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _38056_, clk);
  dff _79774_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _38057_, clk);
  dff _79775_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _38058_, clk);
  dff _79776_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _38059_, clk);
  dff _79777_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _38060_, clk);
  dff _79778_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _38061_, clk);
  dff _79779_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _38062_, clk);
  dff _79780_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _38063_, clk);
  dff _79781_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _37688_, clk);
  dff _79782_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _37689_, clk);
  dff _79783_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _37690_, clk);
  dff _79784_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _37691_, clk);
  dff _79785_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _37692_, clk);
  dff _79786_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _37693_, clk);
  dff _79787_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _37694_, clk);
  dff _79788_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _37695_, clk);
  dff _79789_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _37696_, clk);
  dff _79790_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _37697_, clk);
  dff _79791_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _37698_, clk);
  dff _79792_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _37699_, clk);
  dff _79793_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _37700_, clk);
  dff _79794_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _37701_, clk);
  dff _79795_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _37702_, clk);
  dff _79796_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _37703_, clk);
  dff _79797_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _37672_, clk);
  dff _79798_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _37673_, clk);
  dff _79799_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _37674_, clk);
  dff _79800_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _37675_, clk);
  dff _79801_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _37676_, clk);
  dff _79802_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _37677_, clk);
  dff _79803_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _37678_, clk);
  dff _79804_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _37679_, clk);
  dff _79805_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _37680_, clk);
  dff _79806_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _37681_, clk);
  dff _79807_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _37682_, clk);
  dff _79808_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _37683_, clk);
  dff _79809_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _37684_, clk);
  dff _79810_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _37685_, clk);
  dff _79811_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _37686_, clk);
  dff _79812_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _37687_, clk);
  dff _79813_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _37664_, clk);
  dff _79814_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _37665_, clk);
  dff _79815_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _37666_, clk);
  dff _79816_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _37667_, clk);
  dff _79817_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _37668_, clk);
  dff _79818_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _37669_, clk);
  dff _79819_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _37670_, clk);
  dff _79820_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _37671_, clk);
  dff _79821_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _37656_, clk);
  dff _79822_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _37657_, clk);
  dff _79823_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _37658_, clk);
  dff _79824_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _37659_, clk);
  dff _79825_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _37660_, clk);
  dff _79826_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _37661_, clk);
  dff _79827_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _37662_, clk);
  dff _79828_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _37663_, clk);
  dff _79829_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _37648_, clk);
  dff _79830_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _37649_, clk);
  dff _79831_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _37650_, clk);
  dff _79832_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _37651_, clk);
  dff _79833_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _37652_, clk);
  dff _79834_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _37653_, clk);
  dff _79835_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _37654_, clk);
  dff _79836_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _37655_, clk);
  dff _79837_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _37624_, clk);
  dff _79838_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _37625_, clk);
  dff _79839_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _37626_, clk);
  dff _79840_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _37627_, clk);
  dff _79841_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _37628_, clk);
  dff _79842_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _37629_, clk);
  dff _79843_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _37630_, clk);
  dff _79844_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _37631_, clk);
  dff _79845_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _37640_, clk);
  dff _79846_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _37641_, clk);
  dff _79847_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _37642_, clk);
  dff _79848_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _37643_, clk);
  dff _79849_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _37644_, clk);
  dff _79850_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _37645_, clk);
  dff _79851_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _37646_, clk);
  dff _79852_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _37647_, clk);
  dff _79853_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _37816_, clk);
  dff _79854_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _37817_, clk);
  dff _79855_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _37818_, clk);
  dff _79856_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _37819_, clk);
  dff _79857_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _37820_, clk);
  dff _79858_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _37821_, clk);
  dff _79859_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _37822_, clk);
  dff _79860_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _37823_, clk);
  dff _79861_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _36928_, clk);
  dff _79862_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _36929_, clk);
  dff _79863_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _36930_, clk);
  dff _79864_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _36931_, clk);
  dff _79865_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _36932_, clk);
  dff _79866_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _36933_, clk);
  dff _79867_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _36934_, clk);
  dff _79868_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _36935_, clk);
  dff _79869_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _38536_, clk);
  dff _79870_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _38537_, clk);
  dff _79871_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _38538_, clk);
  dff _79872_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _38539_, clk);
  dff _79873_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _38540_, clk);
  dff _79874_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _38541_, clk);
  dff _79875_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _38542_, clk);
  dff _79876_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _38543_, clk);
  dff _79877_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _38448_, clk);
  dff _79878_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _38449_, clk);
  dff _79879_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _38450_, clk);
  dff _79880_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _38451_, clk);
  dff _79881_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _38452_, clk);
  dff _79882_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _38453_, clk);
  dff _79883_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _38454_, clk);
  dff _79884_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _38455_, clk);
  dff _79885_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _38360_, clk);
  dff _79886_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _38361_, clk);
  dff _79887_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _38362_, clk);
  dff _79888_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _38363_, clk);
  dff _79889_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _38364_, clk);
  dff _79890_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _38365_, clk);
  dff _79891_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _38366_, clk);
  dff _79892_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _38367_, clk);
  dff _79893_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _38800_, clk);
  dff _79894_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _38801_, clk);
  dff _79895_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _38802_, clk);
  dff _79896_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _38803_, clk);
  dff _79897_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _38804_, clk);
  dff _79898_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _38805_, clk);
  dff _79899_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _38806_, clk);
  dff _79900_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _38807_, clk);
  dff _79901_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _38712_, clk);
  dff _79902_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _38713_, clk);
  dff _79903_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _38714_, clk);
  dff _79904_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _38715_, clk);
  dff _79905_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _38716_, clk);
  dff _79906_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _38717_, clk);
  dff _79907_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _38718_, clk);
  dff _79908_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _38719_, clk);
  dff _79909_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _38624_, clk);
  dff _79910_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _38625_, clk);
  dff _79911_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _38626_, clk);
  dff _79912_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _38627_, clk);
  dff _79913_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _38628_, clk);
  dff _79914_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _38629_, clk);
  dff _79915_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _38630_, clk);
  dff _79916_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _38631_, clk);
  dff _79917_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _38920_, clk);
  dff _79918_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _38921_, clk);
  dff _79919_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _38922_, clk);
  dff _79920_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _38923_, clk);
  dff _79921_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _38924_, clk);
  dff _79922_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _38925_, clk);
  dff _79923_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _38926_, clk);
  dff _79924_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _38927_, clk);
  dff _79925_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _38912_, clk);
  dff _79926_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _38913_, clk);
  dff _79927_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _38914_, clk);
  dff _79928_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _38915_, clk);
  dff _79929_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _38916_, clk);
  dff _79930_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _38917_, clk);
  dff _79931_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _38918_, clk);
  dff _79932_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _38919_, clk);
  dff _79933_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _38904_, clk);
  dff _79934_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _38905_, clk);
  dff _79935_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _38906_, clk);
  dff _79936_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _38907_, clk);
  dff _79937_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _38908_, clk);
  dff _79938_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _38909_, clk);
  dff _79939_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _38910_, clk);
  dff _79940_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _38911_, clk);
  dff _79941_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _38896_, clk);
  dff _79942_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _38897_, clk);
  dff _79943_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _38898_, clk);
  dff _79944_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _38899_, clk);
  dff _79945_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _38900_, clk);
  dff _79946_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _38901_, clk);
  dff _79947_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _38902_, clk);
  dff _79948_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _38903_, clk);
  dff _79949_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _38880_, clk);
  dff _79950_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _38881_, clk);
  dff _79951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _38882_, clk);
  dff _79952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _38883_, clk);
  dff _79953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _38884_, clk);
  dff _79954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _38885_, clk);
  dff _79955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _38886_, clk);
  dff _79956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _38887_, clk);
  dff _79957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _38872_, clk);
  dff _79958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _38873_, clk);
  dff _79959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _38874_, clk);
  dff _79960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _38875_, clk);
  dff _79961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _38876_, clk);
  dff _79962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _38877_, clk);
  dff _79963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _38878_, clk);
  dff _79964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _38879_, clk);
  dff _79965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _38864_, clk);
  dff _79966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _38865_, clk);
  dff _79967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _38866_, clk);
  dff _79968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _38867_, clk);
  dff _79969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _38868_, clk);
  dff _79970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _38869_, clk);
  dff _79971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _38870_, clk);
  dff _79972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _38871_, clk);
  dff _79973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _38856_, clk);
  dff _79974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _38857_, clk);
  dff _79975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _38858_, clk);
  dff _79976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _38859_, clk);
  dff _79977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _38860_, clk);
  dff _79978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _38861_, clk);
  dff _79979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _38862_, clk);
  dff _79980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _38863_, clk);
  dff _79981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _38848_, clk);
  dff _79982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _38849_, clk);
  dff _79983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _38850_, clk);
  dff _79984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _38851_, clk);
  dff _79985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _38852_, clk);
  dff _79986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _38853_, clk);
  dff _79987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _38854_, clk);
  dff _79988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _38855_, clk);
  dff _79989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _38840_, clk);
  dff _79990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _38841_, clk);
  dff _79991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _38842_, clk);
  dff _79992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _38843_, clk);
  dff _79993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _38844_, clk);
  dff _79994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _38845_, clk);
  dff _79995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _38846_, clk);
  dff _79996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _38847_, clk);
  dff _79997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _38832_, clk);
  dff _79998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _38833_, clk);
  dff _79999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _38834_, clk);
  dff _80000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _38835_, clk);
  dff _80001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _38836_, clk);
  dff _80002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _38837_, clk);
  dff _80003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _38838_, clk);
  dff _80004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _38839_, clk);
  dff _80005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _38824_, clk);
  dff _80006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _38825_, clk);
  dff _80007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _38826_, clk);
  dff _80008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _38827_, clk);
  dff _80009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _38828_, clk);
  dff _80010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _38829_, clk);
  dff _80011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _38830_, clk);
  dff _80012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _38831_, clk);
  dff _80013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _38816_, clk);
  dff _80014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _38817_, clk);
  dff _80015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _38818_, clk);
  dff _80016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _38819_, clk);
  dff _80017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _38820_, clk);
  dff _80018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _38821_, clk);
  dff _80019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _38822_, clk);
  dff _80020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _38823_, clk);
  dff _80021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _38808_, clk);
  dff _80022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _38809_, clk);
  dff _80023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _38810_, clk);
  dff _80024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _38811_, clk);
  dff _80025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _38812_, clk);
  dff _80026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _38813_, clk);
  dff _80027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _38814_, clk);
  dff _80028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _38815_, clk);
  dff _80029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _38792_, clk);
  dff _80030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _38793_, clk);
  dff _80031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _38794_, clk);
  dff _80032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _38795_, clk);
  dff _80033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _38796_, clk);
  dff _80034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _38797_, clk);
  dff _80035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _38798_, clk);
  dff _80036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _38799_, clk);
  dff _80037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _38784_, clk);
  dff _80038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _38785_, clk);
  dff _80039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _38786_, clk);
  dff _80040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _38787_, clk);
  dff _80041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _38788_, clk);
  dff _80042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _38789_, clk);
  dff _80043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _38790_, clk);
  dff _80044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _38791_, clk);
  dff _80045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _38776_, clk);
  dff _80046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _38777_, clk);
  dff _80047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _38778_, clk);
  dff _80048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _38779_, clk);
  dff _80049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _38780_, clk);
  dff _80050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _38781_, clk);
  dff _80051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _38782_, clk);
  dff _80052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _38783_, clk);
  dff _80053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _38768_, clk);
  dff _80054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _38769_, clk);
  dff _80055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _38770_, clk);
  dff _80056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _38771_, clk);
  dff _80057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _38772_, clk);
  dff _80058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _38773_, clk);
  dff _80059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _38774_, clk);
  dff _80060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _38775_, clk);
  dff _80061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _38760_, clk);
  dff _80062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _38761_, clk);
  dff _80063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _38762_, clk);
  dff _80064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _38763_, clk);
  dff _80065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _38764_, clk);
  dff _80066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _38765_, clk);
  dff _80067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _38766_, clk);
  dff _80068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _38767_, clk);
  dff _80069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _38752_, clk);
  dff _80070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _38753_, clk);
  dff _80071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _38754_, clk);
  dff _80072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _38755_, clk);
  dff _80073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _38756_, clk);
  dff _80074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _38757_, clk);
  dff _80075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _38758_, clk);
  dff _80076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _38759_, clk);
  dff _80077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _38744_, clk);
  dff _80078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _38745_, clk);
  dff _80079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _38746_, clk);
  dff _80080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _38747_, clk);
  dff _80081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _38748_, clk);
  dff _80082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _38749_, clk);
  dff _80083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _38750_, clk);
  dff _80084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _38751_, clk);
  dff _80085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _38736_, clk);
  dff _80086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _38737_, clk);
  dff _80087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _38738_, clk);
  dff _80088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _38739_, clk);
  dff _80089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _38740_, clk);
  dff _80090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _38741_, clk);
  dff _80091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _38742_, clk);
  dff _80092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _38743_, clk);
  dff _80093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _38728_, clk);
  dff _80094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _38729_, clk);
  dff _80095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _38730_, clk);
  dff _80096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _38731_, clk);
  dff _80097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _38732_, clk);
  dff _80098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _38733_, clk);
  dff _80099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _38734_, clk);
  dff _80100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _38735_, clk);
  dff _80101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _38720_, clk);
  dff _80102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _38721_, clk);
  dff _80103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _38722_, clk);
  dff _80104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _38723_, clk);
  dff _80105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _38724_, clk);
  dff _80106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _38725_, clk);
  dff _80107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _38726_, clk);
  dff _80108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _38727_, clk);
  dff _80109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _38704_, clk);
  dff _80110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _38705_, clk);
  dff _80111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _38706_, clk);
  dff _80112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _38707_, clk);
  dff _80113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _38708_, clk);
  dff _80114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _38709_, clk);
  dff _80115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _38710_, clk);
  dff _80116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _38711_, clk);
  dff _80117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _38696_, clk);
  dff _80118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _38697_, clk);
  dff _80119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _38698_, clk);
  dff _80120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _38699_, clk);
  dff _80121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _38700_, clk);
  dff _80122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _38701_, clk);
  dff _80123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _38702_, clk);
  dff _80124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _38703_, clk);
  dff _80125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _38688_, clk);
  dff _80126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _38689_, clk);
  dff _80127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _38690_, clk);
  dff _80128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _38691_, clk);
  dff _80129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _38692_, clk);
  dff _80130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _38693_, clk);
  dff _80131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _38694_, clk);
  dff _80132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _38695_, clk);
  dff _80133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _38680_, clk);
  dff _80134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _38681_, clk);
  dff _80135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _38682_, clk);
  dff _80136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _38683_, clk);
  dff _80137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _38684_, clk);
  dff _80138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _38685_, clk);
  dff _80139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _38686_, clk);
  dff _80140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _38687_, clk);
  dff _80141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _38672_, clk);
  dff _80142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _38673_, clk);
  dff _80143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _38674_, clk);
  dff _80144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _38675_, clk);
  dff _80145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _38676_, clk);
  dff _80146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _38677_, clk);
  dff _80147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _38678_, clk);
  dff _80148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _38679_, clk);
  dff _80149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _38664_, clk);
  dff _80150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _38665_, clk);
  dff _80151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _38666_, clk);
  dff _80152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _38667_, clk);
  dff _80153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _38668_, clk);
  dff _80154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _38669_, clk);
  dff _80155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _38670_, clk);
  dff _80156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _38671_, clk);
  dff _80157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _38656_, clk);
  dff _80158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _38657_, clk);
  dff _80159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _38658_, clk);
  dff _80160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _38659_, clk);
  dff _80161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _38660_, clk);
  dff _80162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _38661_, clk);
  dff _80163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _38662_, clk);
  dff _80164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _38663_, clk);
  dff _80165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _38648_, clk);
  dff _80166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _38649_, clk);
  dff _80167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _38650_, clk);
  dff _80168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _38651_, clk);
  dff _80169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _38652_, clk);
  dff _80170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _38653_, clk);
  dff _80171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _38654_, clk);
  dff _80172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _38655_, clk);
  dff _80173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _38640_, clk);
  dff _80174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _38641_, clk);
  dff _80175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _38642_, clk);
  dff _80176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _38643_, clk);
  dff _80177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _38644_, clk);
  dff _80178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _38645_, clk);
  dff _80179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _38646_, clk);
  dff _80180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _38647_, clk);
  dff _80181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _38632_, clk);
  dff _80182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _38633_, clk);
  dff _80183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _38634_, clk);
  dff _80184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _38635_, clk);
  dff _80185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _38636_, clk);
  dff _80186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _38637_, clk);
  dff _80187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _38638_, clk);
  dff _80188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _38639_, clk);
  dff _80189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _38616_, clk);
  dff _80190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _38617_, clk);
  dff _80191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _38618_, clk);
  dff _80192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _38619_, clk);
  dff _80193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _38620_, clk);
  dff _80194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _38621_, clk);
  dff _80195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _38622_, clk);
  dff _80196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _38623_, clk);
  dff _80197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _38608_, clk);
  dff _80198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _38609_, clk);
  dff _80199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _38610_, clk);
  dff _80200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _38611_, clk);
  dff _80201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _38612_, clk);
  dff _80202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _38613_, clk);
  dff _80203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _38614_, clk);
  dff _80204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _38615_, clk);
  dff _80205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _38600_, clk);
  dff _80206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _38601_, clk);
  dff _80207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _38602_, clk);
  dff _80208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _38603_, clk);
  dff _80209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _38604_, clk);
  dff _80210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _38605_, clk);
  dff _80211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _38606_, clk);
  dff _80212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _38607_, clk);
  dff _80213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _38592_, clk);
  dff _80214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _38593_, clk);
  dff _80215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _38594_, clk);
  dff _80216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _38595_, clk);
  dff _80217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _38596_, clk);
  dff _80218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _38597_, clk);
  dff _80219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _38598_, clk);
  dff _80220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _38599_, clk);
  dff _80221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _38584_, clk);
  dff _80222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _38585_, clk);
  dff _80223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _38586_, clk);
  dff _80224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _38587_, clk);
  dff _80225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _38588_, clk);
  dff _80226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _38589_, clk);
  dff _80227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _38590_, clk);
  dff _80228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _38591_, clk);
  dff _80229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _38576_, clk);
  dff _80230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _38577_, clk);
  dff _80231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _38578_, clk);
  dff _80232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _38579_, clk);
  dff _80233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _38580_, clk);
  dff _80234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _38581_, clk);
  dff _80235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _38582_, clk);
  dff _80236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _38583_, clk);
  dff _80237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _38568_, clk);
  dff _80238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _38569_, clk);
  dff _80239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _38570_, clk);
  dff _80240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _38571_, clk);
  dff _80241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _38572_, clk);
  dff _80242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _38573_, clk);
  dff _80243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _38574_, clk);
  dff _80244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _38575_, clk);
  dff _80245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _38560_, clk);
  dff _80246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _38561_, clk);
  dff _80247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _38562_, clk);
  dff _80248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _38563_, clk);
  dff _80249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _38564_, clk);
  dff _80250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _38565_, clk);
  dff _80251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _38566_, clk);
  dff _80252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _38567_, clk);
  dff _80253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _38552_, clk);
  dff _80254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _38553_, clk);
  dff _80255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _38554_, clk);
  dff _80256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _38555_, clk);
  dff _80257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _38556_, clk);
  dff _80258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _38557_, clk);
  dff _80259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _38558_, clk);
  dff _80260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _38559_, clk);
  dff _80261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _38544_, clk);
  dff _80262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _38545_, clk);
  dff _80263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _38546_, clk);
  dff _80264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _38547_, clk);
  dff _80265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _38548_, clk);
  dff _80266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _38549_, clk);
  dff _80267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _38550_, clk);
  dff _80268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _38551_, clk);
  dff _80269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _38528_, clk);
  dff _80270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _38529_, clk);
  dff _80271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _38530_, clk);
  dff _80272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _38531_, clk);
  dff _80273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _38532_, clk);
  dff _80274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _38533_, clk);
  dff _80275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _38534_, clk);
  dff _80276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _38535_, clk);
  dff _80277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _38520_, clk);
  dff _80278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _38521_, clk);
  dff _80279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _38522_, clk);
  dff _80280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _38523_, clk);
  dff _80281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _38524_, clk);
  dff _80282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _38525_, clk);
  dff _80283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _38526_, clk);
  dff _80284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _38527_, clk);
  dff _80285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _38512_, clk);
  dff _80286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _38513_, clk);
  dff _80287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _38514_, clk);
  dff _80288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _38515_, clk);
  dff _80289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _38516_, clk);
  dff _80290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _38517_, clk);
  dff _80291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _38518_, clk);
  dff _80292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _38519_, clk);
  dff _80293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _38504_, clk);
  dff _80294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _38505_, clk);
  dff _80295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _38506_, clk);
  dff _80296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _38507_, clk);
  dff _80297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _38508_, clk);
  dff _80298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _38509_, clk);
  dff _80299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _38510_, clk);
  dff _80300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _38511_, clk);
  dff _80301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _38496_, clk);
  dff _80302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _38497_, clk);
  dff _80303_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _38498_, clk);
  dff _80304_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _38499_, clk);
  dff _80305_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _38500_, clk);
  dff _80306_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _38501_, clk);
  dff _80307_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _38502_, clk);
  dff _80308_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _38503_, clk);
  dff _80309_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _38488_, clk);
  dff _80310_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _38489_, clk);
  dff _80311_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _38490_, clk);
  dff _80312_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _38491_, clk);
  dff _80313_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _38492_, clk);
  dff _80314_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _38493_, clk);
  dff _80315_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _38494_, clk);
  dff _80316_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _38495_, clk);
  dff _80317_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _38480_, clk);
  dff _80318_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _38481_, clk);
  dff _80319_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _38482_, clk);
  dff _80320_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _38483_, clk);
  dff _80321_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _38484_, clk);
  dff _80322_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _38485_, clk);
  dff _80323_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _38486_, clk);
  dff _80324_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _38487_, clk);
  dff _80325_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _38472_, clk);
  dff _80326_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _38473_, clk);
  dff _80327_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _38474_, clk);
  dff _80328_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _38475_, clk);
  dff _80329_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _38476_, clk);
  dff _80330_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _38477_, clk);
  dff _80331_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _38478_, clk);
  dff _80332_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _38479_, clk);
  dff _80333_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _38464_, clk);
  dff _80334_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _38465_, clk);
  dff _80335_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _38466_, clk);
  dff _80336_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _38467_, clk);
  dff _80337_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _38468_, clk);
  dff _80338_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _38469_, clk);
  dff _80339_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _38470_, clk);
  dff _80340_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _38471_, clk);
  dff _80341_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _38456_, clk);
  dff _80342_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _38457_, clk);
  dff _80343_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _38458_, clk);
  dff _80344_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _38459_, clk);
  dff _80345_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _38460_, clk);
  dff _80346_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _38461_, clk);
  dff _80347_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _38462_, clk);
  dff _80348_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _38463_, clk);
  dff _80349_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _38440_, clk);
  dff _80350_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _38441_, clk);
  dff _80351_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _38442_, clk);
  dff _80352_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _38443_, clk);
  dff _80353_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _38444_, clk);
  dff _80354_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _38445_, clk);
  dff _80355_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _38446_, clk);
  dff _80356_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _38447_, clk);
  dff _80357_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _38432_, clk);
  dff _80358_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _38433_, clk);
  dff _80359_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _38434_, clk);
  dff _80360_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _38435_, clk);
  dff _80361_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _38436_, clk);
  dff _80362_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _38437_, clk);
  dff _80363_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _38438_, clk);
  dff _80364_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _38439_, clk);
  dff _80365_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _38424_, clk);
  dff _80366_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _38425_, clk);
  dff _80367_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _38426_, clk);
  dff _80368_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _38427_, clk);
  dff _80369_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _38428_, clk);
  dff _80370_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _38429_, clk);
  dff _80371_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _38430_, clk);
  dff _80372_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _38431_, clk);
  dff _80373_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _38416_, clk);
  dff _80374_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _38417_, clk);
  dff _80375_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _38418_, clk);
  dff _80376_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _38419_, clk);
  dff _80377_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _38420_, clk);
  dff _80378_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _38421_, clk);
  dff _80379_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _38422_, clk);
  dff _80380_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _38423_, clk);
  dff _80381_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _38408_, clk);
  dff _80382_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _38409_, clk);
  dff _80383_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _38410_, clk);
  dff _80384_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _38411_, clk);
  dff _80385_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _38412_, clk);
  dff _80386_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _38413_, clk);
  dff _80387_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _38414_, clk);
  dff _80388_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _38415_, clk);
  dff _80389_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _38400_, clk);
  dff _80390_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _38401_, clk);
  dff _80391_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _38402_, clk);
  dff _80392_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _38403_, clk);
  dff _80393_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _38404_, clk);
  dff _80394_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _38405_, clk);
  dff _80395_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _38406_, clk);
  dff _80396_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _38407_, clk);
  dff _80397_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _38392_, clk);
  dff _80398_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _38393_, clk);
  dff _80399_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _38394_, clk);
  dff _80400_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _38395_, clk);
  dff _80401_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _38396_, clk);
  dff _80402_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _38397_, clk);
  dff _80403_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _38398_, clk);
  dff _80404_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _38399_, clk);
  dff _80405_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _38384_, clk);
  dff _80406_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _38385_, clk);
  dff _80407_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _38386_, clk);
  dff _80408_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _38387_, clk);
  dff _80409_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _38388_, clk);
  dff _80410_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _38389_, clk);
  dff _80411_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _38390_, clk);
  dff _80412_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _38391_, clk);
  dff _80413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _38376_, clk);
  dff _80414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _38377_, clk);
  dff _80415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _38378_, clk);
  dff _80416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _38379_, clk);
  dff _80417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _38380_, clk);
  dff _80418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _38381_, clk);
  dff _80419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _38382_, clk);
  dff _80420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _38383_, clk);
  dff _80421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _38368_, clk);
  dff _80422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _38369_, clk);
  dff _80423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _38370_, clk);
  dff _80424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _38371_, clk);
  dff _80425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _38372_, clk);
  dff _80426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _38373_, clk);
  dff _80427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _38374_, clk);
  dff _80428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _38375_, clk);
  dff _80429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _38352_, clk);
  dff _80430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _38353_, clk);
  dff _80431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _38354_, clk);
  dff _80432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _38355_, clk);
  dff _80433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _38356_, clk);
  dff _80434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _38357_, clk);
  dff _80435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _38358_, clk);
  dff _80436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _38359_, clk);
  dff _80437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _38344_, clk);
  dff _80438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _38345_, clk);
  dff _80439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _38346_, clk);
  dff _80440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _38347_, clk);
  dff _80441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _38348_, clk);
  dff _80442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _38349_, clk);
  dff _80443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _38350_, clk);
  dff _80444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _38351_, clk);
  dff _80445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _38336_, clk);
  dff _80446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _38337_, clk);
  dff _80447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _38338_, clk);
  dff _80448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _38339_, clk);
  dff _80449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _38340_, clk);
  dff _80450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _38341_, clk);
  dff _80451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _38342_, clk);
  dff _80452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _38343_, clk);
  dff _80453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _38328_, clk);
  dff _80454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _38329_, clk);
  dff _80455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _38330_, clk);
  dff _80456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _38331_, clk);
  dff _80457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _38332_, clk);
  dff _80458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _38333_, clk);
  dff _80459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _38334_, clk);
  dff _80460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _38335_, clk);
  dff _80461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _38320_, clk);
  dff _80462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _38321_, clk);
  dff _80463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _38322_, clk);
  dff _80464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _38323_, clk);
  dff _80465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _38324_, clk);
  dff _80466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _38325_, clk);
  dff _80467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _38326_, clk);
  dff _80468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _38327_, clk);
  dff _80469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _38256_, clk);
  dff _80470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _38257_, clk);
  dff _80471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _38258_, clk);
  dff _80472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _38259_, clk);
  dff _80473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _38260_, clk);
  dff _80474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _38261_, clk);
  dff _80475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _38262_, clk);
  dff _80476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _38263_, clk);
  dff _80477_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _38168_, clk);
  dff _80478_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _38169_, clk);
  dff _80479_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _38170_, clk);
  dff _80480_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _38171_, clk);
  dff _80481_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _38172_, clk);
  dff _80482_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _38173_, clk);
  dff _80483_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _38174_, clk);
  dff _80484_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _38175_, clk);
  dff _80485_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _38080_, clk);
  dff _80486_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _38081_, clk);
  dff _80487_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _38082_, clk);
  dff _80488_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _38083_, clk);
  dff _80489_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _38084_, clk);
  dff _80490_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _38085_, clk);
  dff _80491_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _38086_, clk);
  dff _80492_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _38087_, clk);
  dff _80493_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _37992_, clk);
  dff _80494_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _37993_, clk);
  dff _80495_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _37994_, clk);
  dff _80496_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _37995_, clk);
  dff _80497_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _37996_, clk);
  dff _80498_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _37997_, clk);
  dff _80499_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _37998_, clk);
  dff _80500_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _37999_, clk);
  dff _80501_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _37904_, clk);
  dff _80502_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _37905_, clk);
  dff _80503_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _37906_, clk);
  dff _80504_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _37907_, clk);
  dff _80505_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _37908_, clk);
  dff _80506_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _37909_, clk);
  dff _80507_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _37910_, clk);
  dff _80508_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _37911_, clk);
  dff _80509_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _37808_, clk);
  dff _80510_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _37809_, clk);
  dff _80511_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _37810_, clk);
  dff _80512_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _37811_, clk);
  dff _80513_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _37812_, clk);
  dff _80514_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _37813_, clk);
  dff _80515_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _37814_, clk);
  dff _80516_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _37815_, clk);
  dff _80517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _37720_, clk);
  dff _80518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _37721_, clk);
  dff _80519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _37722_, clk);
  dff _80520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _37723_, clk);
  dff _80521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _37724_, clk);
  dff _80522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _37725_, clk);
  dff _80523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _37726_, clk);
  dff _80524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _37727_, clk);
  dff _80525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _37632_, clk);
  dff _80526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _37633_, clk);
  dff _80527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _37634_, clk);
  dff _80528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _37635_, clk);
  dff _80529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _37636_, clk);
  dff _80530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _37637_, clk);
  dff _80531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _37638_, clk);
  dff _80532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _37639_, clk);
  dff _80533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _37544_, clk);
  dff _80534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _37545_, clk);
  dff _80535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _37546_, clk);
  dff _80536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _37547_, clk);
  dff _80537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _37548_, clk);
  dff _80538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _37549_, clk);
  dff _80539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _37550_, clk);
  dff _80540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _37551_, clk);
  dff _80541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _37456_, clk);
  dff _80542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _37457_, clk);
  dff _80543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _37458_, clk);
  dff _80544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _37459_, clk);
  dff _80545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _37460_, clk);
  dff _80546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _37461_, clk);
  dff _80547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _37462_, clk);
  dff _80548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _37463_, clk);
  dff _80549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _37368_, clk);
  dff _80550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _37369_, clk);
  dff _80551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _37370_, clk);
  dff _80552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _37371_, clk);
  dff _80553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _37372_, clk);
  dff _80554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _37373_, clk);
  dff _80555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _37374_, clk);
  dff _80556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _37375_, clk);
  dff _80557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _37280_, clk);
  dff _80558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _37281_, clk);
  dff _80559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _37282_, clk);
  dff _80560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _37283_, clk);
  dff _80561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _37284_, clk);
  dff _80562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _37285_, clk);
  dff _80563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _37286_, clk);
  dff _80564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _37287_, clk);
  dff _80565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _37192_, clk);
  dff _80566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _37193_, clk);
  dff _80567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _37194_, clk);
  dff _80568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _37195_, clk);
  dff _80569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _37196_, clk);
  dff _80570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _37197_, clk);
  dff _80571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _37198_, clk);
  dff _80572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _37199_, clk);
  dff _80573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _37104_, clk);
  dff _80574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _37105_, clk);
  dff _80575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _37106_, clk);
  dff _80576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _37107_, clk);
  dff _80577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _37108_, clk);
  dff _80578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _37109_, clk);
  dff _80579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _37110_, clk);
  dff _80580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _37111_, clk);
  dff _80581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _37016_, clk);
  dff _80582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _37017_, clk);
  dff _80583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _37018_, clk);
  dff _80584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _37019_, clk);
  dff _80585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _37020_, clk);
  dff _80586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _37021_, clk);
  dff _80587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _37022_, clk);
  dff _80588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _37023_, clk);
  dff _80589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _38976_, clk);
  dff _80590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _38977_, clk);
  dff _80591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _38978_, clk);
  dff _80592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _38979_, clk);
  dff _80593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _38980_, clk);
  dff _80594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _38981_, clk);
  dff _80595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _38982_, clk);
  dff _80596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _38983_, clk);
  dff _80597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _38888_, clk);
  dff _80598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _38889_, clk);
  dff _80599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _38890_, clk);
  dff _80600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _38891_, clk);
  dff _80601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _38892_, clk);
  dff _80602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _38893_, clk);
  dff _80603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _38894_, clk);
  dff _80604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _38895_, clk);
  dff _80605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _38048_, clk);
  dff _80606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _38049_, clk);
  dff _80607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _38050_, clk);
  dff _80608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _38051_, clk);
  dff _80609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _38052_, clk);
  dff _80610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _38053_, clk);
  dff _80611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _38054_, clk);
  dff _80612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _38055_, clk);
  dff _80613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _37976_, clk);
  dff _80614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _37977_, clk);
  dff _80615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _37978_, clk);
  dff _80616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _37979_, clk);
  dff _80617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _37980_, clk);
  dff _80618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _37981_, clk);
  dff _80619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _37982_, clk);
  dff _80620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _37983_, clk);
  dff _80621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _37856_, clk);
  dff _80622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _37857_, clk);
  dff _80623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _37858_, clk);
  dff _80624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _37859_, clk);
  dff _80625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _37860_, clk);
  dff _80626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _37861_, clk);
  dff _80627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _37862_, clk);
  dff _80628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _37863_, clk);
  dff _80629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _37848_, clk);
  dff _80630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _37849_, clk);
  dff _80631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _37850_, clk);
  dff _80632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _37851_, clk);
  dff _80633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _37852_, clk);
  dff _80634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _37853_, clk);
  dff _80635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _37854_, clk);
  dff _80636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _37855_, clk);
  dff _80637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _37840_, clk);
  dff _80638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _37841_, clk);
  dff _80639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _37842_, clk);
  dff _80640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _37843_, clk);
  dff _80641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _37844_, clk);
  dff _80642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _37845_, clk);
  dff _80643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _37846_, clk);
  dff _80644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _37847_, clk);
  dff _80645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _37832_, clk);
  dff _80646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _37833_, clk);
  dff _80647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _37834_, clk);
  dff _80648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _37835_, clk);
  dff _80649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _37836_, clk);
  dff _80650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _37837_, clk);
  dff _80651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _37838_, clk);
  dff _80652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _37839_, clk);
  dff _80653_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _37824_, clk);
  dff _80654_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _37825_, clk);
  dff _80655_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _37826_, clk);
  dff _80656_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _37827_, clk);
  dff _80657_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _37828_, clk);
  dff _80658_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _37829_, clk);
  dff _80659_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _37830_, clk);
  dff _80660_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _37831_, clk);
  dff _80661_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _37800_, clk);
  dff _80662_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _37801_, clk);
  dff _80663_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _37802_, clk);
  dff _80664_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _37803_, clk);
  dff _80665_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _37804_, clk);
  dff _80666_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _37805_, clk);
  dff _80667_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _37806_, clk);
  dff _80668_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _37807_, clk);
  dff _80669_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _37792_, clk);
  dff _80670_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _37793_, clk);
  dff _80671_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _37794_, clk);
  dff _80672_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _37795_, clk);
  dff _80673_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _37796_, clk);
  dff _80674_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _37797_, clk);
  dff _80675_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _37798_, clk);
  dff _80676_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _37799_, clk);
  dff _80677_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _37784_, clk);
  dff _80678_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _37785_, clk);
  dff _80679_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _37786_, clk);
  dff _80680_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _37787_, clk);
  dff _80681_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _37788_, clk);
  dff _80682_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _37789_, clk);
  dff _80683_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _37790_, clk);
  dff _80684_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _37791_, clk);
  dff _80685_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _37776_, clk);
  dff _80686_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _37777_, clk);
  dff _80687_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _37778_, clk);
  dff _80688_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _37779_, clk);
  dff _80689_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _37780_, clk);
  dff _80690_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _37781_, clk);
  dff _80691_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _37782_, clk);
  dff _80692_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _37783_, clk);
  dff _80693_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _37768_, clk);
  dff _80694_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _37769_, clk);
  dff _80695_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _37770_, clk);
  dff _80696_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _37771_, clk);
  dff _80697_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _37772_, clk);
  dff _80698_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _37773_, clk);
  dff _80699_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _37774_, clk);
  dff _80700_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _37775_, clk);
  dff _80701_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _37760_, clk);
  dff _80702_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _37761_, clk);
  dff _80703_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _37762_, clk);
  dff _80704_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _37763_, clk);
  dff _80705_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _37764_, clk);
  dff _80706_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _37765_, clk);
  dff _80707_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _37766_, clk);
  dff _80708_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _37767_, clk);
  dff _80709_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _37752_, clk);
  dff _80710_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _37753_, clk);
  dff _80711_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _37754_, clk);
  dff _80712_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _37755_, clk);
  dff _80713_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _37756_, clk);
  dff _80714_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _37757_, clk);
  dff _80715_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _37758_, clk);
  dff _80716_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _37759_, clk);
  dff _80717_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _37744_, clk);
  dff _80718_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _37745_, clk);
  dff _80719_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _37746_, clk);
  dff _80720_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _37747_, clk);
  dff _80721_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _37748_, clk);
  dff _80722_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _37749_, clk);
  dff _80723_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _37750_, clk);
  dff _80724_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _37751_, clk);
  dff _80725_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _37736_, clk);
  dff _80726_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _37737_, clk);
  dff _80727_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _37738_, clk);
  dff _80728_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _37739_, clk);
  dff _80729_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _37740_, clk);
  dff _80730_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _37741_, clk);
  dff _80731_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _37742_, clk);
  dff _80732_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _37743_, clk);
  dff _80733_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _37728_, clk);
  dff _80734_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _37729_, clk);
  dff _80735_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _37730_, clk);
  dff _80736_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _37731_, clk);
  dff _80737_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _37732_, clk);
  dff _80738_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _37733_, clk);
  dff _80739_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _37734_, clk);
  dff _80740_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _37735_, clk);
  dff _80741_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _37712_, clk);
  dff _80742_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _37713_, clk);
  dff _80743_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _37714_, clk);
  dff _80744_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _37715_, clk);
  dff _80745_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _37716_, clk);
  dff _80746_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _37717_, clk);
  dff _80747_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _37718_, clk);
  dff _80748_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _37719_, clk);
  dff _80749_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _37392_, clk);
  dff _80750_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _37393_, clk);
  dff _80751_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _37394_, clk);
  dff _80752_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _37395_, clk);
  dff _80753_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _37396_, clk);
  dff _80754_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _37397_, clk);
  dff _80755_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _37398_, clk);
  dff _80756_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _37399_, clk);
  dff _80757_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _37512_, clk);
  dff _80758_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _37513_, clk);
  dff _80759_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _37514_, clk);
  dff _80760_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _37515_, clk);
  dff _80761_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _37516_, clk);
  dff _80762_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _37517_, clk);
  dff _80763_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _37518_, clk);
  dff _80764_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _37519_, clk);
  dff _80765_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _37384_, clk);
  dff _80766_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _37385_, clk);
  dff _80767_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _37386_, clk);
  dff _80768_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _37387_, clk);
  dff _80769_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _37388_, clk);
  dff _80770_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _37389_, clk);
  dff _80771_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _37390_, clk);
  dff _80772_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _37391_, clk);
  dff _80773_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _37504_, clk);
  dff _80774_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _37505_, clk);
  dff _80775_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _37506_, clk);
  dff _80776_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _37507_, clk);
  dff _80777_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _37508_, clk);
  dff _80778_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _37509_, clk);
  dff _80779_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _37510_, clk);
  dff _80780_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _37511_, clk);
  dff _80781_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _37376_, clk);
  dff _80782_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _37377_, clk);
  dff _80783_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _37378_, clk);
  dff _80784_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _37379_, clk);
  dff _80785_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _37380_, clk);
  dff _80786_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _37381_, clk);
  dff _80787_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _37382_, clk);
  dff _80788_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _37383_, clk);
  dff _80789_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _37496_, clk);
  dff _80790_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _37497_, clk);
  dff _80791_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _37498_, clk);
  dff _80792_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _37499_, clk);
  dff _80793_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _37500_, clk);
  dff _80794_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _37501_, clk);
  dff _80795_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _37502_, clk);
  dff _80796_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _37503_, clk);
  dff _80797_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _37360_, clk);
  dff _80798_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _37361_, clk);
  dff _80799_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _37362_, clk);
  dff _80800_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _37363_, clk);
  dff _80801_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _37364_, clk);
  dff _80802_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _37365_, clk);
  dff _80803_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _37366_, clk);
  dff _80804_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _37367_, clk);
  dff _80805_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _37488_, clk);
  dff _80806_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _37489_, clk);
  dff _80807_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _37490_, clk);
  dff _80808_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _37491_, clk);
  dff _80809_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _37492_, clk);
  dff _80810_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _37493_, clk);
  dff _80811_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _37494_, clk);
  dff _80812_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _37495_, clk);
  dff _80813_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _37352_, clk);
  dff _80814_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _37353_, clk);
  dff _80815_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _37354_, clk);
  dff _80816_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _37355_, clk);
  dff _80817_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _37356_, clk);
  dff _80818_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _37357_, clk);
  dff _80819_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _37358_, clk);
  dff _80820_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _37359_, clk);
  dff _80821_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _37344_, clk);
  dff _80822_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _37345_, clk);
  dff _80823_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _37346_, clk);
  dff _80824_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _37347_, clk);
  dff _80825_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _37348_, clk);
  dff _80826_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _37349_, clk);
  dff _80827_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _37350_, clk);
  dff _80828_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _37351_, clk);
  dff _80829_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _37336_, clk);
  dff _80830_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _37337_, clk);
  dff _80831_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _37338_, clk);
  dff _80832_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _37339_, clk);
  dff _80833_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _37340_, clk);
  dff _80834_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _37341_, clk);
  dff _80835_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _37342_, clk);
  dff _80836_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _37343_, clk);
  dff _80837_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _37328_, clk);
  dff _80838_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _37329_, clk);
  dff _80839_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _37330_, clk);
  dff _80840_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _37331_, clk);
  dff _80841_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _37332_, clk);
  dff _80842_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _37333_, clk);
  dff _80843_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _37334_, clk);
  dff _80844_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _37335_, clk);
  dff _80845_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _37320_, clk);
  dff _80846_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _37321_, clk);
  dff _80847_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _37322_, clk);
  dff _80848_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _37323_, clk);
  dff _80849_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _37324_, clk);
  dff _80850_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _37325_, clk);
  dff _80851_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _37326_, clk);
  dff _80852_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _37327_, clk);
  dff _80853_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _37312_, clk);
  dff _80854_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _37313_, clk);
  dff _80855_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _37314_, clk);
  dff _80856_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _37315_, clk);
  dff _80857_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _37316_, clk);
  dff _80858_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _37317_, clk);
  dff _80859_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _37318_, clk);
  dff _80860_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _37319_, clk);
  dff _80861_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _37304_, clk);
  dff _80862_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _37305_, clk);
  dff _80863_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _37306_, clk);
  dff _80864_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _37307_, clk);
  dff _80865_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _37308_, clk);
  dff _80866_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _37309_, clk);
  dff _80867_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _37310_, clk);
  dff _80868_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _37311_, clk);
  dff _80869_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _37296_, clk);
  dff _80870_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _37297_, clk);
  dff _80871_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _37298_, clk);
  dff _80872_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _37299_, clk);
  dff _80873_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _37300_, clk);
  dff _80874_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _37301_, clk);
  dff _80875_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _37302_, clk);
  dff _80876_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _37303_, clk);
  dff _80877_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _37288_, clk);
  dff _80878_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _37289_, clk);
  dff _80879_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _37290_, clk);
  dff _80880_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _37291_, clk);
  dff _80881_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _37292_, clk);
  dff _80882_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _37293_, clk);
  dff _80883_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _37294_, clk);
  dff _80884_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _37295_, clk);
  dff _80885_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _37248_, clk);
  dff _80886_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _37249_, clk);
  dff _80887_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _37250_, clk);
  dff _80888_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _37251_, clk);
  dff _80889_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _37252_, clk);
  dff _80890_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _37253_, clk);
  dff _80891_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _37254_, clk);
  dff _80892_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _37255_, clk);
  dff _80893_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _36992_, clk);
  dff _80894_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _36993_, clk);
  dff _80895_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _36994_, clk);
  dff _80896_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _36995_, clk);
  dff _80897_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _36996_, clk);
  dff _80898_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _36997_, clk);
  dff _80899_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _36998_, clk);
  dff _80900_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _36999_, clk);
  dff _80901_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _36984_, clk);
  dff _80902_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _36985_, clk);
  dff _80903_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _36986_, clk);
  dff _80904_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _36987_, clk);
  dff _80905_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _36988_, clk);
  dff _80906_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _36989_, clk);
  dff _80907_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _36990_, clk);
  dff _80908_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _36991_, clk);
  dff _80909_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _36976_, clk);
  dff _80910_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _36977_, clk);
  dff _80911_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _36978_, clk);
  dff _80912_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _36979_, clk);
  dff _80913_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _36980_, clk);
  dff _80914_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _36981_, clk);
  dff _80915_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _36982_, clk);
  dff _80916_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _36983_, clk);
  dff _80917_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _36968_, clk);
  dff _80918_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _36969_, clk);
  dff _80919_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _36970_, clk);
  dff _80920_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _36971_, clk);
  dff _80921_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _36972_, clk);
  dff _80922_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _36973_, clk);
  dff _80923_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _36974_, clk);
  dff _80924_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _36975_, clk);
  dff _80925_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _36960_, clk);
  dff _80926_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _36961_, clk);
  dff _80927_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _36962_, clk);
  dff _80928_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _36963_, clk);
  dff _80929_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _36964_, clk);
  dff _80930_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _36965_, clk);
  dff _80931_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _36966_, clk);
  dff _80932_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _36967_, clk);
  dff _80933_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _37176_, clk);
  dff _80934_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _37177_, clk);
  dff _80935_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _37178_, clk);
  dff _80936_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _37179_, clk);
  dff _80937_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _37180_, clk);
  dff _80938_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _37181_, clk);
  dff _80939_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _37182_, clk);
  dff _80940_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _37183_, clk);
  dff _80941_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _36952_, clk);
  dff _80942_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _36953_, clk);
  dff _80943_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _36954_, clk);
  dff _80944_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _36955_, clk);
  dff _80945_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _36956_, clk);
  dff _80946_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _36957_, clk);
  dff _80947_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _36958_, clk);
  dff _80948_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _36959_, clk);
  dff _80949_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _36944_, clk);
  dff _80950_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _36945_, clk);
  dff _80951_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _36946_, clk);
  dff _80952_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _36947_, clk);
  dff _80953_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _36948_, clk);
  dff _80954_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _36949_, clk);
  dff _80955_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _36950_, clk);
  dff _80956_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _36951_, clk);
  dff _80957_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _36936_, clk);
  dff _80958_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _36937_, clk);
  dff _80959_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _36938_, clk);
  dff _80960_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _36939_, clk);
  dff _80961_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _36940_, clk);
  dff _80962_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _36941_, clk);
  dff _80963_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _36942_, clk);
  dff _80964_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _36943_, clk);
  dff _80965_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _38968_, clk);
  dff _80966_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _38969_, clk);
  dff _80967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _38970_, clk);
  dff _80968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _38971_, clk);
  dff _80969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _38972_, clk);
  dff _80970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _38973_, clk);
  dff _80971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _38974_, clk);
  dff _80972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _38975_, clk);
  dff _80973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _38960_, clk);
  dff _80974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _38961_, clk);
  dff _80975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _38962_, clk);
  dff _80976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _38963_, clk);
  dff _80977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _38964_, clk);
  dff _80978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _38965_, clk);
  dff _80979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _38966_, clk);
  dff _80980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _38967_, clk);
  dff _80981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _37168_, clk);
  dff _80982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _37169_, clk);
  dff _80983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _37170_, clk);
  dff _80984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _37171_, clk);
  dff _80985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _37172_, clk);
  dff _80986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _37173_, clk);
  dff _80987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _37174_, clk);
  dff _80988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _37175_, clk);
  dff _80989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _38952_, clk);
  dff _80990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _38953_, clk);
  dff _80991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _38954_, clk);
  dff _80992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _38955_, clk);
  dff _80993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _38956_, clk);
  dff _80994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _38957_, clk);
  dff _80995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _38958_, clk);
  dff _80996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _38959_, clk);
  dff _80997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _38944_, clk);
  dff _80998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _38945_, clk);
  dff _80999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _38946_, clk);
  dff _81000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _38947_, clk);
  dff _81001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _38948_, clk);
  dff _81002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _38949_, clk);
  dff _81003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _38950_, clk);
  dff _81004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _38951_, clk);
  dff _81005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _37160_, clk);
  dff _81006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _37161_, clk);
  dff _81007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _37162_, clk);
  dff _81008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _37163_, clk);
  dff _81009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _37164_, clk);
  dff _81010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _37165_, clk);
  dff _81011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _37166_, clk);
  dff _81012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _37167_, clk);
  dff _81013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _38936_, clk);
  dff _81014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _38937_, clk);
  dff _81015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _38938_, clk);
  dff _81016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _38939_, clk);
  dff _81017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _38940_, clk);
  dff _81018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _38941_, clk);
  dff _81019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _38942_, clk);
  dff _81020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _38943_, clk);
  dff _81021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _38928_, clk);
  dff _81022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _38929_, clk);
  dff _81023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _38930_, clk);
  dff _81024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _38931_, clk);
  dff _81025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _38932_, clk);
  dff _81026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _38933_, clk);
  dff _81027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _38934_, clk);
  dff _81028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _38935_, clk);
  dff _81029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _38232_, clk);
  dff _81030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _38233_, clk);
  dff _81031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _38234_, clk);
  dff _81032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _38235_, clk);
  dff _81033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _38236_, clk);
  dff _81034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _38237_, clk);
  dff _81035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _38238_, clk);
  dff _81036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _38239_, clk);
  dff _81037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _38240_, clk);
  dff _81038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _38241_, clk);
  dff _81039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _38242_, clk);
  dff _81040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _38243_, clk);
  dff _81041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _38244_, clk);
  dff _81042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _38245_, clk);
  dff _81043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _38246_, clk);
  dff _81044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _38247_, clk);
  dff _81045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _38136_, clk);
  dff _81046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _38137_, clk);
  dff _81047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _38138_, clk);
  dff _81048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _38139_, clk);
  dff _81049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _38140_, clk);
  dff _81050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _38141_, clk);
  dff _81051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _38142_, clk);
  dff _81052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _38143_, clk);
  dff _81053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _38144_, clk);
  dff _81054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _38145_, clk);
  dff _81055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _38146_, clk);
  dff _81056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _38147_, clk);
  dff _81057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _38148_, clk);
  dff _81058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _38149_, clk);
  dff _81059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _38150_, clk);
  dff _81060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _38151_, clk);
  dff _81061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _37944_, clk);
  dff _81062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _37945_, clk);
  dff _81063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _37946_, clk);
  dff _81064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _37947_, clk);
  dff _81065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _37948_, clk);
  dff _81066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _37949_, clk);
  dff _81067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _37950_, clk);
  dff _81068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _37951_, clk);
  dff _81069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _37616_, clk);
  dff _81070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _37617_, clk);
  dff _81071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _37618_, clk);
  dff _81072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _37619_, clk);
  dff _81073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _37620_, clk);
  dff _81074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _37621_, clk);
  dff _81075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _37622_, clk);
  dff _81076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _37623_, clk);
  dff _81077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _37552_, clk);
  dff _81078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _37553_, clk);
  dff _81079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _37554_, clk);
  dff _81080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _37555_, clk);
  dff _81081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _37556_, clk);
  dff _81082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _37557_, clk);
  dff _81083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _37558_, clk);
  dff _81084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _37559_, clk);
  dff _81085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _37152_, clk);
  dff _81086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _37153_, clk);
  dff _81087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _37154_, clk);
  dff _81088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _37155_, clk);
  dff _81089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _37156_, clk);
  dff _81090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _37157_, clk);
  dff _81091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _37158_, clk);
  dff _81092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _37159_, clk);
  dff _81093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _37144_, clk);
  dff _81094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _37145_, clk);
  dff _81095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _37146_, clk);
  dff _81096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _37147_, clk);
  dff _81097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _37148_, clk);
  dff _81098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _37149_, clk);
  dff _81099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _37150_, clk);
  dff _81100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _37151_, clk);
  dff _81101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _37608_, clk);
  dff _81102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _37609_, clk);
  dff _81103_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _37610_, clk);
  dff _81104_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _37611_, clk);
  dff _81105_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _37612_, clk);
  dff _81106_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _37613_, clk);
  dff _81107_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _37614_, clk);
  dff _81108_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _37615_, clk);
  dff _81109_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _37592_, clk);
  dff _81110_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _37593_, clk);
  dff _81111_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _37594_, clk);
  dff _81112_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _37595_, clk);
  dff _81113_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _37596_, clk);
  dff _81114_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _37597_, clk);
  dff _81115_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _37598_, clk);
  dff _81116_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _37599_, clk);
  dff _81117_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _37600_, clk);
  dff _81118_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _37601_, clk);
  dff _81119_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _37602_, clk);
  dff _81120_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _37603_, clk);
  dff _81121_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _37604_, clk);
  dff _81122_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _37605_, clk);
  dff _81123_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _37606_, clk);
  dff _81124_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _37607_, clk);
  dff _81125_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _37576_, clk);
  dff _81126_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _37577_, clk);
  dff _81127_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _37578_, clk);
  dff _81128_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _37579_, clk);
  dff _81129_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _37580_, clk);
  dff _81130_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _37581_, clk);
  dff _81131_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _37582_, clk);
  dff _81132_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _37583_, clk);
  dff _81133_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _37584_, clk);
  dff _81134_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _37585_, clk);
  dff _81135_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _37586_, clk);
  dff _81136_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _37587_, clk);
  dff _81137_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _37588_, clk);
  dff _81138_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _37589_, clk);
  dff _81139_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _37590_, clk);
  dff _81140_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _37591_, clk);
  dff _81141_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _37560_, clk);
  dff _81142_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _37561_, clk);
  dff _81143_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _37562_, clk);
  dff _81144_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _37563_, clk);
  dff _81145_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _37564_, clk);
  dff _81146_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _37565_, clk);
  dff _81147_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _37566_, clk);
  dff _81148_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _37567_, clk);
  dff _81149_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _37568_, clk);
  dff _81150_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _37569_, clk);
  dff _81151_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _37570_, clk);
  dff _81152_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _37571_, clk);
  dff _81153_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _37572_, clk);
  dff _81154_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _37573_, clk);
  dff _81155_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _37574_, clk);
  dff _81156_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _37575_, clk);
  dff _81157_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _37536_, clk);
  dff _81158_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _37537_, clk);
  dff _81159_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _37538_, clk);
  dff _81160_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _37539_, clk);
  dff _81161_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _37540_, clk);
  dff _81162_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _37541_, clk);
  dff _81163_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _37542_, clk);
  dff _81164_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _37543_, clk);
  dff _81165_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _37528_, clk);
  dff _81166_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _37529_, clk);
  dff _81167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _37530_, clk);
  dff _81168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _37531_, clk);
  dff _81169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _37532_, clk);
  dff _81170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _37533_, clk);
  dff _81171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _37534_, clk);
  dff _81172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _37535_, clk);
  dff _81173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _37520_, clk);
  dff _81174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _37521_, clk);
  dff _81175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _37522_, clk);
  dff _81176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _37523_, clk);
  dff _81177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _37524_, clk);
  dff _81178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _37525_, clk);
  dff _81179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _37526_, clk);
  dff _81180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _37527_, clk);
  dff _81181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _37232_, clk);
  dff _81182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _37233_, clk);
  dff _81183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _37234_, clk);
  dff _81184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _37235_, clk);
  dff _81185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _37236_, clk);
  dff _81186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _37237_, clk);
  dff _81187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _37238_, clk);
  dff _81188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _37239_, clk);
  dff _81189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _37240_, clk);
  dff _81190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _37241_, clk);
  dff _81191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _37242_, clk);
  dff _81192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _37243_, clk);
  dff _81193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _37244_, clk);
  dff _81194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _37245_, clk);
  dff _81195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _37246_, clk);
  dff _81196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _37247_, clk);
  dff _81197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _37224_, clk);
  dff _81198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _37225_, clk);
  dff _81199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _37226_, clk);
  dff _81200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _37227_, clk);
  dff _81201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _37228_, clk);
  dff _81202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _37229_, clk);
  dff _81203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _37230_, clk);
  dff _81204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _37231_, clk);
  dff _81205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _37216_, clk);
  dff _81206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _37217_, clk);
  dff _81207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _37218_, clk);
  dff _81208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _37219_, clk);
  dff _81209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _37220_, clk);
  dff _81210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _37221_, clk);
  dff _81211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _37222_, clk);
  dff _81212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _37223_, clk);
  dff _81213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _37208_, clk);
  dff _81214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _37209_, clk);
  dff _81215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _37210_, clk);
  dff _81216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _37211_, clk);
  dff _81217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _37212_, clk);
  dff _81218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _37213_, clk);
  dff _81219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _37214_, clk);
  dff _81220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _37215_, clk);
  dff _81221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [0], _38312_, clk);
  dff _81222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [1], _38313_, clk);
  dff _81223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [2], _38314_, clk);
  dff _81224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [3], _38315_, clk);
  dff _81225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [4], _38316_, clk);
  dff _81226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [5], _38317_, clk);
  dff _81227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [6], _38318_, clk);
  dff _81228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [7], _38319_, clk);
  dff _81229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _38304_, clk);
  dff _81230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _38305_, clk);
  dff _81231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _38306_, clk);
  dff _81232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _38307_, clk);
  dff _81233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _38308_, clk);
  dff _81234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _38309_, clk);
  dff _81235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _38310_, clk);
  dff _81236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _38311_, clk);
  dff _81237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _38288_, clk);
  dff _81238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _38289_, clk);
  dff _81239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _38290_, clk);
  dff _81240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _38291_, clk);
  dff _81241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _38292_, clk);
  dff _81242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _38293_, clk);
  dff _81243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _38294_, clk);
  dff _81244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _38295_, clk);
  dff _81245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _38296_, clk);
  dff _81246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _38297_, clk);
  dff _81247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _38298_, clk);
  dff _81248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _38299_, clk);
  dff _81249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _38300_, clk);
  dff _81250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _38301_, clk);
  dff _81251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _38302_, clk);
  dff _81252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _38303_, clk);
  dff _81253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _38280_, clk);
  dff _81254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _38281_, clk);
  dff _81255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _38282_, clk);
  dff _81256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _38283_, clk);
  dff _81257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _38284_, clk);
  dff _81258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _38285_, clk);
  dff _81259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _38286_, clk);
  dff _81260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _38287_, clk);
  dff _81261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _38272_, clk);
  dff _81262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _38273_, clk);
  dff _81263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _38274_, clk);
  dff _81264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _38275_, clk);
  dff _81265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _38276_, clk);
  dff _81266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _38277_, clk);
  dff _81267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _38278_, clk);
  dff _81268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _38279_, clk);
  dff _81269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _38248_, clk);
  dff _81270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _38249_, clk);
  dff _81271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _38250_, clk);
  dff _81272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _38251_, clk);
  dff _81273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _38252_, clk);
  dff _81274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _38253_, clk);
  dff _81275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _38254_, clk);
  dff _81276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _38255_, clk);
  dff _81277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _38264_, clk);
  dff _81278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _38265_, clk);
  dff _81279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _38266_, clk);
  dff _81280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _38267_, clk);
  dff _81281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _38268_, clk);
  dff _81282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _38269_, clk);
  dff _81283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _38270_, clk);
  dff _81284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _38271_, clk);
  dff _81285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _38224_, clk);
  dff _81286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _38225_, clk);
  dff _81287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _38226_, clk);
  dff _81288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _38227_, clk);
  dff _81289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _38228_, clk);
  dff _81290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _38229_, clk);
  dff _81291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _38230_, clk);
  dff _81292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _38231_, clk);
  dff _81293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _38216_, clk);
  dff _81294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _38217_, clk);
  dff _81295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _38218_, clk);
  dff _81296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _38219_, clk);
  dff _81297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _38220_, clk);
  dff _81298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _38221_, clk);
  dff _81299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _38222_, clk);
  dff _81300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _38223_, clk);
  dff _81301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _38200_, clk);
  dff _81302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _38201_, clk);
  dff _81303_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _38202_, clk);
  dff _81304_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _38203_, clk);
  dff _81305_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _38204_, clk);
  dff _81306_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _38205_, clk);
  dff _81307_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _38206_, clk);
  dff _81308_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _38207_, clk);
  dff _81309_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _38208_, clk);
  dff _81310_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _38209_, clk);
  dff _81311_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _38210_, clk);
  dff _81312_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _38211_, clk);
  dff _81313_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _38212_, clk);
  dff _81314_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _38213_, clk);
  dff _81315_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _38214_, clk);
  dff _81316_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _38215_, clk);
  dff _81317_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _38192_, clk);
  dff _81318_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _38193_, clk);
  dff _81319_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _38194_, clk);
  dff _81320_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _38195_, clk);
  dff _81321_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _38196_, clk);
  dff _81322_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _38197_, clk);
  dff _81323_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _38198_, clk);
  dff _81324_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _38199_, clk);
  dff _81325_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _38184_, clk);
  dff _81326_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _38185_, clk);
  dff _81327_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _38186_, clk);
  dff _81328_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _38187_, clk);
  dff _81329_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _38188_, clk);
  dff _81330_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _38189_, clk);
  dff _81331_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _38190_, clk);
  dff _81332_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _38191_, clk);
  dff _81333_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _38176_, clk);
  dff _81334_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _38177_, clk);
  dff _81335_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _38178_, clk);
  dff _81336_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _38179_, clk);
  dff _81337_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _38180_, clk);
  dff _81338_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _38181_, clk);
  dff _81339_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _38182_, clk);
  dff _81340_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _38183_, clk);
  dff _81341_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _38160_, clk);
  dff _81342_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _38161_, clk);
  dff _81343_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _38162_, clk);
  dff _81344_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _38163_, clk);
  dff _81345_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _38164_, clk);
  dff _81346_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _38165_, clk);
  dff _81347_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _38166_, clk);
  dff _81348_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _38167_, clk);
  dff _81349_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _38152_, clk);
  dff _81350_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _38153_, clk);
  dff _81351_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _38154_, clk);
  dff _81352_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _38155_, clk);
  dff _81353_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _38156_, clk);
  dff _81354_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _38157_, clk);
  dff _81355_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _38158_, clk);
  dff _81356_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _38159_, clk);
  dff _81357_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _38120_, clk);
  dff _81358_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _38121_, clk);
  dff _81359_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _38122_, clk);
  dff _81360_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _38123_, clk);
  dff _81361_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _38124_, clk);
  dff _81362_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _38125_, clk);
  dff _81363_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _38126_, clk);
  dff _81364_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _38127_, clk);
  dff _81365_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _38128_, clk);
  dff _81366_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _38129_, clk);
  dff _81367_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _38130_, clk);
  dff _81368_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _38131_, clk);
  dff _81369_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _38132_, clk);
  dff _81370_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _38133_, clk);
  dff _81371_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _38134_, clk);
  dff _81372_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _38135_, clk);
  dff _81373_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _38112_, clk);
  dff _81374_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _38113_, clk);
  dff _81375_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _38114_, clk);
  dff _81376_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _38115_, clk);
  dff _81377_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _38116_, clk);
  dff _81378_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _38117_, clk);
  dff _81379_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _38118_, clk);
  dff _81380_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _38119_, clk);
  dff _81381_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _38104_, clk);
  dff _81382_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _38105_, clk);
  dff _81383_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _38106_, clk);
  dff _81384_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _38107_, clk);
  dff _81385_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _38108_, clk);
  dff _81386_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _38109_, clk);
  dff _81387_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _38110_, clk);
  dff _81388_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _38111_, clk);
  dff _81389_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _38096_, clk);
  dff _81390_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _38097_, clk);
  dff _81391_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _38098_, clk);
  dff _81392_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _38099_, clk);
  dff _81393_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _38100_, clk);
  dff _81394_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _38101_, clk);
  dff _81395_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _38102_, clk);
  dff _81396_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _38103_, clk);
  dff _81397_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _38088_, clk);
  dff _81398_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _38089_, clk);
  dff _81399_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _38090_, clk);
  dff _81400_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _38091_, clk);
  dff _81401_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _38092_, clk);
  dff _81402_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _38093_, clk);
  dff _81403_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _38094_, clk);
  dff _81404_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _38095_, clk);
  dff _81405_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _38072_, clk);
  dff _81406_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _38073_, clk);
  dff _81407_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _38074_, clk);
  dff _81408_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _38075_, clk);
  dff _81409_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _38076_, clk);
  dff _81410_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _38077_, clk);
  dff _81411_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _38078_, clk);
  dff _81412_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _38079_, clk);
  dff _81413_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _38040_, clk);
  dff _81414_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _38041_, clk);
  dff _81415_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _38042_, clk);
  dff _81416_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _38043_, clk);
  dff _81417_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _38044_, clk);
  dff _81418_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _38045_, clk);
  dff _81419_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _38046_, clk);
  dff _81420_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _38047_, clk);
  dff _81421_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _38032_, clk);
  dff _81422_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _38033_, clk);
  dff _81423_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _38034_, clk);
  dff _81424_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _38035_, clk);
  dff _81425_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _38036_, clk);
  dff _81426_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _38037_, clk);
  dff _81427_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _38038_, clk);
  dff _81428_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _38039_, clk);
  dff _81429_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _38024_, clk);
  dff _81430_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _38025_, clk);
  dff _81431_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _38026_, clk);
  dff _81432_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _38027_, clk);
  dff _81433_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _38028_, clk);
  dff _81434_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _38029_, clk);
  dff _81435_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _38030_, clk);
  dff _81436_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _38031_, clk);
  dff _81437_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _37936_, clk);
  dff _81438_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _37937_, clk);
  dff _81439_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _37938_, clk);
  dff _81440_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _37939_, clk);
  dff _81441_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _37940_, clk);
  dff _81442_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _37941_, clk);
  dff _81443_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _37942_, clk);
  dff _81444_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _37943_, clk);
  dff _81445_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _37968_, clk);
  dff _81446_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _37969_, clk);
  dff _81447_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _37970_, clk);
  dff _81448_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _37971_, clk);
  dff _81449_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _37972_, clk);
  dff _81450_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _37973_, clk);
  dff _81451_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _37974_, clk);
  dff _81452_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _37975_, clk);
  dff _81453_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _37952_, clk);
  dff _81454_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _37953_, clk);
  dff _81455_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _37954_, clk);
  dff _81456_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _37955_, clk);
  dff _81457_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _37956_, clk);
  dff _81458_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _37957_, clk);
  dff _81459_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _37958_, clk);
  dff _81460_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _37959_, clk);
  dff _81461_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _37960_, clk);
  dff _81462_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _37961_, clk);
  dff _81463_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _37962_, clk);
  dff _81464_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _37963_, clk);
  dff _81465_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _37964_, clk);
  dff _81466_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _37965_, clk);
  dff _81467_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _37966_, clk);
  dff _81468_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _37967_, clk);
  dff _81469_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _38984_[0], clk);
  dff _81470_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _38984_[1], clk);
  dff _81471_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _38984_[2], clk);
  dff _81472_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _38984_[3], clk);
  dff _81473_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _38984_[4], clk);
  dff _81474_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _38984_[5], clk);
  dff _81475_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _38984_[6], clk);
  dff _81476_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _38984_[7], clk);
  dff _81477_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0], clk);
  dff _81478_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1], clk);
  dff _81479_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2], clk);
  dff _81480_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3], clk);
  dff _81481_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4], clk);
  dff _81482_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5], clk);
  dff _81483_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6], clk);
  dff _81484_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7], clk);
  dff _81485_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8], clk);
  dff _81486_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9], clk);
  dff _81487_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10], clk);
  dff _81488_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11], clk);
  dff _81489_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12], clk);
  dff _81490_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13], clk);
  dff _81491_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14], clk);
  dff _81492_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15], clk);
  dff _81493_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16], clk);
  dff _81494_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17], clk);
  dff _81495_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18], clk);
  dff _81496_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19], clk);
  dff _81497_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20], clk);
  dff _81498_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21], clk);
  dff _81499_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22], clk);
  dff _81500_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23], clk);
  dff _81501_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24], clk);
  dff _81502_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25], clk);
  dff _81503_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26], clk);
  dff _81504_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27], clk);
  dff _81505_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28], clk);
  dff _81506_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29], clk);
  dff _81507_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30], clk);
  dff _81508_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31], clk);
  dff _81509_ (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1, clk);
  dff _81510_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _38985_, clk);
  dff _81511_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _38986_[0], clk);
  dff _81512_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _38986_[1], clk);
  dff _81513_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _38986_[2], clk);
  dff _81514_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _38986_[3], clk);
  dff _81515_ (\oc8051_top_1.oc8051_sfr1.bit_out , _38987_, clk);
  dff _81516_ (\oc8051_top_1.oc8051_sfr1.wait_data , _38988_, clk);
  dff _81517_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _38989_[0], clk);
  dff _81518_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _38989_[1], clk);
  dff _81519_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _38989_[2], clk);
  dff _81520_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _38989_[3], clk);
  dff _81521_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _38989_[4], clk);
  dff _81522_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _38989_[5], clk);
  dff _81523_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _38989_[6], clk);
  dff _81524_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _38989_[7], clk);
  dff _81525_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _38990_, clk);
  dff _81526_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _38991_[0], clk);
  dff _81527_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _38991_[1], clk);
  dff _81528_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _38991_[2], clk);
  dff _81529_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _38991_[3], clk);
  dff _81530_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _38991_[4], clk);
  dff _81531_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _38991_[5], clk);
  dff _81532_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _38991_[6], clk);
  dff _81533_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _38991_[7], clk);
  dff _81534_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _38992_[0], clk);
  dff _81535_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _38992_[1], clk);
  dff _81536_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _38992_[2], clk);
  dff _81537_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _38992_[3], clk);
  dff _81538_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _38992_[4], clk);
  dff _81539_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _38992_[5], clk);
  dff _81540_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _38992_[6], clk);
  dff _81541_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _38992_[7], clk);
  dff _81542_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _38993_[0], clk);
  dff _81543_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _38993_[1], clk);
  dff _81544_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _38993_[2], clk);
  dff _81545_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _38993_[3], clk);
  dff _81546_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _38993_[4], clk);
  dff _81547_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _38993_[5], clk);
  dff _81548_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _38993_[6], clk);
  dff _81549_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _38993_[7], clk);
  dff _81550_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _38994_[0], clk);
  dff _81551_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _38994_[1], clk);
  dff _81552_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _38994_[2], clk);
  dff _81553_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _38994_[3], clk);
  dff _81554_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _38994_[4], clk);
  dff _81555_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _38994_[5], clk);
  dff _81556_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _38994_[6], clk);
  dff _81557_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _38994_[7], clk);
  dff _81558_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _38995_, clk);
  dff _81559_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _38996_, clk);
  dff _81560_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0, clk);
  dff _81561_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _38997_, clk);
  dff _81562_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _38998_[0], clk);
  dff _81563_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _38998_[1], clk);
  dff _81564_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _38998_[2], clk);
  dff _81565_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _38998_[3], clk);
  dff _81566_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _38998_[4], clk);
  dff _81567_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _38998_[5], clk);
  dff _81568_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _38998_[6], clk);
  dff _81569_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _38998_[7], clk);
  dff _81570_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _38999_[0], clk);
  dff _81571_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _38999_[1], clk);
  dff _81572_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _39000_, clk);
  dff _81573_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _39001_[0], clk);
  dff _81574_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _39001_[1], clk);
  dff _81575_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _39001_[2], clk);
  dff _81576_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _39002_[0], clk);
  dff _81577_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _39002_[1], clk);
  dff _81578_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _39002_[2], clk);
  dff _81579_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _39003_[0], clk);
  dff _81580_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _39003_[1], clk);
  dff _81581_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _39004_[0], clk);
  dff _81582_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _39004_[1], clk);
  dff _81583_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _39005_, clk);
  dff _81584_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _39006_, clk);
  dff _81585_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _39007_, clk);
  dff _81586_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _39008_, clk);
  dff _81587_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _39009_[0], clk);
  dff _81588_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _39009_[1], clk);
  dff _81589_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _39009_[2], clk);
  dff _81590_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _39009_[3], clk);
  dff _81591_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _39010_[0], clk);
  dff _81592_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _39010_[1], clk);
  dff _81593_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _39010_[2], clk);
  dff _81594_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _39010_[3], clk);
  dff _81595_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _39010_[4], clk);
  dff _81596_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _39010_[5], clk);
  dff _81597_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _39010_[6], clk);
  dff _81598_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _39010_[7], clk);
  dff _81599_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _39011_[0], clk);
  dff _81600_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _39011_[1], clk);
  dff _81601_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _39011_[2], clk);
  dff _81602_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _39011_[3], clk);
  dff _81603_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _39011_[4], clk);
  dff _81604_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _39011_[5], clk);
  dff _81605_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _39011_[6], clk);
  dff _81606_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _39011_[7], clk);
  dff _81607_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _39012_[0], clk);
  dff _81608_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _39012_[1], clk);
  dff _81609_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _39012_[2], clk);
  dff _81610_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _39012_[3], clk);
  dff _81611_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _39012_[4], clk);
  dff _81612_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _39012_[5], clk);
  dff _81613_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _39012_[6], clk);
  dff _81614_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _39012_[7], clk);
  dff _81615_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _39013_[0], clk);
  dff _81616_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _39013_[1], clk);
  dff _81617_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _39013_[2], clk);
  dff _81618_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _39013_[3], clk);
  dff _81619_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _39013_[4], clk);
  dff _81620_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _39013_[5], clk);
  dff _81621_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _39013_[6], clk);
  dff _81622_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _39013_[7], clk);
  dff _81623_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _39014_[0], clk);
  dff _81624_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _39014_[1], clk);
  dff _81625_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _39014_[2], clk);
  dff _81626_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _39014_[3], clk);
  dff _81627_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _39014_[4], clk);
  dff _81628_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _39014_[5], clk);
  dff _81629_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _39014_[6], clk);
  dff _81630_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _39014_[7], clk);
  dff _81631_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _39015_[0], clk);
  dff _81632_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _39015_[1], clk);
  dff _81633_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _39015_[2], clk);
  dff _81634_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _39015_[3], clk);
  dff _81635_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _39015_[4], clk);
  dff _81636_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _39015_[5], clk);
  dff _81637_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _39015_[6], clk);
  dff _81638_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _39015_[7], clk);
  dff _81639_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _39016_[0], clk);
  dff _81640_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _39016_[1], clk);
  dff _81641_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _39016_[2], clk);
  dff _81642_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _39016_[3], clk);
  dff _81643_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _39016_[4], clk);
  dff _81644_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _39016_[5], clk);
  dff _81645_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _39016_[6], clk);
  dff _81646_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _39017_, clk);
  dff _81647_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _39018_[0], clk);
  dff _81648_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _39018_[1], clk);
  dff _81649_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _39018_[2], clk);
  dff _81650_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _39018_[3], clk);
  dff _81651_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _39018_[4], clk);
  dff _81652_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _39018_[5], clk);
  dff _81653_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _39018_[6], clk);
  dff _81654_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _39018_[7], clk);
  dff _81655_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _39019_, clk);
  dff _81656_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _39020_, clk);
  dff _81657_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _39021_[0], clk);
  dff _81658_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _39021_[1], clk);
  dff _81659_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _39021_[2], clk);
  dff _81660_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _39021_[3], clk);
  dff _81661_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _39021_[4], clk);
  dff _81662_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _39021_[5], clk);
  dff _81663_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _39021_[6], clk);
  dff _81664_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _39021_[7], clk);
  dff _81665_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _39022_[0], clk);
  dff _81666_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _39022_[1], clk);
  dff _81667_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _39022_[2], clk);
  dff _81668_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _39022_[3], clk);
  dff _81669_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _39022_[4], clk);
  dff _81670_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _39022_[5], clk);
  dff _81671_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _39022_[6], clk);
  dff _81672_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _39022_[7], clk);
  dff _81673_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _39023_, clk);
  dff _81674_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _39024_, clk);
  dff _81675_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _39025_[0], clk);
  dff _81676_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _39025_[1], clk);
  dff _81677_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _39025_[2], clk);
  dff _81678_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _39025_[3], clk);
  dff _81679_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _39025_[4], clk);
  dff _81680_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _39025_[5], clk);
  dff _81681_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _39025_[6], clk);
  dff _81682_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _39025_[7], clk);
  dff _81683_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _39026_[0], clk);
  dff _81684_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _39026_[1], clk);
  dff _81685_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _39026_[2], clk);
  dff _81686_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _39026_[3], clk);
  dff _81687_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _39026_[4], clk);
  dff _81688_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _39026_[5], clk);
  dff _81689_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _39026_[6], clk);
  dff _81690_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _39026_[7], clk);
  dff _81691_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _39027_, clk);
  dff _81692_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _39028_[0], clk);
  dff _81693_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _39028_[1], clk);
  dff _81694_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _39028_[2], clk);
  dff _81695_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _39028_[3], clk);
  dff _81696_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _39028_[4], clk);
  dff _81697_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _39028_[5], clk);
  dff _81698_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _39028_[6], clk);
  dff _81699_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _39028_[7], clk);
  dff _81700_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _39029_, clk);
  dff _81701_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _39030_, clk);
  dff _81702_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _39031_, clk);
  dff _81703_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _39032_, clk);
  dff _81704_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _39033_[0], clk);
  dff _81705_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _39033_[1], clk);
  dff _81706_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _39033_[2], clk);
  dff _81707_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _39033_[3], clk);
  dff _81708_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _39033_[4], clk);
  dff _81709_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _39033_[5], clk);
  dff _81710_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _39033_[6], clk);
  dff _81711_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _39033_[7], clk);
  dff _81712_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _39034_[0], clk);
  dff _81713_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _39034_[1], clk);
  dff _81714_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _39034_[2], clk);
  dff _81715_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _39034_[3], clk);
  dff _81716_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _39034_[4], clk);
  dff _81717_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _39034_[5], clk);
  dff _81718_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _39034_[6], clk);
  dff _81719_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _39034_[7], clk);
  dff _81720_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _39035_, clk);
  dff _81721_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _39036_[0], clk);
  dff _81722_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _39036_[1], clk);
  dff _81723_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _39036_[2], clk);
  dff _81724_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _39036_[3], clk);
  dff _81725_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _39036_[4], clk);
  dff _81726_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _39036_[5], clk);
  dff _81727_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _39036_[6], clk);
  dff _81728_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _39036_[7], clk);
  dff _81729_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _39037_[0], clk);
  dff _81730_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _39037_[1], clk);
  dff _81731_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _39037_[2], clk);
  dff _81732_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _39037_[3], clk);
  dff _81733_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _39037_[4], clk);
  dff _81734_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _39037_[5], clk);
  dff _81735_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _39037_[6], clk);
  dff _81736_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _39037_[7], clk);
  dff _81737_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _39038_, clk);
  dff _81738_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _39039_[0], clk);
  dff _81739_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _39039_[1], clk);
  dff _81740_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _39039_[2], clk);
  dff _81741_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _39039_[3], clk);
  dff _81742_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _39039_[4], clk);
  dff _81743_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _39039_[5], clk);
  dff _81744_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _39039_[6], clk);
  dff _81745_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _39039_[7], clk);
  dff _81746_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _39049_[0], clk);
  dff _81747_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _39049_[1], clk);
  dff _81748_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _39049_[2], clk);
  dff _81749_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _39049_[3], clk);
  dff _81750_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _39049_[4], clk);
  dff _81751_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _39049_[5], clk);
  dff _81752_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _39049_[6], clk);
  dff _81753_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _39049_[7], clk);
  dff _81754_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _39049_[8], clk);
  dff _81755_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _39049_[9], clk);
  dff _81756_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _39049_[10], clk);
  dff _81757_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _39049_[11], clk);
  dff _81758_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _39040_, clk);
  dff _81759_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _39041_, clk);
  dff _81760_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _39042_, clk);
  dff _81761_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _39043_, clk);
  dff _81762_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _39044_, clk);
  dff _81763_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _39045_, clk);
  dff _81764_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _39046_[0], clk);
  dff _81765_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _39046_[1], clk);
  dff _81766_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _39047_[0], clk);
  dff _81767_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _39047_[1], clk);
  dff _81768_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _39047_[2], clk);
  dff _81769_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _39047_[3], clk);
  dff _81770_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _39048_[0], clk);
  dff _81771_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _39048_[1], clk);
  dff _81772_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _39048_[2], clk);
  dff _81773_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _39048_[3], clk);
  dff _81774_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _39048_[4], clk);
  dff _81775_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _39048_[5], clk);
  dff _81776_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _39048_[6], clk);
  dff _81777_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _39048_[7], clk);
  dff _81778_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _39050_, clk);
  dff _81779_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _39051_, clk);
  dff _81780_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _39052_, clk);
  dff _81781_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _39053_, clk);
  dff _81782_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _39054_, clk);
  dff _81783_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _39055_[0], clk);
  dff _81784_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _39055_[1], clk);
  dff _81785_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _39055_[2], clk);
  dff _81786_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _39055_[3], clk);
  dff _81787_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _39056_[0], clk);
  dff _81788_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _39056_[1], clk);
  dff _81789_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _39056_[2], clk);
  dff _81790_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _39056_[3], clk);
  dff _81791_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _39056_[4], clk);
  dff _81792_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _39056_[5], clk);
  dff _81793_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _39056_[6], clk);
  dff _81794_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _39056_[7], clk);
  dff _81795_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _39056_[8], clk);
  dff _81796_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _39056_[9], clk);
  dff _81797_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _39056_[10], clk);
  dff _81798_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _39057_[0], clk);
  dff _81799_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _39057_[1], clk);
  dff _81800_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _39057_[2], clk);
  dff _81801_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _39057_[3], clk);
  dff _81802_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _39057_[4], clk);
  dff _81803_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _39057_[5], clk);
  dff _81804_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _39057_[6], clk);
  dff _81805_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _39057_[7], clk);
  dff _81806_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _39058_[0], clk);
  dff _81807_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _39058_[1], clk);
  dff _81808_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _39058_[2], clk);
  dff _81809_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _39058_[3], clk);
  dff _81810_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _39058_[4], clk);
  dff _81811_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _39058_[5], clk);
  dff _81812_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _39058_[6], clk);
  dff _81813_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _39058_[7], clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 );
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 );
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 );
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 );
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 );
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 );
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.uart_int , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr );
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tc2_int , \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
